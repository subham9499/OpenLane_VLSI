* NGSPICE file created from Turn_Controller.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt Turn_Controller vdd gnd clock ped_Hori_Interrupt ped_Vert_Interrupt police_Interrupt
+ traffic_Street_0[0] traffic_Street_0[1] traffic_Street_0[2] traffic_Street_0[3]
+ traffic_Street_1[0] traffic_Street_1[1] traffic_Street_1[2] traffic_Street_1[3]
+ address[0] address[1] address[2] address[3] address[4] address[5] address[6] read_Write
+ enable street north_South[0] north_South[1] west_East[0] west_East[1] pedestrian_Hori_Street
+ pedestrian_Vert_Street traffic_Street[0] traffic_Street[1] traffic_Street[2] traffic_Street[3]
XFILL_9_6_0 gnd vdd FILL
XFILL_17_5_0 gnd vdd FILL
XAOI21X1_609 BUFX4_72/Y NOR2X1_231/B NOR2X1_721/Y gnd AOI21X1_609/Y vdd AOI21X1
XFILL_50_3_0 gnd vdd FILL
XFILL_41_3_0 gnd vdd FILL
XFILL_42_8_1 gnd vdd FILL
XOAI21X1_371 BUFX4_470/Y NAND2X1_2/Y NAND2X1_89/Y gnd DFFPOSX1_45/D vdd OAI21X1
XOAI21X1_382 BUFX4_294/Y BUFX4_299/Y NOR2X1_449/A gnd OAI21X1_382/Y vdd OAI21X1
XOAI21X1_360 BUFX4_188/Y BUFX4_197/Y NAND2X1_198/A gnd OAI21X1_361/C vdd OAI21X1
XINVX1_402 INVX1_402/A gnd INVX1_402/Y vdd INVX1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_393 BUFX4_448/Y BUFX4_294/Y NOR2X1_505/A gnd OAI21X1_393/Y vdd OAI21X1
XINVX1_413 INVX1_413/A gnd INVX1_413/Y vdd INVX1
XINVX1_424 INVX1_424/A gnd INVX1_424/Y vdd INVX1
XINVX1_435 INVX1_435/A gnd INVX1_435/Y vdd INVX1
XINVX1_457 INVX1_457/A gnd INVX1_457/Y vdd INVX1
XINVX1_446 INVX1_446/A gnd INVX1_446/Y vdd INVX1
XFILL_49_4_0 gnd vdd FILL
XFILL_32_3_0 gnd vdd FILL
XFILL_33_8_1 gnd vdd FILL
XAOI21X1_406 BUFX4_106/Y INVX1_362/Y BUFX4_265/Y gnd AOI21X1_406/Y vdd AOI21X1
XAOI21X1_439 INVX1_46/Y BUFX4_271/Y AOI21X1_439/C gnd AOI21X1_439/Y vdd AOI21X1
XAOI21X1_428 NAND2X1_7/A BUFX4_347/Y BUFX4_146/Y gnd OAI21X1_979/C vdd AOI21X1
XAOI21X1_417 BUFX4_283/Y INVX1_380/Y AOI21X1_417/C gnd AOI21X1_417/Y vdd AOI21X1
XFILL_23_3_0 gnd vdd FILL
XFILL_24_8_1 gnd vdd FILL
XFILL_7_9_1 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XMUX2X1_17 INVX1_22/Y BUFX4_442/Y MUX2X1_18/S gnd MUX2X1_17/Y vdd MUX2X1
XMUX2X1_28 INVX1_36/Y BUFX4_70/Y MUX2X1_29/S gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_39 INVX1_49/Y MUX2X1_39/B MUX2X1_42/S gnd MUX2X1_39/Y vdd MUX2X1
XFILL_15_8_1 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XOAI21X1_190 BUFX4_136/Y BUFX4_127/Y OAI21X1_190/C gnd OAI21X1_191/C vdd OAI21X1
XDFFPOSX1_509 NOR2X1_721/A CLKBUF1_16/Y AOI21X1_609/Y gnd vdd DFFPOSX1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_232 INVX1_232/A gnd INVX1_232/Y vdd INVX1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XINVX1_276 INVX1_276/A gnd INVX1_276/Y vdd INVX1
XINVX1_265 INVX1_265/A gnd INVX1_265/Y vdd INVX1
XINVX1_298 INVX1_298/A gnd INVX1_298/Y vdd INVX1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XNAND2X1_32 INVX8_12/A INVX4_5/Y gnd NAND2X1_32/Y vdd NAND2X1
XNAND2X1_21 NOR2X1_4/Y NOR2X1_10/Y gnd BUFX4_449/A vdd NAND2X1
XNAND2X1_10 NOR2X1_12/Y NOR2X1_6/Y gnd MUX2X1_18/S vdd NAND2X1
XNAND2X1_43 INVX8_18/A INVX4_2/Y gnd MUX2X1_70/S vdd NAND2X1
XNAND2X1_54 INVX8_19/A INVX4_5/Y gnd MUX2X1_81/S vdd NAND2X1
XNAND2X1_76 INVX8_25/A INVX4_3/Y gnd NAND2X1_76/Y vdd NAND2X1
XNAND2X1_65 INVX8_22/A INVX4_4/Y gnd MUX2X1_353/S vdd NAND2X1
XNAND2X1_98 traffic_Street_1[1] AOI21X1_7/B gnd NAND2X1_98/Y vdd NAND2X1
XNAND2X1_87 NAND2X1_87/A NAND2X1_2/Y gnd NAND2X1_87/Y vdd NAND2X1
XNOR2X1_601 NOR2X1_601/A BUFX4_225/Y gnd NOR2X1_601/Y vdd NOR2X1
XFILL_42_2 gnd vdd FILL
XNOR2X1_634 NOR2X1_634/A NOR2X1_65/Y gnd NOR2X1_634/Y vdd NOR2X1
XNOR2X1_623 BUFX4_39/Y MUX2X1_266/Y gnd NOR2X1_623/Y vdd NOR2X1
XNOR2X1_612 NOR2X1_204/A AND2X2_22/A gnd OAI22X1_87/D vdd NOR2X1
XNOR2X1_667 NOR2X1_667/A AOI21X1_72/B gnd NOR2X1_667/Y vdd NOR2X1
XNOR2X1_678 NOR2X1_678/A MUX2X1_94/S gnd NOR2X1_678/Y vdd NOR2X1
XNOR2X1_656 NOR2X1_656/A NOR2X1_107/B gnd NOR2X1_656/Y vdd NOR2X1
XNOR2X1_645 NOR2X1_645/A MUX2X1_55/S gnd NOR2X1_645/Y vdd NOR2X1
XFILL_35_1 gnd vdd FILL
XNOR2X1_689 NOR2X1_689/A MUX2X1_340/S gnd NOR2X1_689/Y vdd NOR2X1
XAOI21X1_203 NAND3X1_5/B NAND3X1_5/C NAND3X1_5/A gnd OAI21X1_441/A vdd AOI21X1
XAOI21X1_225 AOI21X1_225/A NOR2X1_341/B INVX1_198/Y gnd AOI21X1_225/Y vdd AOI21X1
XAOI21X1_214 NAND2X1_168/A INVX2_15/A INVX1_192/Y gnd OAI21X1_463/C vdd AOI21X1
XAOI21X1_236 NOR3X1_9/Y AND2X2_10/Y AOI21X1_235/Y gnd AOI21X1_236/Y vdd AOI21X1
XAOI21X1_258 BUFX4_237/Y NOR2X1_655/A BUFX4_85/Y gnd OAI21X1_569/C vdd AOI21X1
XAOI21X1_247 AND2X2_46/B INVX1_220/Y BUFX4_74/Y gnd AOI21X1_247/Y vdd AOI21X1
XAOI21X1_269 BUFX4_91/Y OAI21X1_588/Y AOI21X1_268/Y gnd OAI22X1_5/C vdd AOI21X1
XAOI22X1_30 AOI22X1_30/A AOI22X1_30/B AOI22X1_30/C BUFX4_171/Y gnd AOI22X1_30/Y vdd
+ AOI22X1
XOAI21X1_1420 BUFX4_119/Y BUFX4_408/Y OAI21X1_1116/B gnd OAI21X1_1421/C vdd OAI21X1
XOAI21X1_1431 NAND2X1_66/Y BUFX4_437/Y OAI21X1_1431/C gnd OAI21X1_1431/Y vdd OAI21X1
XOAI21X1_1442 BUFX4_60/Y BUFX4_435/Y OAI21X1_957/B gnd OAI21X1_1442/Y vdd OAI21X1
XOAI21X1_1464 NAND2X1_70/Y MUX2X1_29/B OAI21X1_1463/Y gnd OAI21X1_1464/Y vdd OAI21X1
XOAI21X1_1453 NAND2X1_69/Y MUX2X1_29/B OAI21X1_1453/C gnd DFFPOSX1_293/D vdd OAI21X1
XOAI21X1_1475 BUFX4_132/Y BUFX4_162/Y INVX1_319/A gnd OAI21X1_1475/Y vdd OAI21X1
XOAI21X1_1497 BUFX4_386/Y BUFX4_456/Y INVX1_265/A gnd OAI21X1_1498/C vdd OAI21X1
XOAI21X1_1486 BUFX4_66/Y NAND2X1_74/Y OAI21X1_1486/C gnd OAI21X1_1486/Y vdd OAI21X1
XDFFPOSX1_1027 INVX1_141/A CLKBUF1_57/Y MUX2X1_128/Y gnd vdd DFFPOSX1
XDFFPOSX1_1005 NOR2X1_518/A CLKBUF1_79/Y OAI21X1_293/Y gnd vdd DFFPOSX1
XDFFPOSX1_1016 NOR2X1_460/A CLKBUF1_60/Y AOI21X1_145/Y gnd vdd DFFPOSX1
XDFFPOSX1_1038 INVX1_445/A CLKBUF1_64/Y OAI21X1_319/Y gnd vdd DFFPOSX1
XDFFPOSX1_1049 NOR2X1_248/A CLKBUF1_67/Y AOI21X1_158/Y gnd vdd DFFPOSX1
XOAI22X1_3 OAI22X1_3/A INVX4_12/A OAI22X1_3/C OAI22X1_3/D gnd AND2X2_16/A vdd OAI22X1
XFILL_47_7_1 gnd vdd FILL
XFILL_46_2_0 gnd vdd FILL
XFILL_30_6_1 gnd vdd FILL
XDFFPOSX1_306 INVX1_250/A CLKBUF1_97/Y DFFPOSX1_306/D gnd vdd DFFPOSX1
XDFFPOSX1_317 INVX1_413/A CLKBUF1_48/Y MUX2X1_287/Y gnd vdd DFFPOSX1
XDFFPOSX1_328 INVX1_370/A CLKBUF1_74/Y DFFPOSX1_328/D gnd vdd DFFPOSX1
XDFFPOSX1_339 NOR2X1_656/A CLKBUF1_87/Y AOI21X1_544/Y gnd vdd DFFPOSX1
XFILL_37_2_0 gnd vdd FILL
XFILL_38_7_1 gnd vdd FILL
XBUFX4_382 BUFX4_384/A gnd INVX4_3/A vdd BUFX4
XBUFX4_360 BUFX4_26/Y gnd BUFX4_360/Y vdd BUFX4
XBUFX4_371 INVX8_14/Y gnd BUFX4_371/Y vdd BUFX4
XNOR2X1_442 OAI21X1_12/C BUFX4_246/Y gnd NOR2X1_442/Y vdd NOR2X1
XNOR2X1_420 BUFX4_112/Y NOR2X1_420/B gnd NOR2X1_420/Y vdd NOR2X1
XBUFX4_393 INVX8_28/Y gnd BUFX4_393/Y vdd BUFX4
XNOR2X1_431 NOR2X1_431/A BUFX4_331/Y gnd NOR2X1_431/Y vdd NOR2X1
XNOR2X1_464 NOR2X1_464/A AND2X2_22/A gnd OAI22X1_33/D vdd NOR2X1
XNOR2X1_475 NOR2X1_475/A NOR2X1_475/B gnd NOR2X1_475/Y vdd NOR2X1
XNOR2X1_453 NOR2X1_453/A BUFX4_287/Y gnd NOR2X1_453/Y vdd NOR2X1
XNOR2X1_486 NOR2X1_486/A BUFX4_350/Y gnd NOR2X1_486/Y vdd NOR2X1
XNOR2X1_497 BUFX4_39/Y MUX2X1_244/Y gnd NOR2X1_497/Y vdd NOR2X1
XFILL_20_1_0 gnd vdd FILL
XFILL_21_6_1 gnd vdd FILL
XOAI21X1_915 BUFX4_365/Y INVX1_346/Y OAI21X1_915/C gnd OAI21X1_915/Y vdd OAI21X1
XOAI21X1_904 BUFX4_345/Y OAI21X1_274/C BUFX4_152/Y gnd OAI22X1_35/C vdd OAI21X1
XOAI21X1_948 INVX1_372/Y BUFX4_274/Y NAND2X1_283/Y gnd MUX2X1_233/B vdd OAI21X1
XOAI21X1_926 INVX1_356/Y BUFX4_93/Y BUFX4_263/Y gnd OAI21X1_926/Y vdd OAI21X1
XOAI21X1_937 BUFX4_35/Y INVX1_365/Y BUFX4_328/Y gnd OAI21X1_937/Y vdd OAI21X1
XOAI21X1_959 OAI21X1_959/A AOI21X1_417/Y BUFX4_33/Y gnd AOI21X1_420/A vdd OAI21X1
XMUX2X1_404 INVX1_270/Y BUFX4_442/Y MUX2X1_406/S gnd MUX2X1_404/Y vdd MUX2X1
XDFFPOSX1_851 OAI21X1_686/A CLKBUF1_53/Y OAI21X1_177/Y gnd vdd DFFPOSX1
XOAI21X1_1283 BUFX4_124/Y BUFX4_43/Y OAI21X1_741/B gnd OAI21X1_1283/Y vdd OAI21X1
XOAI21X1_1272 NAND2X1_30/Y BUFX4_321/Y OAI21X1_1272/C gnd DFFPOSX1_241/D vdd OAI21X1
XDFFPOSX1_840 INVX1_98/A CLKBUF1_17/Y MUX2X1_85/Y gnd vdd DFFPOSX1
XOAI21X1_1261 OAI21X1_1260/Y AND2X2_55/Y BUFX4_32/Y gnd AOI21X1_511/C vdd OAI21X1
XOAI21X1_1250 OAI21X1_254/C BUFX4_244/Y AND2X2_33/B gnd OAI22X1_89/B vdd OAI21X1
XDFFPOSX1_873 NOR2X1_147/A CLKBUF1_32/Y AOI21X1_87/Y gnd vdd DFFPOSX1
XDFFPOSX1_862 NOR2X1_598/A CLKBUF1_32/Y AOI21X1_83/Y gnd vdd DFFPOSX1
XOAI21X1_1294 BUFX4_120/Y BUFX4_479/Y INVX1_350/A gnd OAI21X1_1294/Y vdd OAI21X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XDFFPOSX1_884 OAI21X1_194/C CLKBUF1_33/Y OAI21X1_195/Y gnd vdd DFFPOSX1
XINVX2_23 INVX2_23/A gnd INVX2_23/Y vdd INVX2
XDFFPOSX1_895 NOR2X1_159/A CLKBUF1_45/Y AOI21X1_95/Y gnd vdd DFFPOSX1
XFILL_4_7_1 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XFILL_29_7_1 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 BUFX4_450/Y BUFX4_293/Y INVX1_273/A gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XDFFPOSX1_103 NOR2X1_452/A CLKBUF1_91/Y AOI21X1_190/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 AND2X2_46/A CLKBUF1_100/Y OAI21X1_434/Y gnd vdd DFFPOSX1
XDFFPOSX1_125 NOR2X1_610/A CLKBUF1_100/Y OAI21X1_428/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 INVX1_180/A CLKBUF1_77/Y MUX2X1_166/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 INVX1_235/A CLKBUF1_41/Y MUX2X1_346/Y gnd vdd DFFPOSX1
XDFFPOSX1_147 NOR2X1_417/B CLKBUF1_24/Y DFFPOSX1_147/D gnd vdd DFFPOSX1
XDFFPOSX1_169 NOR2X1_545/A CLKBUF1_26/Y AOI21X1_569/Y gnd vdd DFFPOSX1
XNAND2X1_217 NOR2X1_164/A BUFX4_287/Y gnd NAND2X1_217/Y vdd NAND2X1
XNAND2X1_206 OAI21X1_429/C BUFX4_250/Y gnd OAI21X1_651/C vdd NAND2X1
XNAND2X1_239 BUFX4_289/Y NAND2X1_239/B gnd OAI21X1_774/C vdd NAND2X1
XNAND2X1_228 AND2X2_52/A NAND2X1_228/B gnd OAI21X1_724/C vdd NAND2X1
XBUFX4_190 INVX8_9/Y gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_250 BUFX4_308/Y BUFX4_136/Y gnd NOR2X1_733/B vdd NOR2X1
XNOR2X1_261 NOR2X1_261/A NOR2X1_261/B gnd NOR2X1_261/Y vdd NOR2X1
XNOR2X1_272 NOR2X1_272/A MUX2X1_410/S gnd NOR2X1_272/Y vdd NOR2X1
XNOR2X1_283 NOR2X1_283/A NOR2X1_30/B gnd NOR2X1_283/Y vdd NOR2X1
XNOR2X1_294 NOR2X1_294/A NOR2X1_47/B gnd NOR2X1_294/Y vdd NOR2X1
XOAI21X1_712 BUFX4_370/Y NOR2X1_97/A BUFX4_156/Y gnd OAI21X1_714/B vdd OAI21X1
XOAI21X1_701 BUFX4_334/Y NOR2X1_66/A BUFX4_157/Y gnd OAI22X1_17/C vdd OAI21X1
XOAI21X1_723 AOI22X1_18/Y NOR2X1_624/A OAI21X1_723/C gnd OAI21X1_723/Y vdd OAI21X1
XOAI21X1_734 BUFX4_257/Y INVX1_299/Y AOI21X1_322/Y gnd OAI21X1_734/Y vdd OAI21X1
XOAI21X1_745 OAI21X1_744/Y AOI21X1_327/Y BUFX4_169/Y gnd OAI21X1_745/Y vdd OAI21X1
XOAI21X1_767 BUFX4_329/Y NOR2X1_679/A AOI21X1_337/Y gnd OAI21X1_767/Y vdd OAI21X1
XOAI21X1_756 BUFX4_367/Y OAI21X1_756/B OAI21X1_756/C gnd OAI21X1_757/C vdd OAI21X1
XOAI21X1_789 OAI21X1_788/Y AND2X2_30/Y OAI21X1_787/Y gnd MUX2X1_215/B vdd OAI21X1
XOAI21X1_778 BUFX4_223/Y OAI21X1_778/B AOI21X1_340/Y gnd OAI21X1_778/Y vdd OAI21X1
XMUX2X1_223 MUX2X1_223/A MUX2X1_222/Y BUFX4_51/Y gnd MUX2X1_223/Y vdd MUX2X1
XMUX2X1_212 MUX2X1_212/A MUX2X1_212/B BUFX4_76/Y gnd MUX2X1_213/B vdd MUX2X1
XMUX2X1_201 MUX2X1_201/A MUX2X1_201/B BUFX4_88/Y gnd MUX2X1_203/B vdd MUX2X1
XOAI21X1_1091 AND2X2_29/A OAI21X1_1091/B BUFX4_88/Y gnd OAI22X1_49/B vdd OAI21X1
XMUX2X1_256 MUX2X1_256/A OAI22X1_49/Y BUFX4_41/Y gnd MUX2X1_256/Y vdd MUX2X1
XMUX2X1_234 MUX2X1_233/Y MUX2X1_234/B INVX8_30/A gnd MUX2X1_234/Y vdd MUX2X1
XOAI21X1_1080 INVX1_408/Y BUFX4_260/Y BUFX4_85/Y gnd AOI21X1_460/C vdd OAI21X1
XMUX2X1_245 NOR2X1_166/A MUX2X1_245/B INVX8_30/A gnd MUX2X1_245/Y vdd MUX2X1
XDFFPOSX1_670 NOR2X1_43/A CLKBUF1_4/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XMUX2X1_278 INVX1_447/Y BUFX4_317/Y MUX2X1_42/S gnd MUX2X1_278/Y vdd MUX2X1
XDFFPOSX1_692 INVX1_43/A CLKBUF1_94/Y MUX2X1_35/Y gnd vdd DFFPOSX1
XMUX2X1_267 BUFX4_421/Y INVX1_304/Y NOR2X1_54/Y gnd MUX2X1_267/Y vdd MUX2X1
XMUX2X1_289 BUFX4_318/Y INVX1_414/Y MUX2X1_50/S gnd MUX2X1_289/Y vdd MUX2X1
XDFFPOSX1_681 INVX1_39/A CLKBUF1_51/Y MUX2X1_31/Y gnd vdd DFFPOSX1
XFILL_44_5_1 gnd vdd FILL
XFILL_43_0_0 gnd vdd FILL
XBUFX4_41 BUFX4_33/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_52 BUFX4_54/A gnd BUFX4_52/Y vdd BUFX4
XBUFX4_30 BUFX4_28/A gnd BUFX4_30/Y vdd BUFX4
XBUFX4_74 BUFX4_11/Y gnd BUFX4_74/Y vdd BUFX4
XBUFX4_96 BUFX4_14/Y gnd BUFX4_96/Y vdd BUFX4
XBUFX4_63 INVX8_4/Y gnd BUFX4_63/Y vdd BUFX4
XBUFX4_85 BUFX4_85/A gnd BUFX4_85/Y vdd BUFX4
XFILL_34_0_0 gnd vdd FILL
XFILL_35_5_1 gnd vdd FILL
XOR2X2_4 traffic_Street_0[0] traffic_Street_0[1] gnd OR2X2_4/Y vdd OR2X2
XXNOR2X1_6 XOR2X1_3/A XNOR2X1_6/B gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_1_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_26_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX8_11 traffic_Street_1[0] gnd INVX8_11/Y vdd INVX8
XINVX8_33 INVX8_33/A gnd INVX8_33/Y vdd INVX8
XINVX8_22 INVX8_22/A gnd INVX8_22/Y vdd INVX8
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOAI21X1_520 OAI21X1_520/A NOR2X1_335/Y AOI22X1_7/Y gnd OAI21X1_520/Y vdd OAI21X1
XOAI21X1_531 INVX1_212/Y XNOR2X1_5/B NAND2X1_122/B gnd OAI21X1_531/Y vdd OAI21X1
XOAI21X1_553 BUFX4_342/Y NOR2X1_640/A AOI21X1_248/Y gnd NAND3X1_71/C vdd OAI21X1
XOAI21X1_542 INVX1_214/Y NOR3X1_10/Y OAI21X1_541/Y gnd AOI21X1_246/C vdd OAI21X1
XOAI21X1_564 INVX1_228/Y BUFX4_232/Y OAI21X1_564/C gnd MUX2X1_177/A vdd OAI21X1
XOAI21X1_575 INVX1_237/Y BUFX4_244/Y BUFX4_88/Y gnd AOI21X1_261/C vdd OAI21X1
XOAI21X1_586 OAI21X1_585/Y NOR2X1_372/Y BUFX4_39/Y gnd OAI22X1_5/A vdd OAI21X1
XOAI21X1_597 INVX1_256/Y BUFX4_266/Y BUFX4_97/Y gnd OAI21X1_598/B vdd OAI21X1
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_50_3_1 gnd vdd FILL
XFILL_41_3_1 gnd vdd FILL
XOAI21X1_350 INVX4_3/A BUFX4_199/Y OAI21X1_350/C gnd OAI21X1_351/C vdd OAI21X1
XOAI21X1_383 OAI21X1_11/A BUFX4_173/Y OAI21X1_382/Y gnd OAI21X1_383/Y vdd OAI21X1
XOAI21X1_361 MUX2X1_39/B NAND2X1_85/Y OAI21X1_361/C gnd DFFPOSX1_38/D vdd OAI21X1
XOAI21X1_372 BUFX4_209/Y NAND2X1_6/B NAND2X1_90/Y gnd DFFPOSX1_50/D vdd OAI21X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd NOR3X1_4/C vdd AND2X2
XOAI21X1_394 OAI21X1_24/A BUFX4_372/Y OAI21X1_393/Y gnd DFFPOSX1_92/D vdd OAI21X1
XINVX1_425 INVX1_425/A gnd INVX1_425/Y vdd INVX1
XINVX1_403 INVX1_403/A gnd INVX1_403/Y vdd INVX1
XINVX1_414 INVX1_414/A gnd INVX1_414/Y vdd INVX1
XINVX1_447 INVX1_447/A gnd INVX1_447/Y vdd INVX1
XINVX1_436 INVX1_436/A gnd INVX1_436/Y vdd INVX1
XINVX1_458 INVX1_458/A gnd INVX1_458/Y vdd INVX1
XFILL_49_4_1 gnd vdd FILL
XFILL_32_3_1 gnd vdd FILL
XAOI21X1_407 BUFX4_35/Y AOI21X1_407/B OAI21X1_936/Y gnd OAI22X1_39/B vdd AOI21X1
XAOI21X1_418 BUFX4_340/Y INVX1_381/Y AOI21X1_418/C gnd OAI21X1_962/A vdd AOI21X1
XAOI21X1_429 NAND2X1_363/A BUFX4_347/Y BUFX4_82/Y gnd OAI21X1_980/C vdd AOI21X1
XFILL_23_3_1 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XMUX2X1_18 INVX1_24/Y MUX2X1_18/B MUX2X1_18/S gnd MUX2X1_18/Y vdd MUX2X1
XMUX2X1_29 INVX1_37/Y MUX2X1_29/B MUX2X1_29/S gnd MUX2X1_29/Y vdd MUX2X1
XFILL_14_3_1 gnd vdd FILL
XAOI22X1_1 AND2X2_2/B AND2X2_2/A AOI22X1_1/C AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XOAI21X1_180 BUFX4_385/Y BUFX4_129/Y INVX1_393/A gnd OAI21X1_180/Y vdd OAI21X1
XOAI21X1_191 BUFX4_467/Y NAND2X1_58/Y OAI21X1_191/C gnd OAI21X1_191/Y vdd OAI21X1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XINVX1_266 INVX1_266/A gnd INVX1_266/Y vdd INVX1
XINVX1_277 INVX1_277/A gnd INVX1_277/Y vdd INVX1
XINVX1_299 INVX1_299/A gnd INVX1_299/Y vdd INVX1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XNAND2X1_11 NAND2X1_11/A OAI21X1_7/B gnd OAI21X1_6/C vdd NAND2X1
XNAND2X1_22 INVX8_5/A INVX4_4/Y gnd OAI21X1_24/A vdd NAND2X1
XNAND2X1_33 traffic_Street_1[1] NOR2X1_76/B gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_55 INVX8_19/A INVX8_9/A gnd MUX2X1_84/S vdd NAND2X1
XNAND2X1_77 INVX8_25/A INVX8_8/A gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_44 INVX8_18/A INVX8_6/A gnd NAND2X1_44/Y vdd NAND2X1
XNAND2X1_66 INVX8_22/A INVX4_5/Y gnd NAND2X1_66/Y vdd NAND2X1
XNAND2X1_99 MUX2X1_57/A NOR2X1_299/Y gnd NOR2X1_300/B vdd NAND2X1
XNAND2X1_88 NOR2X1_509/A NAND2X1_2/Y gnd NAND2X1_88/Y vdd NAND2X1
XNOR2X1_635 NOR2X1_635/A NOR2X1_65/Y gnd NOR2X1_635/Y vdd NOR2X1
XNOR2X1_602 NOR2X1_269/A BUFX4_333/Y gnd NOR2X1_602/Y vdd NOR2X1
XNOR2X1_624 NOR2X1_624/A OAI22X1_94/Y gnd NOR2X1_624/Y vdd NOR2X1
XNOR2X1_613 NOR2X1_613/A BUFX4_341/Y gnd NOR2X1_613/Y vdd NOR2X1
XNOR2X1_668 NOR2X1_668/A AOI21X1_72/B gnd NOR2X1_668/Y vdd NOR2X1
XNOR2X1_657 NOR2X1_657/A NOR2X1_107/B gnd NOR2X1_657/Y vdd NOR2X1
XNOR2X1_646 NOR2X1_646/A NOR2X1_92/B gnd NOR2X1_646/Y vdd NOR2X1
XFILL_35_2 gnd vdd FILL
XNOR2X1_679 NOR2X1_679/A MUX2X1_94/S gnd NOR2X1_679/Y vdd NOR2X1
XFILL_28_1 gnd vdd FILL
XAOI21X1_204 NAND3X1_5/B NAND3X1_5/C AND2X2_3/B gnd NAND2X1_106/B vdd AOI21X1
XAOI21X1_215 NAND2X1_117/Y AOI21X1_215/B AOI21X1_215/C gnd OR2X2_5/B vdd AOI21X1
XAOI21X1_237 AOI22X1_6/Y AOI21X1_237/B INVX1_207/Y gnd AOI21X1_237/Y vdd AOI21X1
XAOI21X1_226 AND2X2_9/Y OAI21X1_483/Y NOR3X1_13/B gnd NAND3X1_54/C vdd AOI21X1
XAOI21X1_248 BUFX4_342/Y INVX1_221/Y BUFX4_148/Y gnd AOI21X1_248/Y vdd AOI21X1
XAOI22X1_31 AOI22X1_31/A AOI22X1_31/B AOI22X1_31/C INVX8_33/A gnd AOI22X1_31/Y vdd
+ AOI22X1
XAOI21X1_259 BUFX4_48/Y AOI22X1_12/Y INVX8_33/A gnd AOI22X1_14/A vdd AOI21X1
XAOI22X1_20 AOI22X1_20/A AOI22X1_20/B BUFX4_168/Y AOI22X1_20/D gnd AOI22X1_20/Y vdd
+ AOI22X1
XOAI21X1_1421 NAND2X1_62/Y BUFX4_320/Y OAI21X1_1421/C gnd OAI21X1_1421/Y vdd OAI21X1
XOAI21X1_1410 BUFX4_449/Y BUFX4_404/Y NAND2X1_281/B gnd OAI21X1_1411/C vdd OAI21X1
XOAI21X1_1432 BUFX4_123/Y BUFX4_141/Y INVX1_306/A gnd OAI21X1_1432/Y vdd OAI21X1
XOAI21X1_1443 BUFX4_70/Y NAND2X1_68/Y OAI21X1_1442/Y gnd DFFPOSX1_284/D vdd OAI21X1
XOAI21X1_1465 BUFX4_451/Y BUFX4_162/Y INVX1_252/A gnd OAI21X1_1465/Y vdd OAI21X1
XOAI21X1_1454 INVX1_258/Y NOR2X1_188/B NAND2X1_358/Y gnd OAI21X1_1454/Y vdd OAI21X1
XOAI21X1_1498 NAND2X1_76/Y BUFX4_440/Y OAI21X1_1498/C gnd OAI21X1_1498/Y vdd OAI21X1
XOAI21X1_1476 BUFX4_429/Y NAND2X1_73/Y OAI21X1_1475/Y gnd OAI21X1_1476/Y vdd OAI21X1
XOAI21X1_1487 BUFX4_188/Y BUFX4_161/Y AND2X2_52/B gnd OAI21X1_1488/C vdd OAI21X1
XDFFPOSX1_1006 NOR2X1_621/A CLKBUF1_18/Y OAI21X1_295/Y gnd vdd DFFPOSX1
XDFFPOSX1_1017 NOR2X1_230/A CLKBUF1_67/Y AOI21X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_1028 INVX1_142/A CLKBUF1_34/Y MUX2X1_129/Y gnd vdd DFFPOSX1
XDFFPOSX1_1039 NOR2X1_241/A CLKBUF1_36/Y AOI21X1_152/Y gnd vdd DFFPOSX1
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B OAI22X1_4/C OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XFILL_46_2_1 gnd vdd FILL
XDFFPOSX1_307 INVX1_312/A CLKBUF1_56/Y DFFPOSX1_307/D gnd vdd DFFPOSX1
XDFFPOSX1_329 NOR2X1_539/B CLKBUF1_48/Y AOI21X1_551/Y gnd vdd DFFPOSX1
XDFFPOSX1_318 OAI21X1_590/B CLKBUF1_17/Y DFFPOSX1_318/D gnd vdd DFFPOSX1
XFILL_37_2_1 gnd vdd FILL
XBUFX4_372 INVX8_14/Y gnd BUFX4_372/Y vdd BUFX4
XBUFX4_361 BUFX4_29/Y gnd BUFX4_361/Y vdd BUFX4
XBUFX4_350 BUFX4_26/Y gnd BUFX4_350/Y vdd BUFX4
XNOR2X1_410 NOR2X1_410/A BUFX4_339/Y gnd OAI22X1_19/A vdd NOR2X1
XNOR2X1_443 NOR2X1_443/A BUFX4_247/Y gnd NOR2X1_443/Y vdd NOR2X1
XBUFX4_394 INVX8_28/Y gnd BUFX4_394/Y vdd BUFX4
XNOR2X1_432 NOR2X1_720/A BUFX4_155/Y gnd NOR2X1_432/Y vdd NOR2X1
XNOR2X1_421 BUFX4_277/Y NOR2X1_421/B gnd NOR2X1_421/Y vdd NOR2X1
XBUFX4_383 BUFX4_384/A gnd BUFX4_383/Y vdd BUFX4
XNOR2X1_465 INVX1_128/A BUFX4_340/Y gnd OAI22X1_33/A vdd NOR2X1
XNOR2X1_476 BUFX4_41/Y NOR2X1_475/Y gnd NOR2X1_476/Y vdd NOR2X1
XNOR2X1_454 NOR2X1_454/A BUFX4_350/Y gnd NOR2X1_454/Y vdd NOR2X1
XNOR2X1_487 BUFX4_34/Y NOR2X1_487/B gnd NOR2X1_487/Y vdd NOR2X1
XNOR2X1_498 AND2X2_23/A NOR2X1_498/B gnd NOR2X1_498/Y vdd NOR2X1
XOAI21X1_916 INVX1_348/Y BUFX4_253/Y BUFX4_88/Y gnd OAI21X1_916/Y vdd OAI21X1
XOAI21X1_905 NOR2X1_219/A BUFX4_244/Y BUFX4_84/Y gnd OAI22X1_35/B vdd OAI21X1
XOAI21X1_949 INVX1_373/Y BUFX4_276/Y NAND2X1_284/Y gnd MUX2X1_233/A vdd OAI21X1
XFILL_20_1_1 gnd vdd FILL
XOAI21X1_927 INVX1_357/Y BUFX4_96/Y BUFX4_353/Y gnd OAI21X1_928/A vdd OAI21X1
XOAI21X1_938 OAI21X1_937/Y NOR2X1_477/Y BUFX4_147/Y gnd OAI22X1_39/A vdd OAI21X1
XMUX2X1_405 INVX1_328/Y BUFX4_426/Y MUX2X1_406/S gnd MUX2X1_405/Y vdd MUX2X1
XOAI21X1_1240 BUFX4_364/Y NOR2X1_297/A BUFX4_149/Y gnd OAI22X1_85/C vdd OAI21X1
XOAI21X1_1251 BUFX4_344/Y NOR2X1_200/A BUFX4_151/Y gnd OAI22X1_90/C vdd OAI21X1
XDFFPOSX1_830 NOR2X1_593/A CLKBUF1_2/Y OAI21X1_167/Y gnd vdd DFFPOSX1
XDFFPOSX1_841 INVX1_99/A CLKBUF1_26/Y MUX2X1_86/Y gnd vdd DFFPOSX1
XOAI21X1_1273 BUFX4_448/Y BUFX4_43/Y INVX1_223/A gnd OAI21X1_1274/C vdd OAI21X1
XOAI21X1_1262 NOR2X1_623/Y AOI21X1_511/Y BUFX4_202/Y gnd NAND3X1_82/C vdd OAI21X1
XOAI21X1_1284 NAND2X1_32/Y BUFX4_421/Y OAI21X1_1283/Y gnd DFFPOSX1_143/D vdd OAI21X1
XDFFPOSX1_863 OAI21X1_184/C CLKBUF1_31/Y OAI21X1_185/Y gnd vdd DFFPOSX1
XDFFPOSX1_874 NOR2X1_599/A CLKBUF1_93/Y AOI21X1_88/Y gnd vdd DFFPOSX1
XOAI21X1_1295 NAND2X1_36/Y BUFX4_63/Y OAI21X1_1294/Y gnd OAI21X1_1295/Y vdd OAI21X1
XDFFPOSX1_852 NAND2X1_259/A CLKBUF1_85/Y OAI21X1_179/Y gnd vdd DFFPOSX1
XINVX2_24 INVX2_24/A gnd INVX2_24/Y vdd INVX2
XINVX2_13 BUFX2_3/A gnd INVX2_13/Y vdd INVX2
XDFFPOSX1_896 NOR2X1_160/A CLKBUF1_33/Y AOI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_885 INVX1_397/A CLKBUF1_12/Y OAI21X1_197/Y gnd vdd DFFPOSX1
XFILL_3_2_1 gnd vdd FILL
XFILL_28_2_1 gnd vdd FILL
XFILL_40_9_0 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XAOI21X1_590 BUFX4_420/Y NOR2X1_188/B NOR2X1_702/Y gnd AOI21X1_590/Y vdd AOI21X1
XFILL_19_2_1 gnd vdd FILL
XFILL_31_9_0 gnd vdd FILL
XDFFPOSX1_104 NOR2X1_288/A CLKBUF1_30/Y AOI21X1_191/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 INVX1_181/A CLKBUF1_4/Y MUX2X1_167/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 NOR2X1_294/A CLKBUF1_81/Y AOI21X1_197/Y gnd vdd DFFPOSX1
XDFFPOSX1_137 NOR2X1_611/A CLKBUF1_87/Y OAI21X1_436/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 NOR2X1_474/B CLKBUF1_28/Y DFFPOSX1_148/D gnd vdd DFFPOSX1
XDFFPOSX1_159 NOR2X1_693/A CLKBUF1_39/Y AOI21X1_581/Y gnd vdd DFFPOSX1
XNAND2X1_207 NOR2X1_251/A AND2X2_27/A gnd OAI21X1_655/C vdd NAND2X1
XNAND2X1_218 NOR2X1_154/A BUFX4_289/Y gnd NAND2X1_218/Y vdd NAND2X1
XNAND2X1_229 BUFX4_247/Y NOR2X1_647/A gnd OAI21X1_725/C vdd NAND2X1
XBUFX4_180 INVX8_13/Y gnd BUFX4_180/Y vdd BUFX4
XBUFX4_191 INVX8_9/Y gnd BUFX4_191/Y vdd BUFX4
XNOR2X1_251 NOR2X1_251/A NOR2X1_733/B gnd NOR2X1_251/Y vdd NOR2X1
XNOR2X1_240 BUFX4_311/Y BUFX4_56/Y gnd NOR2X1_727/B vdd NOR2X1
XNOR2X1_273 NOR2X1_273/A MUX2X1_410/S gnd NOR2X1_273/Y vdd NOR2X1
XNOR2X1_284 NOR2X1_284/A NOR2X1_30/B gnd NOR2X1_284/Y vdd NOR2X1
XNOR2X1_262 NOR2X1_262/A NOR2X1_261/B gnd NOR2X1_262/Y vdd NOR2X1
XFILL_22_9_0 gnd vdd FILL
XNOR2X1_295 NOR2X1_295/A NOR2X1_47/B gnd NOR2X1_295/Y vdd NOR2X1
XOAI21X1_713 INVX1_73/A BUFX4_362/Y OAI21X1_713/C gnd OAI21X1_714/C vdd OAI21X1
XOAI21X1_702 OAI21X1_83/C BUFX4_229/Y BUFX4_93/Y gnd OAI22X1_17/B vdd OAI21X1
XOAI21X1_724 INVX1_291/Y BUFX4_246/Y OAI21X1_724/C gnd MUX2X1_208/B vdd OAI21X1
XOAI21X1_735 INVX1_300/Y BUFX4_259/Y AND2X2_33/B gnd OAI21X1_736/A vdd OAI21X1
XOAI21X1_746 OAI21X1_746/A AOI21X1_328/Y BUFX4_390/Y gnd OAI21X1_746/Y vdd OAI21X1
XOAI21X1_757 NOR2X1_421/Y OAI21X1_757/B OAI21X1_757/C gnd OAI21X1_757/Y vdd OAI21X1
XOAI21X1_768 NOR2X1_427/Y OAI21X1_768/B OAI21X1_767/Y gnd OAI21X1_768/Y vdd OAI21X1
XOAI21X1_779 BUFX4_224/Y NOR2X1_714/A BUFX4_79/Y gnd OAI21X1_779/Y vdd OAI21X1
XMUX2X1_202 MUX2X1_202/A MUX2X1_202/B BUFX4_89/Y gnd MUX2X1_202/Y vdd MUX2X1
XMUX2X1_213 MUX2X1_213/A MUX2X1_213/B BUFX4_415/Y gnd MUX2X1_213/Y vdd MUX2X1
XOAI21X1_1081 BUFX4_32/Y OAI21X1_1078/Y NAND2X1_331/Y gnd OAI21X1_1081/Y vdd OAI21X1
XMUX2X1_224 MUX2X1_224/A MUX2X1_224/B BUFX4_116/Y gnd AND2X2_35/A vdd MUX2X1
XMUX2X1_235 MUX2X1_235/A MUX2X1_235/B BUFX4_37/Y gnd MUX2X1_235/Y vdd MUX2X1
XMUX2X1_246 MUX2X1_246/A MUX2X1_246/B BUFX4_410/Y gnd NOR2X1_498/B vdd MUX2X1
XOAI21X1_1070 AOI21X1_456/Y AOI21X1_457/Y BUFX4_33/Y gnd AND2X2_48/A vdd OAI21X1
XDFFPOSX1_671 INVX1_275/A CLKBUF1_96/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_660 OAI21X1_45/C CLKBUF1_88/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XMUX2X1_268 BUFX4_321/Y INVX1_412/Y NOR2X1_54/Y gnd MUX2X1_268/Y vdd MUX2X1
XDFFPOSX1_693 INVX1_44/A CLKBUF1_70/Y MUX2X1_36/Y gnd vdd DFFPOSX1
XOAI21X1_1092 INVX1_413/Y BUFX4_89/Y BUFX4_330/Y gnd AOI21X1_466/C vdd OAI21X1
XMUX2X1_257 MUX2X1_257/A MUX2X1_257/B BUFX4_112/Y gnd AND2X2_50/A vdd MUX2X1
XDFFPOSX1_682 INVX1_40/A CLKBUF1_100/Y MUX2X1_32/Y gnd vdd DFFPOSX1
XMUX2X1_279 BUFX4_445/Y INVX1_221/Y MUX2X1_45/S gnd MUX2X1_279/Y vdd MUX2X1
XFILL_43_0_1 gnd vdd FILL
XFILL_13_9_0 gnd vdd FILL
XBUFX4_20 address[0] gnd BUFX4_20/Y vdd BUFX4
XBUFX4_42 BUFX4_46/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_31 BUFX4_33/A gnd BUFX4_31/Y vdd BUFX4
XBUFX4_53 BUFX4_54/A gnd BUFX4_53/Y vdd BUFX4
XBUFX4_64 INVX8_4/Y gnd BUFX4_64/Y vdd BUFX4
XBUFX4_86 BUFX4_82/A gnd BUFX4_86/Y vdd BUFX4
XBUFX4_75 BUFX4_75/A gnd INVX8_32/A vdd BUFX4
XBUFX4_97 BUFX4_14/Y gnd BUFX4_97/Y vdd BUFX4
XFILL_34_0_1 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 XNOR2X1_7/A XNOR2X1_7/B gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX8_12 INVX8_12/A gnd BUFX4_46/A vdd INVX8
XINVX8_23 INVX8_23/A gnd INVX8_23/Y vdd INVX8
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XOAI21X1_510 NAND3X1_50/Y NOR2X1_334/B INVX1_208/Y gnd OAI21X1_510/Y vdd OAI21X1
XOAI21X1_521 XNOR2X1_4/B OR2X2_6/A AND2X2_10/Y gnd OAI21X1_522/C vdd OAI21X1
XOAI21X1_532 OR2X2_1/Y traffic_Street_1[0] traffic_Street_1[3] gnd NAND2X1_161/A vdd
+ OAI21X1
XOAI21X1_543 INVX4_12/Y INVX1_213/Y OAI21X1_497/A gnd INVX1_215/A vdd OAI21X1
XOAI21X1_554 BUFX4_352/Y NOR2X1_625/A BUFX4_157/Y gnd NOR2X1_364/B vdd OAI21X1
XOAI21X1_565 NOR2X1_366/Y NOR2X1_367/Y BUFX4_328/Y gnd OAI21X1_565/Y vdd OAI21X1
XOAI21X1_576 BUFX4_337/Y INVX1_239/Y BUFX4_151/Y gnd OAI21X1_577/A vdd OAI21X1
XOAI21X1_587 BUFX4_356/Y OAI21X1_587/B BUFX4_154/Y gnd AOI21X1_268/C vdd OAI21X1
XOAI21X1_598 NOR2X1_373/Y OAI21X1_598/B OAI21X1_598/C gnd MUX2X1_181/A vdd OAI21X1
XDFFPOSX1_490 INVX1_432/A CLKBUF1_65/Y MUX2X1_380/Y gnd vdd DFFPOSX1
XFILL_8_1_1 gnd vdd FILL
XFILL_45_8_0 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XFILL_36_8_0 gnd vdd FILL
XFILL_2_8_0 gnd vdd FILL
XFILL_27_8_0 gnd vdd FILL
XFILL_10_7_0 gnd vdd FILL
XOAI21X1_340 BUFX4_194/Y BUFX4_309/Y AND2X2_49/A gnd OAI21X1_340/Y vdd OAI21X1
XOAI21X1_351 NAND2X1_82/Y MUX2X1_83/B OAI21X1_351/C gnd OAI21X1_351/Y vdd OAI21X1
XOAI21X1_362 BUFX4_188/Y BUFX4_197/Y INVX1_339/A gnd OAI21X1_362/Y vdd OAI21X1
XOAI21X1_373 BUFX4_178/Y NAND2X1_6/B NAND2X1_91/Y gnd DFFPOSX1_51/D vdd OAI21X1
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_395 BUFX4_450/Y BUFX4_293/Y NOR2X1_606/A gnd OAI21X1_395/Y vdd OAI21X1
XOAI21X1_384 BUFX4_294/Y BUFX4_299/Y NOR2X1_503/A gnd OAI21X1_384/Y vdd OAI21X1
XINVX1_404 INVX1_404/A gnd INVX1_404/Y vdd INVX1
XINVX1_426 INVX1_426/A gnd INVX1_426/Y vdd INVX1
XINVX1_415 INVX1_415/A gnd INVX1_415/Y vdd INVX1
XINVX1_459 INVX1_459/A gnd INVX1_459/Y vdd INVX1
XINVX1_437 INVX1_437/A gnd INVX1_437/Y vdd INVX1
XINVX1_448 INVX1_448/A gnd INVX1_448/Y vdd INVX1
XFILL_18_8_0 gnd vdd FILL
XAOI21X1_419 BUFX4_285/Y INVX1_382/Y AOI21X1_419/C gnd OAI21X1_962/B vdd AOI21X1
XAOI21X1_408 BUFX4_35/Y NOR2X1_648/A OAI21X1_939/Y gnd OAI22X1_39/C vdd AOI21X1
XMUX2X1_19 INVX1_25/Y BUFX4_71/Y MUX2X1_18/S gnd MUX2X1_19/Y vdd MUX2X1
XFILL_42_6_0 gnd vdd FILL
XAOI22X1_2 traffic_Street_1[3] OR2X2_1/Y AOI22X1_2/C AOI22X1_2/D gnd AOI22X1_2/Y vdd
+ AOI22X1
XOAI21X1_181 NAND2X1_57/Y MUX2X1_82/B OAI21X1_180/Y gnd OAI21X1_181/Y vdd OAI21X1
XOAI21X1_170 BUFX4_128/Y BUFX4_297/Y INVX1_337/A gnd OAI21X1_171/C vdd OAI21X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XOAI21X1_192 BUFX4_387/Y BUFX4_408/Y INVX1_287/A gnd OAI21X1_192/Y vdd OAI21X1
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XINVX1_212 AOI22X1_7/C gnd INVX1_212/Y vdd INVX1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XINVX1_267 INVX1_267/A gnd INVX1_267/Y vdd INVX1
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XINVX1_256 INVX1_256/A gnd INVX1_256/Y vdd INVX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XNAND2X1_34 traffic_Street_1[3] NOR2X1_76/B gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_12 INVX1_330/A OAI21X1_7/B gnd OAI21X1_7/C vdd NAND2X1
XNAND2X1_23 NOR2X1_4/Y NOR2X1_12/Y gnd BUFX4_124/A vdd NAND2X1
XNAND2X1_56 INVX8_20/A INVX4_2/Y gnd NAND2X1_56/Y vdd NAND2X1
XNAND2X1_45 INVX8_18/A INVX4_3/Y gnd MUX2X1_71/S vdd NAND2X1
XNAND2X1_67 INVX8_23/A INVX4_2/Y gnd MUX2X1_360/S vdd NAND2X1
XNAND2X1_89 NAND2X1_89/A NAND2X1_2/Y gnd NAND2X1_89/Y vdd NAND2X1
XNAND2X1_78 INVX8_26/A INVX4_2/Y gnd NAND2X1_78/Y vdd NAND2X1
XNOR2X1_603 BUFX4_231/Y INVX1_166/Y gnd NOR2X1_603/Y vdd NOR2X1
XNOR2X1_625 NOR2X1_625/A NOR2X1_54/Y gnd NOR2X1_625/Y vdd NOR2X1
XNOR2X1_614 BUFX4_413/Y NOR2X1_614/B gnd OAI22X1_91/B vdd NOR2X1
XNOR2X1_669 NOR2X1_669/A AOI21X1_72/B gnd NOR2X1_669/Y vdd NOR2X1
XNOR2X1_636 NOR2X1_523/A NOR2X1_70/Y gnd NOR2X1_636/Y vdd NOR2X1
XNOR2X1_658 AND2X2_22/B AOI21X1_62/B gnd NOR2X1_658/Y vdd NOR2X1
XNOR2X1_647 NOR2X1_647/A NOR2X1_92/B gnd NOR2X1_647/Y vdd NOR2X1
XFILL_35_3 gnd vdd FILL
XFILL_33_6_0 gnd vdd FILL
XAOI21X1_216 NAND3X1_27/Y OAI21X1_468/Y NOR3X1_3/B gnd AOI21X1_219/B vdd AOI21X1
XAOI21X1_205 NAND3X1_6/C NAND3X1_28/C INVX4_8/Y gnd NOR3X1_2/B vdd AOI21X1
XAOI21X1_238 INVX1_207/A AOI21X1_238/B OAI21X1_510/Y gnd NAND3X1_65/C vdd AOI21X1
XAOI21X1_227 NAND3X1_64/C NOR2X1_327/Y AOI21X1_227/C gnd OAI21X1_492/A vdd AOI21X1
XAOI21X1_249 BUFX4_76/Y OAI21X1_555/Y NOR2X1_364/Y gnd AOI21X1_249/Y vdd AOI21X1
XAOI22X1_21 AOI22X1_21/A AOI22X1_21/B AOI22X1_21/C BUFX4_205/Y gnd AOI22X1_21/Y vdd
+ AOI22X1
XAOI22X1_32 BUFX4_166/Y AOI22X1_32/B AND2X2_48/Y AOI22X1_32/D gnd OAI22X1_48/B vdd
+ AOI22X1
XAOI22X1_10 INVX1_214/Y NOR3X1_10/Y AOI22X1_9/C AOI22X1_10/D gnd AOI22X1_10/Y vdd
+ AOI22X1
XOAI21X1_1411 NAND2X1_61/Y BUFX4_73/Y OAI21X1_1411/C gnd DFFPOSX1_176/D vdd OAI21X1
XOAI21X1_1400 BUFX4_143/Y BUFX4_403/Y OAI21X1_756/B gnd OAI21X1_1401/C vdd OAI21X1
XOAI21X1_1422 BUFX4_383/Y BUFX4_141/Y INVX1_234/A gnd OAI21X1_1423/C vdd OAI21X1
XOAI21X1_1444 BUFX4_61/Y BUFX4_433/Y OAI21X1_1153/B gnd OAI21X1_1444/Y vdd OAI21X1
XOAI21X1_1466 NAND2X1_72/Y BUFX4_445/Y OAI21X1_1465/Y gnd OAI21X1_1466/Y vdd OAI21X1
XOAI21X1_1455 INVX1_380/Y NOR2X1_188/B NAND2X1_359/Y gnd DFFPOSX1_445/D vdd OAI21X1
XOAI21X1_1433 NAND2X1_66/Y BUFX4_420/Y OAI21X1_1432/Y gnd OAI21X1_1433/Y vdd OAI21X1
XOAI21X1_1499 BUFX4_389/Y BUFX4_458/Y NOR2X1_434/A gnd OAI21X1_1500/C vdd OAI21X1
XOAI21X1_1477 BUFX4_135/Y BUFX4_160/Y AOI21X1_414/B gnd OAI21X1_1478/C vdd OAI21X1
XOAI21X1_1488 BUFX4_324/Y NAND2X1_74/Y OAI21X1_1488/C gnd DFFPOSX1_494/D vdd OAI21X1
XFILL_24_6_0 gnd vdd FILL
XDFFPOSX1_1007 NOR2X1_223/A CLKBUF1_60/Y AOI21X1_140/Y gnd vdd DFFPOSX1
XDFFPOSX1_1018 NOR2X1_231/A CLKBUF1_89/Y AOI21X1_147/Y gnd vdd DFFPOSX1
XDFFPOSX1_1029 INVX1_143/A CLKBUF1_52/Y MUX2X1_130/Y gnd vdd DFFPOSX1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B OAI22X1_5/C BUFX4_39/Y gnd OAI22X1_5/Y vdd OAI22X1
XFILL_7_7_0 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XDFFPOSX1_308 INVX1_372/A CLKBUF1_56/Y DFFPOSX1_308/D gnd vdd DFFPOSX1
XDFFPOSX1_319 OAI21X1_760/B CLKBUF1_16/Y OAI21X1_1353/Y gnd vdd DFFPOSX1
XBUFX4_340 BUFX4_25/Y gnd BUFX4_340/Y vdd BUFX4
XBUFX4_362 BUFX4_25/Y gnd BUFX4_362/Y vdd BUFX4
XNOR2X1_400 NOR2X1_400/A BUFX4_226/Y gnd OAI22X1_16/D vdd NOR2X1
XBUFX4_351 BUFX4_29/Y gnd BUFX4_351/Y vdd BUFX4
XBUFX4_373 INVX8_14/Y gnd MUX2X1_61/B vdd BUFX4
XFILL_40_1 gnd vdd FILL
XNOR2X1_422 BUFX4_278/Y NOR2X1_422/B gnd NOR2X1_422/Y vdd NOR2X1
XBUFX4_395 INVX8_18/Y gnd BUFX4_395/Y vdd BUFX4
XNOR2X1_433 BUFX4_81/Y NOR2X1_716/A gnd NOR2X1_433/Y vdd NOR2X1
XNOR2X1_411 NOR2X1_411/A NOR2X1_411/B gnd NOR2X1_411/Y vdd NOR2X1
XBUFX4_384 BUFX4_384/A gnd BUFX4_384/Y vdd BUFX4
XNOR2X1_444 OAI21X1_77/C BUFX4_250/Y gnd NOR2X1_445/A vdd NOR2X1
XNOR2X1_455 NAND2X1_87/A BUFX4_222/Y gnd NOR2X1_455/Y vdd NOR2X1
XNOR2X1_477 BUFX4_413/Y INVX1_364/Y gnd NOR2X1_477/Y vdd NOR2X1
XNOR2X1_466 NOR2X1_466/A BUFX4_241/Y gnd OAI22X1_34/D vdd NOR2X1
XNOR2X1_499 NOR2X1_499/A AND2X2_25/B gnd NOR2X1_500/A vdd NOR2X1
XNOR2X1_488 BUFX4_206/Y NOR2X1_487/Y gnd NOR2X1_488/Y vdd NOR2X1
XOAI21X1_906 OAI22X1_35/Y BUFX4_38/Y BUFX4_202/Y gnd OAI22X1_36/D vdd OAI21X1
XOAI21X1_917 NOR2X1_471/Y OAI21X1_916/Y OAI21X1_915/Y gnd NAND2X1_277/B vdd OAI21X1
XOAI21X1_928 OAI21X1_928/A AND2X2_39/Y BUFX4_38/Y gnd OAI22X1_38/A vdd OAI21X1
XOAI21X1_939 BUFX4_35/Y INVX1_366/Y AND2X2_29/A gnd OAI21X1_939/Y vdd OAI21X1
XOAI21X1_1230 INVX1_162/Y BUFX4_332/Y AOI21X1_505/Y gnd NAND3X1_81/B vdd OAI21X1
XOAI21X1_1252 OAI21X1_262/C BUFX4_246/Y BUFX4_108/Y gnd OAI22X1_90/B vdd OAI21X1
XDFFPOSX1_842 INVX1_100/A CLKBUF1_62/Y MUX2X1_87/Y gnd vdd DFFPOSX1
XOAI21X1_1274 NAND2X1_31/Y BUFX4_442/Y OAI21X1_1274/C gnd OAI21X1_1274/Y vdd OAI21X1
XDFFPOSX1_831 NOR2X1_394/A CLKBUF1_75/Y AOI21X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_820 AND2X2_34/B CLKBUF1_75/Y OAI21X1_155/Y gnd vdd DFFPOSX1
XMUX2X1_406 INVX1_460/Y BUFX4_63/Y MUX2X1_406/S gnd MUX2X1_406/Y vdd MUX2X1
XOAI21X1_1263 BUFX4_48/Y OAI22X1_91/Y NAND3X1_82/Y gnd OAI22X1_93/B vdd OAI21X1
XOAI21X1_1241 NOR2X1_298/A AND2X2_51/B BUFX4_104/Y gnd OAI22X1_85/B vdd OAI21X1
XDFFPOSX1_875 INVX1_108/A CLKBUF1_41/Y MUX2X1_95/Y gnd vdd DFFPOSX1
XOAI21X1_1285 BUFX4_124/Y BUFX4_46/Y OAI21X1_933/B gnd OAI21X1_1285/Y vdd OAI21X1
XDFFPOSX1_853 INVX1_393/A CLKBUF1_31/Y OAI21X1_181/Y gnd vdd DFFPOSX1
XDFFPOSX1_864 NAND2X1_257/A CLKBUF1_5/Y OAI21X1_187/Y gnd vdd DFFPOSX1
XOAI21X1_1296 INVX4_5/A NOR2X1_74/B AOI21X1_466/B gnd OAI21X1_1297/C vdd OAI21X1
XINVX2_25 INVX2_25/A gnd INVX2_25/Y vdd INVX2
XDFFPOSX1_897 MUX2X1_247/A CLKBUF1_71/Y AOI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_886 OAI21X1_198/C CLKBUF1_12/Y OAI21X1_199/Y gnd vdd DFFPOSX1
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XFILL_40_9_1 gnd vdd FILL
XAOI21X1_580 BUFX4_320/Y NOR2X1_167/B NOR2X1_692/Y gnd AOI21X1_580/Y vdd AOI21X1
XAOI21X1_591 BUFX4_444/Y NOR2X1_703/B NOR2X1_703/Y gnd AOI21X1_591/Y vdd AOI21X1
XFILL_47_5_0 gnd vdd FILL
XFILL_31_9_1 gnd vdd FILL
XFILL_30_4_0 gnd vdd FILL
XDFFPOSX1_105 NOR2X1_289/A CLKBUF1_40/Y AOI21X1_192/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NOR2X1_295/A CLKBUF1_6/Y AOI21X1_198/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 INVX1_182/A CLKBUF1_46/Y MUX2X1_168/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 NOR2X1_522/B CLKBUF1_28/Y DFFPOSX1_149/D gnd vdd DFFPOSX1
XDFFPOSX1_138 NOR2X1_400/A CLKBUF1_43/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XNAND2X1_208 DFFPOSX1_6/Q BUFX4_256/Y gnd OAI21X1_656/C vdd NAND2X1
XNAND2X1_219 NAND2X1_219/A BUFX4_291/Y gnd NAND2X1_219/Y vdd NAND2X1
XFILL_38_5_0 gnd vdd FILL
XBUFX4_170 INVX8_29/Y gnd BUFX4_170/Y vdd BUFX4
XBUFX4_181 INVX8_13/Y gnd MUX2X1_64/B vdd BUFX4
XNOR2X1_252 NOR2X1_252/A NOR2X1_733/B gnd NOR2X1_252/Y vdd NOR2X1
XNOR2X1_241 NOR2X1_241/A NOR2X1_727/B gnd NOR2X1_241/Y vdd NOR2X1
XBUFX4_192 INVX8_9/Y gnd BUFX4_192/Y vdd BUFX4
XNOR2X1_230 NOR2X1_230/A NOR2X1_231/B gnd NOR2X1_230/Y vdd NOR2X1
XNOR2X1_274 NOR2X1_274/A MUX2X1_410/S gnd NOR2X1_274/Y vdd NOR2X1
XNOR2X1_263 NOR2X1_263/A NOR2X1_261/B gnd NOR2X1_263/Y vdd NOR2X1
XNOR2X1_285 NOR2X1_285/A NOR2X1_30/B gnd NOR2X1_285/Y vdd NOR2X1
XFILL_22_9_1 gnd vdd FILL
XNOR2X1_296 NOR2X1_296/A NOR2X1_47/B gnd NOR2X1_296/Y vdd NOR2X1
XOAI21X1_714 NOR2X1_408/Y OAI21X1_714/B OAI21X1_714/C gnd OAI21X1_715/A vdd OAI21X1
XOAI21X1_703 OAI22X1_17/Y BUFX4_41/Y BUFX4_169/Y gnd NOR2X1_405/B vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XOAI21X1_736 OAI21X1_736/A AND2X2_28/Y OAI21X1_734/Y gnd OAI21X1_736/Y vdd OAI21X1
XOAI21X1_747 BUFX4_392/Y AOI22X1_19/Y OAI21X1_746/Y gnd AOI21X1_339/B vdd OAI21X1
XOAI21X1_725 INVX1_292/Y BUFX4_248/Y OAI21X1_725/C gnd MUX2X1_208/A vdd OAI21X1
XOAI21X1_758 BUFX4_40/Y AOI21X1_334/Y OAI21X1_758/C gnd AOI22X1_20/D vdd OAI21X1
XOAI21X1_769 OAI21X1_768/Y BUFX4_39/Y BUFX4_207/Y gnd OAI21X1_769/Y vdd OAI21X1
XMUX2X1_214 MUX2X1_214/A MUX2X1_214/B BUFX4_80/Y gnd MUX2X1_214/Y vdd MUX2X1
XMUX2X1_203 MUX2X1_202/Y MUX2X1_203/B BUFX4_40/Y gnd MUX2X1_203/Y vdd MUX2X1
XOAI21X1_1060 BUFX4_348/Y NOR2X1_199/A BUFX4_147/Y gnd NOR2X1_512/B vdd OAI21X1
XDFFPOSX1_650 OAI21X1_33/C CLKBUF1_103/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XMUX2X1_236 MUX2X1_236/A MUX2X1_236/B BUFX4_118/Y gnd MUX2X1_236/Y vdd MUX2X1
XMUX2X1_225 MUX2X1_225/A MUX2X1_225/B INVX8_32/A gnd MUX2X1_225/Y vdd MUX2X1
XOAI21X1_1071 INVX1_139/Y BUFX4_250/Y NAND2X1_329/Y gnd MUX2X1_254/B vdd OAI21X1
XOAI21X1_1082 OAI21X1_1081/Y BUFX4_170/Y BUFX4_49/Y gnd OAI22X1_48/C vdd OAI21X1
XMUX2X1_247 MUX2X1_247/A MUX2X1_247/B BUFX4_411/Y gnd MUX2X1_247/Y vdd MUX2X1
XDFFPOSX1_661 OAI21X1_47/C CLKBUF1_88/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XMUX2X1_269 BUFX4_442/Y INVX1_222/Y NOR2X1_57/Y gnd MUX2X1_269/Y vdd MUX2X1
XOAI21X1_1093 INVX1_414/Y BUFX4_91/Y BUFX4_268/Y gnd AOI21X1_467/C vdd OAI21X1
XDFFPOSX1_683 OAI21X1_59/C CLKBUF1_81/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_672 NOR2X1_440/A CLKBUF1_51/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XMUX2X1_258 MUX2X1_258/A MUX2X1_258/B BUFX4_38/Y gnd MUX2X1_258/Y vdd MUX2X1
XDFFPOSX1_694 NOR2X1_59/A CLKBUF1_70/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XFILL_4_5_0 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_13_9_1 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XINVX8_1 traffic_Street_0[3] gnd INVX8_1/Y vdd INVX8
XBUFX4_10 clock gnd BUFX4_10/Y vdd BUFX4
XBUFX4_43 BUFX4_46/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 address[0] gnd BUFX4_21/Y vdd BUFX4
XBUFX4_32 BUFX4_33/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_65 INVX8_4/Y gnd BUFX4_65/Y vdd BUFX4
XBUFX4_76 BUFX4_11/Y gnd BUFX4_76/Y vdd BUFX4
XBUFX4_87 BUFX4_87/A gnd BUFX4_87/Y vdd BUFX4
XBUFX4_54 BUFX4_54/A gnd BUFX4_54/Y vdd BUFX4
XBUFX4_98 BUFX4_14/Y gnd BUFX4_98/Y vdd BUFX4
XFILL_10_2 gnd vdd FILL
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XXNOR2X1_8 XNOR2X1_8/A INVX2_4/A gnd XNOR2X1_8/Y vdd XNOR2X1
XINVX8_13 traffic_Street_1[1] gnd INVX8_13/Y vdd INVX8
XINVX8_24 INVX8_24/A gnd INVX8_24/Y vdd INVX8
XOAI21X1_500 BUFX4_306/Y INVX4_11/Y AND2X2_10/Y gnd OAI21X1_500/Y vdd OAI21X1
XOAI21X1_522 NOR2X1_331/Y OR2X2_6/Y OAI21X1_522/C gnd NAND3X1_58/B vdd OAI21X1
XOAI21X1_511 AOI21X1_237/Y OAI21X1_510/Y AOI22X1_5/D gnd NAND3X1_51/C vdd OAI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XOAI21X1_533 AOI22X1_9/D AOI22X1_9/C NOR2X1_347/Y gnd NAND3X1_66/A vdd OAI21X1
XOAI21X1_544 NOR2X1_357/B INVX1_217/Y INVX1_218/A gnd NAND2X1_167/A vdd OAI21X1
XOAI21X1_555 INVX1_222/Y BUFX4_224/Y NAND2X1_170/Y gnd OAI21X1_555/Y vdd OAI21X1
XOAI21X1_566 BUFX4_328/Y OAI21X1_566/B OAI21X1_565/Y gnd AOI21X1_255/B vdd OAI21X1
XOAI21X1_599 BUFX4_369/Y OAI21X1_599/B BUFX4_147/Y gnd AOI21X1_275/C vdd OAI21X1
XOAI21X1_577 OAI21X1_577/A NOR2X1_369/Y BUFX4_414/Y gnd OAI22X1_4/C vdd OAI21X1
XOAI21X1_588 INVX1_247/Y BUFX4_253/Y NAND2X1_176/Y gnd OAI21X1_588/Y vdd OAI21X1
XDFFPOSX1_491 AND2X2_23/B CLKBUF1_54/Y OAI21X1_1482/Y gnd vdd DFFPOSX1
XDFFPOSX1_480 OAI21X1_778/B CLKBUF1_44/Y DFFPOSX1_480/D gnd vdd DFFPOSX1
XFILL_45_8_1 gnd vdd FILL
XFILL_44_3_0 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_36_8_1 gnd vdd FILL
XFILL_2_8_1 gnd vdd FILL
XFILL_27_8_1 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_10_7_1 gnd vdd FILL
XOAI21X1_341 MUX2X1_86/B NAND2X1_81/Y OAI21X1_340/Y gnd DFFPOSX1_8/D vdd OAI21X1
XOAI21X1_330 NOR2X1_84/B BUFX4_308/Y INVX1_340/A gnd OAI21X1_330/Y vdd OAI21X1
XOAI21X1_363 MUX2X1_40/B NAND2X1_85/Y OAI21X1_362/Y gnd OAI21X1_363/Y vdd OAI21X1
XOAI21X1_374 BUFX4_375/Y NAND2X1_6/B NAND2X1_92/Y gnd DFFPOSX1_52/D vdd OAI21X1
XOAI21X1_352 INVX4_5/A BUFX4_197/Y INVX1_276/A gnd OAI21X1_353/C vdd OAI21X1
XINVX1_416 INVX1_416/A gnd INVX1_416/Y vdd INVX1
XOAI21X1_396 OAI21X1_24/A BUFX4_470/Y OAI21X1_395/Y gnd DFFPOSX1_93/D vdd OAI21X1
XOAI21X1_385 OAI21X1_11/A BUFX4_375/Y OAI21X1_384/Y gnd DFFPOSX1_76/D vdd OAI21X1
XINVX1_405 INVX1_405/A gnd INVX1_405/Y vdd INVX1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XINVX1_427 INVX1_427/A gnd INVX1_427/Y vdd INVX1
XINVX1_449 INVX1_449/A gnd INVX1_449/Y vdd INVX1
XINVX1_438 INVX1_438/A gnd INVX1_438/Y vdd INVX1
XFILL_9_4_0 gnd vdd FILL
XFILL_18_8_1 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XAOI21X1_409 BUFX4_51/Y OAI22X1_39/Y INVX8_33/A gnd AOI22X1_25/D vdd AOI21X1
XFILL_50_1_0 gnd vdd FILL
XFILL_41_1_0 gnd vdd FILL
XFILL_42_6_1 gnd vdd FILL
XAOI22X1_3 AND2X2_5/B AND2X2_5/A AOI22X1_3/C AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_171 NAND2X1_56/Y MUX2X1_49/A OAI21X1_171/C gnd OAI21X1_171/Y vdd OAI21X1
XOAI21X1_182 INVX4_3/A BUFX4_128/Y OAI21X1_182/C gnd OAI21X1_183/C vdd OAI21X1
XOAI21X1_160 BUFX4_454/Y BUFX4_186/Y OAI21X1_160/C gnd OAI21X1_161/C vdd OAI21X1
XINVX1_235 INVX1_235/A gnd INVX1_235/Y vdd INVX1
XINVX1_202 OAI22X1_2/D gnd INVX1_202/Y vdd INVX1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XOAI21X1_193 NAND2X1_59/Y AND2X2_2/B OAI21X1_192/Y gnd OAI21X1_193/Y vdd OAI21X1
XINVX1_213 OAI22X1_3/A gnd INVX1_213/Y vdd INVX1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XFILL_49_2_0 gnd vdd FILL
XNAND2X1_24 INVX8_5/A INVX4_5/Y gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_13 NAND2X1_13/A OAI21X1_7/B gnd OAI21X1_8/C vdd NAND2X1
XNAND2X1_57 INVX8_20/A INVX4_3/Y gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_46 INVX8_18/A INVX4_4/Y gnd MUX2X1_76/S vdd NAND2X1
XNAND2X1_35 INVX8_16/A INVX8_6/A gnd MUX2X1_42/S vdd NAND2X1
XNAND2X1_68 INVX8_23/A INVX8_6/A gnd NAND2X1_68/Y vdd NAND2X1
XNAND2X1_79 INVX8_26/A INVX4_3/Y gnd NAND2X1_79/Y vdd NAND2X1
XNOR2X1_604 NOR2X1_604/A BUFX4_232/Y gnd NOR2X1_604/Y vdd NOR2X1
XNOR2X1_626 NOR2X1_626/A NOR2X1_54/Y gnd NOR2X1_626/Y vdd NOR2X1
XNOR2X1_615 NOR2X1_615/A BUFX4_241/Y gnd NOR2X1_615/Y vdd NOR2X1
XNOR2X1_637 NOR2X1_637/A NOR2X1_76/B gnd NOR2X1_637/Y vdd NOR2X1
XNOR2X1_659 AND2X2_27/B AOI21X1_62/B gnd NOR2X1_659/Y vdd NOR2X1
XNOR2X1_648 NOR2X1_648/A NOR2X1_92/B gnd NOR2X1_648/Y vdd NOR2X1
XFILL_32_1_0 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XAOI21X1_206 MUX2X1_57/A NAND3X1_5/B AND2X2_3/B gnd NOR3X1_1/B vdd AOI21X1
XAOI21X1_228 NAND3X1_46/Y OAI21X1_500/Y NOR3X1_12/B gnd AOI21X1_231/B vdd AOI21X1
XAOI21X1_239 AOI21X1_236/Y NAND3X1_56/Y NOR2X1_334/A gnd OAI21X1_515/A vdd AOI21X1
XAOI21X1_217 NAND3X1_12/B OR2X2_2/Y INVX2_14/Y gnd NOR3X1_8/A vdd AOI21X1
XAOI22X1_11 AOI22X1_11/A AOI22X1_11/B AOI22X1_11/C BUFX4_167/Y gnd AOI22X1_11/Y vdd
+ AOI22X1
XAOI22X1_33 AOI22X1_33/A AOI22X1_33/B OAI22X1_42/Y INVX4_13/Y gnd AOI22X1_33/Y vdd
+ AOI22X1
XAOI22X1_22 AOI22X1_22/A BUFX4_168/Y AOI22X1_22/C AOI22X1_22/D gnd MUX2X1_223/A vdd
+ AOI22X1
XOAI21X1_1401 BUFX4_422/Y NAND2X1_60/Y OAI21X1_1401/C gnd OAI21X1_1401/Y vdd OAI21X1
XOAI21X1_1412 BUFX4_452/Y BUFX4_403/Y NOR2X1_536/B gnd OAI21X1_1413/C vdd OAI21X1
XOAI21X1_1423 NAND2X1_64/Y BUFX4_437/Y OAI21X1_1423/C gnd DFFPOSX1_210/D vdd OAI21X1
XOAI21X1_1445 MUX2X1_29/B NAND2X1_68/Y OAI21X1_1444/Y gnd OAI21X1_1445/Y vdd OAI21X1
XNOR3X1_1 INVX4_8/A NOR3X1_1/B AND2X2_3/Y gnd NOR3X1_2/A vdd NOR3X1
XOAI21X1_1434 BUFX4_123/Y BUFX4_140/Y AND2X2_40/B gnd OAI21X1_1435/C vdd OAI21X1
XOAI21X1_1456 INVX1_428/Y NOR2X1_188/B NAND2X1_360/Y gnd OAI21X1_1456/Y vdd OAI21X1
XOAI21X1_1489 BUFX4_456/Y BUFX4_298/Y INVX1_264/A gnd OAI21X1_1489/Y vdd OAI21X1
XOAI21X1_1478 BUFX4_72/Y NAND2X1_73/Y OAI21X1_1478/C gnd DFFPOSX1_485/D vdd OAI21X1
XOAI21X1_1467 BUFX4_451/Y BUFX4_164/Y OAI21X1_778/B gnd OAI21X1_1468/C vdd OAI21X1
XFILL_24_6_1 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XDFFPOSX1_1008 NOR2X1_224/A CLKBUF1_89/Y AOI21X1_141/Y gnd vdd DFFPOSX1
XDFFPOSX1_1019 INVX1_137/A CLKBUF1_16/Y MUX2X1_124/Y gnd vdd DFFPOSX1
XOAI22X1_6 OAI22X1_6/A OAI22X1_6/B OAI22X1_6/C OAI22X1_6/D gnd OAI22X1_6/Y vdd OAI22X1
XFILL_7_7_1 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_309 NOR2X1_542/B CLKBUF1_2/Y DFFPOSX1_309/D gnd vdd DFFPOSX1
XBUFX4_330 BUFX4_29/Y gnd BUFX4_330/Y vdd BUFX4
XBUFX4_341 BUFX4_25/Y gnd BUFX4_341/Y vdd BUFX4
XBUFX4_363 BUFX4_28/Y gnd BUFX4_363/Y vdd BUFX4
XBUFX4_352 BUFX4_28/Y gnd BUFX4_352/Y vdd BUFX4
XNOR2X1_401 NOR2X1_61/A BUFX4_352/Y gnd NOR2X1_401/Y vdd NOR2X1
XBUFX4_385 BUFX4_384/A gnd BUFX4_385/Y vdd BUFX4
XNOR2X1_423 NOR2X1_423/A BUFX4_327/Y gnd NOR2X1_423/Y vdd NOR2X1
XNOR2X1_434 NOR2X1_434/A BUFX4_155/Y gnd NOR2X1_434/Y vdd NOR2X1
XBUFX4_374 INVX8_14/Y gnd MUX2X1_57/A vdd BUFX4
XBUFX4_396 INVX8_18/Y gnd BUFX4_396/Y vdd BUFX4
XNOR2X1_412 BUFX4_100/Y NOR2X1_412/B gnd NOR2X1_412/Y vdd NOR2X1
XFILL_40_2 gnd vdd FILL
XNOR2X1_467 NOR2X1_467/A BUFX4_362/Y gnd OAI22X1_34/A vdd NOR2X1
XNOR2X1_445 NOR2X1_445/A NOR2X1_445/B gnd NOR2X1_445/Y vdd NOR2X1
XNOR2X1_456 INVX1_160/A BUFX4_347/Y gnd NOR2X1_456/Y vdd NOR2X1
XFILL_33_1 gnd vdd FILL
XNOR2X1_478 BUFX4_414/Y INVX1_367/Y gnd NOR2X1_478/Y vdd NOR2X1
XNOR2X1_489 BUFX4_235/Y INVX1_16/Y gnd NOR2X1_489/Y vdd NOR2X1
XOAI21X1_907 OAI21X1_907/A OAI21X1_907/B address[6] gnd OAI21X1_907/Y vdd OAI21X1
XOAI21X1_918 BUFX4_255/Y INVX1_349/Y AOI21X1_395/Y gnd OAI21X1_918/Y vdd OAI21X1
XOAI21X1_929 INVX1_358/Y BUFX4_97/Y AND2X2_23/A gnd AOI21X1_402/C vdd OAI21X1
XOAI21X1_1220 OAI22X1_79/Y BUFX4_39/Y BUFX4_201/Y gnd OAI22X1_80/A vdd OAI21X1
XOAI21X1_1231 INVX1_158/Y BUFX4_346/Y AOI21X1_506/Y gnd NAND3X1_81/C vdd OAI21X1
XMUX2X1_407 INVX1_461/Y MUX2X1_4/B MUX2X1_406/S gnd MUX2X1_407/Y vdd MUX2X1
XDFFPOSX1_832 NOR2X1_127/A CLKBUF1_23/Y AOI21X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_821 INVX1_395/A CLKBUF1_17/Y OAI21X1_157/Y gnd vdd DFFPOSX1
XOAI21X1_1264 OAI22X1_93/Y INVX4_14/Y street gnd OAI22X1_94/B vdd OAI21X1
XOAI21X1_1242 OAI22X1_85/Y BUFX4_31/Y BUFX4_205/Y gnd OAI22X1_86/D vdd OAI21X1
XOAI21X1_1253 BUFX4_357/Y NOR2X1_226/A BUFX4_155/Y gnd OAI22X1_92/C vdd OAI21X1
XDFFPOSX1_810 NOR2X1_582/A CLKBUF1_77/Y AOI21X1_65/Y gnd vdd DFFPOSX1
XOAI21X1_1286 NAND2X1_32/Y BUFX4_64/Y OAI21X1_1285/Y gnd OAI21X1_1286/Y vdd OAI21X1
XDFFPOSX1_843 NOR2X1_396/A CLKBUF1_31/Y OAI21X1_169/Y gnd vdd DFFPOSX1
XOAI21X1_1275 BUFX4_448/Y BUFX4_45/Y NOR2X1_417/B gnd OAI21X1_1275/Y vdd OAI21X1
XDFFPOSX1_865 NAND2X1_301/A CLKBUF1_32/Y OAI21X1_189/Y gnd vdd DFFPOSX1
XDFFPOSX1_854 OAI21X1_182/C CLKBUF1_5/Y OAI21X1_183/Y gnd vdd DFFPOSX1
XOAI21X1_1297 NAND2X1_36/Y BUFX4_318/Y OAI21X1_1297/C gnd OAI21X1_1297/Y vdd OAI21X1
XDFFPOSX1_876 INVX1_109/A CLKBUF1_59/Y MUX2X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_898 NOR2X1_162/A CLKBUF1_101/Y AOI21X1_98/Y gnd vdd DFFPOSX1
XINVX2_26 INVX2_26/A gnd INVX2_26/Y vdd INVX2
XDFFPOSX1_887 NAND2X1_219/A CLKBUF1_7/Y OAI21X1_201/Y gnd vdd DFFPOSX1
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XAOI21X1_570 BUFX4_422/Y MUX2X1_96/S NOR2X1_682/Y gnd AOI21X1_570/Y vdd AOI21X1
XAOI21X1_581 BUFX4_430/Y NOR2X1_172/B NOR2X1_693/Y gnd AOI21X1_581/Y vdd AOI21X1
XAOI21X1_592 MUX2X1_27/B NOR2X1_703/B NOR2X1_704/Y gnd AOI21X1_592/Y vdd AOI21X1
XFILL_47_5_1 gnd vdd FILL
XFILL_46_0_0 gnd vdd FILL
XFILL_30_4_1 gnd vdd FILL
XDFFPOSX1_117 INVX1_183/A CLKBUF1_95/Y MUX2X1_169/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 NOR2X1_296/A CLKBUF1_99/Y AOI21X1_199/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 NOR2X1_379/A CLKBUF1_77/Y OAI21X1_406/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 INVX1_332/A CLKBUF1_43/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XNAND2X1_209 BUFX4_32/Y OAI22X1_9/Y gnd NAND2X1_209/Y vdd NAND2X1
XFILL_37_0_0 gnd vdd FILL
XFILL_38_5_1 gnd vdd FILL
XBUFX4_171 INVX8_29/Y gnd BUFX4_171/Y vdd BUFX4
XBUFX4_182 INVX8_13/Y gnd MUX2X1_77/B vdd BUFX4
XBUFX4_160 INVX8_24/Y gnd BUFX4_160/Y vdd BUFX4
XBUFX4_193 INVX8_9/Y gnd BUFX4_193/Y vdd BUFX4
XNOR2X1_242 AND2X2_37/A NOR2X1_727/B gnd NOR2X1_242/Y vdd NOR2X1
XNOR2X1_231 NOR2X1_231/A NOR2X1_231/B gnd NOR2X1_231/Y vdd NOR2X1
XNOR2X1_220 NOR2X1_220/A NOR2X1_220/B gnd NOR2X1_220/Y vdd NOR2X1
XNOR2X1_275 NOR2X1_275/A NOR2X1_16/Y gnd NOR2X1_275/Y vdd NOR2X1
XNOR2X1_253 NOR2X1_253/A NOR2X1_733/B gnd NOR2X1_253/Y vdd NOR2X1
XNOR2X1_264 NOR2X1_264/A NOR2X1_261/B gnd NOR2X1_264/Y vdd NOR2X1
XNOR2X1_286 NOR2X1_286/A NOR2X1_33/Y gnd NOR2X1_286/Y vdd NOR2X1
XNOR2X1_297 NOR2X1_297/A NOR2X1_47/B gnd NOR2X1_297/Y vdd NOR2X1
XOAI21X1_704 INVX1_56/Y BUFX4_231/Y NAND2X1_222/Y gnd MUX2X1_205/B vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XOAI21X1_715 OAI21X1_715/A BUFX4_33/Y BUFX4_166/Y gnd AOI21X1_313/C vdd OAI21X1
XOAI21X1_737 INVX1_301/Y BUFX4_260/Y BUFX4_152/Y gnd OAI21X1_737/Y vdd OAI21X1
XOAI21X1_726 NOR2X1_413/Y NOR2X1_414/Y BUFX4_358/Y gnd OAI21X1_727/C vdd OAI21X1
XOAI21X1_748 BUFX4_266/Y INVX1_305/Y AOI21X1_329/Y gnd OAI21X1_748/Y vdd OAI21X1
XOAI21X1_759 BUFX4_327/Y OAI21X1_759/B BUFX4_153/Y gnd OAI22X1_20/C vdd OAI21X1
XMUX2X1_204 MUX2X1_204/A MUX2X1_204/B BUFX4_90/Y gnd MUX2X1_204/Y vdd MUX2X1
XOAI21X1_1061 INVX1_129/Y BUFX4_359/Y NAND2X1_326/Y gnd AOI21X1_454/B vdd OAI21X1
XMUX2X1_226 MUX2X1_226/A MUX2X1_226/B BUFX4_77/Y gnd MUX2X1_226/Y vdd MUX2X1
XOAI21X1_1072 INVX1_143/Y BUFX4_252/Y NAND2X1_330/Y gnd MUX2X1_254/A vdd OAI21X1
XOAI21X1_1050 BUFX4_360/Y INVX1_157/A BUFX4_149/Y gnd NOR2X1_510/B vdd OAI21X1
XDFFPOSX1_640 NOR2X1_443/A CLKBUF1_66/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XMUX2X1_215 MUX2X1_215/A MUX2X1_215/B BUFX4_32/Y gnd MUX2X1_216/B vdd MUX2X1
XMUX2X1_237 MUX2X1_237/A MUX2X1_237/B BUFX4_76/Y gnd MUX2X1_237/Y vdd MUX2X1
XMUX2X1_259 MUX2X1_259/A MUX2X1_259/B INVX8_32/A gnd MUX2X1_259/Y vdd MUX2X1
XDFFPOSX1_651 NOR2X1_34/A CLKBUF1_30/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XOAI21X1_1094 AOI21X1_466/Y AOI21X1_467/Y BUFX4_412/Y gnd NAND2X1_332/B vdd OAI21X1
XOAI21X1_1083 INVX2_2/Y read_Write BUFX2_7/A gnd OAI21X1_1084/C vdd OAI21X1
XDFFPOSX1_684 OAI21X1_61/C CLKBUF1_96/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_673 INVX1_392/A CLKBUF1_96/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XMUX2X1_248 MUX2X1_248/A MUX2X1_248/B AND2X2_33/B gnd MUX2X1_248/Y vdd MUX2X1
XDFFPOSX1_662 AND2X2_51/A CLKBUF1_1/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_695 NOR2X1_61/A CLKBUF1_24/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XFILL_4_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_29_5_1 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_12_4_1 gnd vdd FILL
XINVX8_2 traffic_Street_0[0] gnd INVX8_2/Y vdd INVX8
XBUFX4_11 address[1] gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 BUFX4_46/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_22 address[0] gnd BUFX4_22/Y vdd BUFX4
XBUFX4_33 BUFX4_33/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_77 BUFX4_11/Y gnd BUFX4_77/Y vdd BUFX4
XBUFX4_66 INVX8_4/Y gnd BUFX4_66/Y vdd BUFX4
XBUFX4_55 BUFX4_54/A gnd BUFX4_55/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_88 BUFX4_11/Y gnd BUFX4_88/Y vdd BUFX4
XBUFX4_99 BUFX4_75/A gnd BUFX4_99/Y vdd BUFX4
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XXNOR2X1_9 INVX8_9/A INVX4_1/Y gnd XNOR2X1_9/Y vdd XNOR2X1
XINVX8_25 INVX8_25/A gnd INVX8_25/Y vdd INVX8
XINVX8_14 traffic_Street_1[2] gnd INVX8_14/Y vdd INVX8
XOAI21X1_512 AOI21X1_237/Y OAI21X1_510/Y AND2X2_8/A gnd NAND3X1_53/C vdd OAI21X1
XOAI21X1_523 AOI21X1_237/Y OAI21X1_510/Y XOR2X1_3/A gnd NAND3X1_59/C vdd OAI21X1
XOAI21X1_501 INVX1_187/A AOI22X1_1/Y INVX2_24/A gnd NAND2X1_144/A vdd OAI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XOAI21X1_534 BUFX4_305/Y OAI22X1_2/D OR2X2_2/A gnd OAI21X1_534/Y vdd OAI21X1
XOAI21X1_556 BUFX4_349/Y NOR2X1_632/A BUFX4_159/Y gnd AOI21X1_250/C vdd OAI21X1
XOAI21X1_545 OR2X2_7/A OR2X2_7/B NOR2X1_356/Y gnd OAI21X1_545/Y vdd OAI21X1
XOAI21X1_589 INVX1_248/Y BUFX4_255/Y OAI21X1_589/C gnd OAI21X1_589/Y vdd OAI21X1
XOAI21X1_567 INVX1_230/Y BUFX4_234/Y NAND2X1_175/Y gnd OAI21X1_567/Y vdd OAI21X1
XOAI21X1_578 BUFX4_148/Y OAI21X1_578/B BUFX4_367/Y gnd NOR2X1_371/B vdd OAI21X1
XDFFPOSX1_481 INVX1_374/A CLKBUF1_7/Y OAI21X1_1470/Y gnd vdd DFFPOSX1
XDFFPOSX1_492 NOR2X1_431/A CLKBUF1_44/Y DFFPOSX1_492/D gnd vdd DFFPOSX1
XDFFPOSX1_470 INVX1_433/A CLKBUF1_22/Y MUX2X1_371/Y gnd vdd DFFPOSX1
XFILL_44_3_1 gnd vdd FILL
XFILL_35_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XOAI21X1_331 NAND2X1_80/Y BUFX4_180/Y OAI21X1_330/Y gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_320 BUFX4_389/Y BUFX4_313/Y OAI21X1_320/C gnd OAI21X1_321/C vdd OAI21X1
XOAI21X1_342 BUFX4_194/Y BUFX4_309/Y DFFPOSX1_9/Q gnd OAI21X1_343/C vdd OAI21X1
XOAI21X1_364 BUFX4_191/Y BUFX4_198/Y NAND2X1_325/A gnd OAI21X1_365/C vdd OAI21X1
XOAI21X1_353 NAND2X1_84/Y MUX2X1_39/B OAI21X1_353/C gnd DFFPOSX1_34/D vdd OAI21X1
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XINVX1_406 INVX1_406/A gnd INVX1_406/Y vdd INVX1
XOAI21X1_375 BUFX4_468/Y NAND2X1_6/B NAND2X1_93/Y gnd DFFPOSX1_53/D vdd OAI21X1
XOAI21X1_386 BUFX4_295/Y BUFX4_299/Y NOR2X1_604/A gnd OAI21X1_387/C vdd OAI21X1
XOAI21X1_397 BUFX4_125/Y BUFX4_292/Y INVX1_279/A gnd OAI21X1_397/Y vdd OAI21X1
XINVX1_417 INVX1_417/A gnd INVX1_417/Y vdd INVX1
XINVX1_439 INVX1_439/A gnd INVX1_439/Y vdd INVX1
XINVX1_428 INVX1_428/A gnd INVX1_428/Y vdd INVX1
XFILL_9_4_1 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XFILL_50_1_1 gnd vdd FILL
XFILL_41_1_1 gnd vdd FILL
XAOI22X1_4 NOR3X1_9/Y INVX2_22/Y NOR3X1_10/Y INVX2_21/Y gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_172 BUFX4_130/Y BUFX4_297/Y INVX1_394/A gnd OAI21X1_173/C vdd OAI21X1
XOAI21X1_183 NAND2X1_57/Y MUX2X1_83/B OAI21X1_183/C gnd OAI21X1_183/Y vdd OAI21X1
XOAI21X1_161 NAND2X1_53/Y BUFX4_217/Y OAI21X1_161/C gnd OAI21X1_161/Y vdd OAI21X1
XOAI21X1_150 BUFX4_59/Y BUFX4_183/Y OAI21X1_150/C gnd OAI21X1_151/C vdd OAI21X1
XINVX1_203 INVX1_203/A gnd INVX1_203/Y vdd INVX1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XOAI21X1_194 BUFX4_387/Y BUFX4_407/Y OAI21X1_194/C gnd OAI21X1_194/Y vdd OAI21X1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XINVX1_258 INVX1_258/A gnd INVX1_258/Y vdd INVX1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XNAND2X1_14 NAND2X1_14/A OAI21X1_7/B gnd OAI21X1_9/C vdd NAND2X1
XNAND2X1_25 INVX8_10/A INVX4_2/Y gnd OAI21X1_40/A vdd NAND2X1
XFILL_49_2_1 gnd vdd FILL
XNAND2X1_58 INVX8_20/A INVX8_8/A gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_36 INVX8_16/A INVX4_5/Y gnd NAND2X1_36/Y vdd NAND2X1
XNAND2X1_47 traffic_Street_1[1] NOR2X1_107/B gnd NAND2X1_47/Y vdd NAND2X1
XNAND2X1_69 INVX8_23/A INVX4_3/Y gnd NAND2X1_69/Y vdd NAND2X1
XNOR2X1_605 NOR2X1_281/A BUFX4_343/Y gnd NOR2X1_605/Y vdd NOR2X1
XNOR2X1_616 NOR2X1_616/A BUFX4_345/Y gnd NOR2X1_616/Y vdd NOR2X1
XNOR2X1_627 NOR2X1_627/A NOR2X1_57/Y gnd NOR2X1_627/Y vdd NOR2X1
XNOR2X1_638 NOR2X1_638/A NOR2X1_76/B gnd NOR2X1_638/Y vdd NOR2X1
XNOR2X1_649 NOR2X1_528/A NOR2X1_92/B gnd NOR2X1_649/Y vdd NOR2X1
XFILL_32_1_1 gnd vdd FILL
XAOI21X1_207 NAND3X1_14/B OR2X2_4/Y INVX2_15/A gnd AOI21X1_207/Y vdd AOI21X1
XAOI21X1_229 INVX4_7/Y NOR3X1_7/Y INVX2_24/Y gnd OAI21X1_502/B vdd AOI21X1
XAOI21X1_218 NAND3X1_10/Y NAND3X1_11/C INVX2_14/A gnd NOR3X1_8/B vdd AOI21X1
XAOI22X1_23 BUFX4_400/Y MUX2X1_223/Y AOI22X1_23/C AOI22X1_23/D gnd AOI22X1_23/Y vdd
+ AOI22X1
XAOI22X1_12 BUFX4_202/Y AOI22X1_12/B AOI22X1_12/C AOI22X1_12/D gnd AOI22X1_12/Y vdd
+ AOI22X1
XOAI21X1_1402 BUFX4_142/Y BUFX4_405/Y MUX2X1_231/B gnd OAI21X1_1402/Y vdd OAI21X1
XOAI21X1_1413 NAND2X1_61/Y BUFX4_320/Y OAI21X1_1413/C gnd OAI21X1_1413/Y vdd OAI21X1
XOAI21X1_1446 BUFX4_384/Y BUFX4_434/Y OAI21X1_600/B gnd OAI21X1_1446/Y vdd OAI21X1
XOAI21X1_1435 NAND2X1_66/Y BUFX4_66/Y OAI21X1_1435/C gnd DFFPOSX1_264/D vdd OAI21X1
XOAI21X1_1424 BUFX4_383/Y BUFX4_140/Y OAI21X1_752/B gnd OAI21X1_1425/C vdd OAI21X1
XOAI21X1_1457 BUFX4_126/Y BUFX4_431/Y OAI21X1_603/B gnd OAI21X1_1457/Y vdd OAI21X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XOAI21X1_1479 BUFX4_135/Y BUFX4_160/Y AOI21X1_487/B gnd OAI21X1_1479/Y vdd OAI21X1
XOAI21X1_1468 NAND2X1_72/Y BUFX4_422/Y OAI21X1_1468/C gnd DFFPOSX1_480/D vdd OAI21X1
XFILL_23_1_1 gnd vdd FILL
XDFFPOSX1_1009 NOR2X1_516/A CLKBUF1_67/Y AOI21X1_142/Y gnd vdd DFFPOSX1
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_43_9_0 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XBUFX4_331 BUFX4_27/Y gnd BUFX4_331/Y vdd BUFX4
XBUFX4_320 INVX8_1/Y gnd BUFX4_320/Y vdd BUFX4
XBUFX4_342 BUFX4_30/Y gnd BUFX4_342/Y vdd BUFX4
XBUFX4_364 BUFX4_26/Y gnd BUFX4_364/Y vdd BUFX4
XBUFX4_353 BUFX4_26/Y gnd BUFX4_353/Y vdd BUFX4
XNOR2X1_402 BUFX4_415/Y OAI22X1_16/Y gnd NOR2X1_405/A vdd NOR2X1
XNOR2X1_424 BUFX4_284/Y NOR2X1_424/B gnd NOR2X1_424/Y vdd NOR2X1
XBUFX4_375 INVX8_14/Y gnd BUFX4_375/Y vdd BUFX4
XBUFX4_386 BUFX4_384/A gnd BUFX4_386/Y vdd BUFX4
XNOR2X1_413 INVX1_450/A BUFX4_158/Y gnd NOR2X1_413/Y vdd NOR2X1
XBUFX4_397 INVX8_18/Y gnd BUFX4_397/Y vdd BUFX4
XFILL_40_3 gnd vdd FILL
XNOR2X1_457 BUFX4_229/Y INVX1_341/Y gnd NOR2X1_457/Y vdd NOR2X1
XNOR2X1_435 BUFX4_82/Y NOR2X1_435/B gnd NOR2X1_435/Y vdd NOR2X1
XNOR2X1_446 INVX1_53/Y BUFX4_152/Y gnd NOR2X1_446/Y vdd NOR2X1
XNOR2X1_468 INVX8_30/A NOR2X1_468/B gnd OAI22X1_36/C vdd NOR2X1
XFILL_34_9_0 gnd vdd FILL
XFILL_26_1 gnd vdd FILL
XNOR2X1_479 BUFX4_268/Y NOR2X1_479/B gnd NOR2X1_479/Y vdd NOR2X1
XOAI21X1_919 INVX1_350/Y BUFX4_257/Y BUFX4_90/Y gnd OAI21X1_920/A vdd OAI21X1
XOAI21X1_908 address[6] AOI22X1_23/Y OAI21X1_907/Y gnd OAI21X1_908/Y vdd OAI21X1
XOAI21X1_1221 OAI22X1_80/Y BUFX4_51/Y BUFX4_402/Y gnd OAI22X1_81/B vdd OAI21X1
XOAI21X1_1210 INVX1_442/Y BUFX4_288/Y BUFX4_93/Y gnd AOI21X1_500/C vdd OAI21X1
XOAI21X1_1265 BUFX4_301/Y BUFX4_45/Y NOR2X1_363/A gnd OAI21X1_1265/Y vdd OAI21X1
XMUX2X1_408 BUFX4_441/Y INVX1_271/Y MUX2X1_410/S gnd MUX2X1_408/Y vdd MUX2X1
XDFFPOSX1_833 NOR2X1_128/A CLKBUF1_90/Y AOI21X1_74/Y gnd vdd DFFPOSX1
XOAI21X1_1232 AOI21X1_504/Y OAI21X1_1229/Y NAND3X1_81/Y gnd AOI21X1_507/B vdd OAI21X1
XDFFPOSX1_822 OAI21X1_158/C CLKBUF1_75/Y OAI21X1_159/Y gnd vdd DFFPOSX1
XOAI21X1_1243 OAI22X1_86/Y BUFX4_392/Y INVX8_33/A gnd OAI22X1_93/D vdd OAI21X1
XOAI21X1_1254 OAI21X1_302/C BUFX4_248/Y BUFX4_109/Y gnd OAI22X1_92/B vdd OAI21X1
XDFFPOSX1_811 NOR2X1_118/A CLKBUF1_89/Y AOI21X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_800 INVX1_90/A CLKBUF1_15/Y OAI21X1_133/Y gnd vdd DFFPOSX1
XOAI21X1_1287 BUFX4_124/Y BUFX4_44/Y OAI21X1_1091/B gnd OAI21X1_1287/Y vdd OAI21X1
XOAI21X1_1276 NAND2X1_31/Y BUFX4_421/Y OAI21X1_1275/Y gnd DFFPOSX1_147/D vdd OAI21X1
XDFFPOSX1_866 OAI21X1_190/C CLKBUF1_32/Y OAI21X1_191/Y gnd vdd DFFPOSX1
XDFFPOSX1_855 NOR2X1_397/A CLKBUF1_69/Y AOI21X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_844 INVX1_337/A CLKBUF1_5/Y OAI21X1_171/Y gnd vdd DFFPOSX1
XOAI21X1_1298 BUFX4_189/Y BUFX4_478/Y AND2X2_21/B gnd OAI21X1_1299/C vdd OAI21X1
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XDFFPOSX1_899 INVX1_286/A CLKBUF1_101/Y OAI21X1_217/Y gnd vdd DFFPOSX1
XDFFPOSX1_877 MUX2X1_246/B CLKBUF1_12/Y AOI21X1_89/Y gnd vdd DFFPOSX1
XDFFPOSX1_888 INVX1_335/A CLKBUF1_8/Y OAI21X1_203/Y gnd vdd DFFPOSX1
XFILL_0_9_0 gnd vdd FILL
XFILL_25_9_0 gnd vdd FILL
XAOI21X1_560 BUFX4_426/Y NOR2X1_137/B NOR2X1_672/Y gnd AOI21X1_560/Y vdd AOI21X1
XAOI21X1_571 BUFX4_320/Y MUX2X1_96/S NOR2X1_683/Y gnd AOI21X1_571/Y vdd AOI21X1
XAOI21X1_593 BUFX4_68/Y NOR2X1_703/B NOR2X1_705/Y gnd AOI21X1_593/Y vdd AOI21X1
XAOI21X1_582 BUFX4_437/Y MUX2X1_102/S NOR2X1_694/Y gnd AOI21X1_582/Y vdd AOI21X1
XFILL_46_0_1 gnd vdd FILL
XFILL_16_9_0 gnd vdd FILL
XDFFPOSX1_107 AOI21X1_382/A CLKBUF1_88/Y OAI21X1_408/Y gnd vdd DFFPOSX1
XDFFPOSX1_118 NOR2X1_290/A CLKBUF1_88/Y AOI21X1_193/Y gnd vdd DFFPOSX1
XCLKBUF1_1 BUFX4_10/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_129 NOR2X1_297/A CLKBUF1_96/Y AOI21X1_200/Y gnd vdd DFFPOSX1
XBUFX4_150 INVX8_32/Y gnd BUFX4_150/Y vdd BUFX4
XBUFX4_161 INVX8_24/Y gnd BUFX4_161/Y vdd BUFX4
XFILL_37_0_1 gnd vdd FILL
XBUFX4_172 INVX8_13/Y gnd MUX2X1_96/A vdd BUFX4
XBUFX4_194 INVX8_9/Y gnd BUFX4_194/Y vdd BUFX4
XBUFX4_183 INVX8_19/Y gnd BUFX4_183/Y vdd BUFX4
XNOR2X1_232 BUFX4_459/Y BUFX4_451/Y gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_243 NOR2X1_243/A NOR2X1_727/B gnd NOR2X1_243/Y vdd NOR2X1
XNOR2X1_221 INVX2_7/Y INVX2_12/Y gnd INVX8_25/A vdd NOR2X1
XNOR2X1_210 BUFX4_161/Y BUFX4_384/Y gnd MUX2X1_120/S vdd NOR2X1
XNOR2X1_276 NOR2X1_276/A NOR2X1_16/Y gnd NOR2X1_276/Y vdd NOR2X1
XNOR2X1_254 DFFPOSX1_1/Q NOR2X1_733/B gnd NOR2X1_254/Y vdd NOR2X1
XNOR2X1_265 BUFX4_198/Y BUFX4_144/Y gnd NOR2X1_737/B vdd NOR2X1
XNOR2X1_287 NOR2X1_452/A NOR2X1_33/Y gnd NOR2X1_287/Y vdd NOR2X1
XNOR2X1_298 NOR2X1_298/A MUX2X1_31/S gnd NOR2X1_298/Y vdd NOR2X1
XOAI21X1_705 INVX1_289/Y BUFX4_233/Y OAI21X1_705/C gnd MUX2X1_205/A vdd OAI21X1
XOAI21X1_738 INVX1_302/Y BUFX4_262/Y BUFX4_108/Y gnd AOI21X1_324/C vdd OAI21X1
XOAI21X1_727 BUFX4_353/Y AOI21X1_318/Y OAI21X1_727/C gnd MUX2X1_209/A vdd OAI21X1
XOAI21X1_716 BUFX4_338/Y NOR2X1_107/A BUFX4_158/Y gnd OAI21X1_716/Y vdd OAI21X1
XOAI21X1_749 INVX1_306/Y BUFX4_268/Y BUFX4_114/Y gnd OAI21X1_750/A vdd OAI21X1
XOAI21X1_1040 BUFX4_349/Y NOR2X1_284/A BUFX4_159/Y gnd OAI22X1_45/C vdd OAI21X1
XMUX2X1_205 MUX2X1_205/A MUX2X1_205/B BUFX4_94/Y gnd MUX2X1_205/Y vdd MUX2X1
XOAI21X1_1062 BUFX4_348/Y OAI21X1_244/C BUFX4_147/Y gnd OAI22X1_47/C vdd OAI21X1
XMUX2X1_227 MUX2X1_227/A MUX2X1_227/B BUFX4_79/Y gnd MUX2X1_227/Y vdd MUX2X1
XMUX2X1_238 MUX2X1_238/A MUX2X1_238/B BUFX4_77/Y gnd MUX2X1_238/Y vdd MUX2X1
XDFFPOSX1_630 NOR2X1_20/A CLKBUF1_21/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_641 NOR2X1_492/A CLKBUF1_66/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XOAI21X1_1051 NAND2X1_92/A BUFX4_226/Y BUFX4_116/Y gnd AOI21X1_451/C vdd OAI21X1
XMUX2X1_216 MUX2X1_216/A MUX2X1_216/B BUFX4_165/Y gnd MUX2X1_216/Y vdd MUX2X1
XOAI21X1_1073 NOR2X1_515/Y NOR2X1_516/Y BUFX4_253/Y gnd NAND3X1_80/B vdd OAI21X1
XDFFPOSX1_652 INVX1_33/A CLKBUF1_30/Y MUX2X1_25/Y gnd vdd DFFPOSX1
XOAI21X1_1084 AOI22X1_33/Y NOR2X1_624/A OAI21X1_1084/C gnd OAI21X1_1084/Y vdd OAI21X1
XDFFPOSX1_674 INVX1_426/A CLKBUF1_87/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XMUX2X1_249 MUX2X1_249/A MUX2X1_249/B BUFX4_110/Y gnd MUX2X1_249/Y vdd MUX2X1
XDFFPOSX1_663 INVX1_34/A CLKBUF1_58/Y MUX2X1_26/Y gnd vdd DFFPOSX1
XOAI21X1_1095 BUFX4_270/Y INVX1_453/A AOI21X1_468/Y gnd OAI21X1_1095/Y vdd OAI21X1
XDFFPOSX1_696 NOR2X1_62/A CLKBUF1_43/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_685 OAI21X1_63/C CLKBUF1_100/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XFILL_3_0_1 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XINVX8_3 traffic_Street_0[1] gnd INVX8_3/Y vdd INVX8
XFILL_40_7_0 gnd vdd FILL
XAOI21X1_390 BUFX4_38/Y OAI22X1_31/Y BUFX4_201/Y gnd OAI21X1_896/C vdd AOI21X1
XBUFX4_34 BUFX4_33/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_23 address[0] gnd BUFX4_23/Y vdd BUFX4
XBUFX4_12 address[1] gnd BUFX4_87/A vdd BUFX4
XFILL_48_8_0 gnd vdd FILL
XBUFX4_67 INVX8_4/Y gnd BUFX4_67/Y vdd BUFX4
XBUFX4_45 BUFX4_46/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_56 INVX8_6/Y gnd BUFX4_56/Y vdd BUFX4
XBUFX4_78 BUFX4_11/Y gnd BUFX4_78/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_89 BUFX4_11/Y gnd BUFX4_89/Y vdd BUFX4
XFILL_31_7_0 gnd vdd FILL
XFILL_39_8_0 gnd vdd FILL
XINVX8_15 traffic_Street_1[3] gnd INVX8_15/Y vdd INVX8
XINVX8_26 INVX8_26/A gnd INVX8_26/Y vdd INVX8
XFILL_22_7_0 gnd vdd FILL
XOAI21X1_502 AOI21X1_230/Y OAI21X1_502/B OAI21X1_502/C gnd NAND3X1_56/C vdd OAI21X1
XOAI21X1_513 NOR2X1_336/B INVX4_10/A AND2X2_8/A gnd NAND3X1_55/C vdd OAI21X1
XOAI21X1_535 BUFX4_305/Y INVX4_11/Y XNOR2X1_6/B gnd OAI21X1_536/C vdd OAI21X1
XOAI21X1_524 NOR2X1_336/B INVX4_10/A XOR2X1_3/A gnd NAND3X1_61/C vdd OAI21X1
XOAI21X1_557 BUFX4_225/Y OAI21X1_557/B BUFX4_77/Y gnd OAI21X1_557/Y vdd OAI21X1
XOAI21X1_546 OR2X2_7/Y INVX1_192/A OAI21X1_545/Y gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_568 BUFX4_235/Y INVX1_452/A BUFX4_84/Y gnd OAI21X1_568/Y vdd OAI21X1
XOAI21X1_579 BUFX4_148/Y NOR2X1_690/A BUFX4_247/Y gnd OAI21X1_579/Y vdd OAI21X1
XDFFPOSX1_460 INVX1_316/A CLKBUF1_49/Y MUX2X1_366/Y gnd vdd DFFPOSX1
XDFFPOSX1_482 INVX1_431/A CLKBUF1_44/Y DFFPOSX1_482/D gnd vdd DFFPOSX1
XDFFPOSX1_471 INVX1_256/A CLKBUF1_10/Y MUX2X1_372/Y gnd vdd DFFPOSX1
XDFFPOSX1_493 AND2X2_41/B CLKBUF1_65/Y OAI21X1_1486/Y gnd vdd DFFPOSX1
XFILL_5_8_0 gnd vdd FILL
XFILL_13_7_0 gnd vdd FILL
XOAI21X1_332 NOR2X1_84/B BUFX4_309/Y INVX1_406/A gnd OAI21X1_333/C vdd OAI21X1
XOAI21X1_310 BUFX4_137/Y BUFX4_455/Y OAI21X1_310/C gnd OAI21X1_310/Y vdd OAI21X1
XOAI21X1_321 NAND2X1_79/Y BUFX4_218/Y OAI21X1_321/C gnd OAI21X1_321/Y vdd OAI21X1
XOAI21X1_343 BUFX4_467/Y NAND2X1_81/Y OAI21X1_343/C gnd DFFPOSX1_9/D vdd OAI21X1
XOAI21X1_365 BUFX4_372/Y NAND2X1_85/Y OAI21X1_365/C gnd OAI21X1_365/Y vdd OAI21X1
XOAI21X1_354 INVX4_5/A BUFX4_198/Y OAI21X1_878/A gnd OAI21X1_355/C vdd OAI21X1
XOAI21X1_387 OAI21X1_11/A BUFX4_468/Y OAI21X1_387/C gnd DFFPOSX1_77/D vdd OAI21X1
XOAI21X1_376 BUFX4_213/Y OAI21X1_7/B NAND2X1_94/Y gnd OAI21X1_376/Y vdd OAI21X1
XOAI21X1_398 NAND2X1_24/Y BUFX4_213/Y OAI21X1_397/Y gnd OAI21X1_398/Y vdd OAI21X1
XINVX1_407 INVX1_407/A gnd INVX1_407/Y vdd INVX1
XINVX1_429 INVX1_429/A gnd INVX1_429/Y vdd INVX1
XINVX1_418 INVX1_418/A gnd INVX1_418/Y vdd INVX1
XDFFPOSX1_290 OAI21X1_600/B CLKBUF1_83/Y DFFPOSX1_290/D gnd vdd DFFPOSX1
XNAND2X1_360 traffic_Street_0[3] NOR2X1_188/B gnd NAND2X1_360/Y vdd NAND2X1
XFILL_45_6_0 gnd vdd FILL
XFILL_36_6_0 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XFILL_27_6_0 gnd vdd FILL
XAOI22X1_5 AND2X2_8/A INVX2_25/Y INVX2_24/A AOI22X1_5/D gnd AOI22X1_5/Y vdd AOI22X1
XFILL_10_5_0 gnd vdd FILL
XOAI21X1_140 BUFX4_121/Y BUFX4_397/Y OAI21X1_140/C gnd OAI21X1_140/Y vdd OAI21X1
XOAI21X1_173 NAND2X1_56/Y MUX2X1_82/B OAI21X1_173/C gnd OAI21X1_173/Y vdd OAI21X1
XOAI21X1_162 BUFX4_454/Y BUFX4_186/Y AOI21X1_378/A gnd OAI21X1_163/C vdd OAI21X1
XOAI21X1_151 MUX2X1_83/B NAND2X1_51/Y OAI21X1_151/C gnd OAI21X1_151/Y vdd OAI21X1
XINVX1_204 OR2X2_6/B gnd INVX1_204/Y vdd INVX1
XOAI21X1_184 BUFX4_133/Y BUFX4_129/Y OAI21X1_184/C gnd OAI21X1_185/C vdd OAI21X1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XOAI21X1_195 NAND2X1_59/Y BUFX4_174/Y OAI21X1_194/Y gnd OAI21X1_195/Y vdd OAI21X1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XINVX1_259 INVX1_259/A gnd INVX1_259/Y vdd INVX1
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XNAND2X1_15 NOR2X1_4/Y NOR2X1_2/Y gnd BUFX4_302/A vdd NAND2X1
XNAND2X1_37 INVX8_16/A INVX8_9/A gnd NAND2X1_37/Y vdd NAND2X1
XNAND2X1_48 INVX8_18/A INVX4_5/Y gnd NAND2X1_48/Y vdd NAND2X1
XNAND2X1_26 INVX8_10/A INVX8_6/A gnd OAI21X1_48/B vdd NAND2X1
XNAND2X1_59 INVX8_21/A INVX4_3/Y gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_190 NOR2X1_23/A AND2X2_46/B gnd NAND2X1_190/Y vdd NAND2X1
XNOR2X1_617 INVX1_126/A AND2X2_47/B gnd OAI22X1_89/D vdd NOR2X1
XNOR2X1_606 NOR2X1_606/A BUFX4_234/Y gnd OAI22X1_84/D vdd NOR2X1
XFILL_18_6_0 gnd vdd FILL
XNOR2X1_628 NOR2X1_628/A NOR2X1_57/Y gnd NOR2X1_628/Y vdd NOR2X1
XNOR2X1_639 NOR2X1_639/A NOR2X1_76/B gnd NOR2X1_639/Y vdd NOR2X1
XAOI21X1_219 NOR3X1_8/Y AOI21X1_219/B OR2X2_5/A gnd NAND3X1_43/B vdd AOI21X1
XAOI21X1_208 NAND2X1_110/Y NAND2X1_111/Y INVX2_15/Y gnd AOI21X1_208/Y vdd AOI21X1
XAOI22X1_13 AOI22X1_13/A AOI22X1_13/B BUFX4_206/Y OAI22X1_5/Y gnd AOI22X1_13/Y vdd
+ AOI22X1
XAOI22X1_24 AOI22X1_24/A AOI22X1_24/B AOI22X1_24/C AOI22X1_24/D gnd NOR2X1_473/B vdd
+ AOI22X1
XOAI21X1_1403 BUFX4_72/Y NAND2X1_60/Y OAI21X1_1402/Y gnd OAI21X1_1403/Y vdd OAI21X1
XOAI21X1_1414 BUFX4_119/Y BUFX4_408/Y OAI21X1_578/B gnd OAI21X1_1415/C vdd OAI21X1
XOAI21X1_1447 NAND2X1_69/Y BUFX4_444/Y OAI21X1_1446/Y gnd DFFPOSX1_290/D vdd OAI21X1
XOAI21X1_1425 NAND2X1_64/Y BUFX4_430/Y OAI21X1_1425/C gnd OAI21X1_1425/Y vdd OAI21X1
XOAI21X1_1436 BUFX4_123/Y BUFX4_138/Y OAI21X1_1436/C gnd OAI21X1_1437/C vdd OAI21X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XOAI21X1_1469 BUFX4_449/Y BUFX4_160/Y INVX1_374/A gnd OAI21X1_1470/C vdd OAI21X1
XOAI21X1_1458 NAND2X1_70/Y BUFX4_444/Y OAI21X1_1457/Y gnd OAI21X1_1458/Y vdd OAI21X1
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C BUFX4_390/Y gnd OAI22X1_8/Y vdd OAI22X1
XFILL_43_9_1 gnd vdd FILL
XFILL_42_4_0 gnd vdd FILL
XAOI21X1_90 BUFX4_465/Y MUX2X1_96/S NOR2X1_152/Y gnd AOI21X1_90/Y vdd AOI21X1
XBUFX4_321 INVX8_1/Y gnd BUFX4_321/Y vdd BUFX4
XBUFX4_310 INVX8_26/Y gnd BUFX4_310/Y vdd BUFX4
XBUFX4_332 BUFX4_28/Y gnd BUFX4_332/Y vdd BUFX4
XBUFX4_343 BUFX4_28/Y gnd BUFX4_343/Y vdd BUFX4
XBUFX4_354 BUFX4_29/Y gnd BUFX4_354/Y vdd BUFX4
XNOR2X1_403 NOR2X1_403/A AND2X2_37/B gnd OAI22X1_17/D vdd NOR2X1
XNOR2X1_425 NOR2X1_425/A BUFX4_325/Y gnd NOR2X1_425/Y vdd NOR2X1
XBUFX4_398 INVX8_18/Y gnd BUFX4_398/Y vdd BUFX4
XBUFX4_365 BUFX4_27/Y gnd BUFX4_365/Y vdd BUFX4
XNOR2X1_414 BUFX4_102/Y NOR2X1_414/B gnd NOR2X1_414/Y vdd NOR2X1
XBUFX4_376 INVX8_14/Y gnd MUX2X1_44/A vdd BUFX4
XBUFX4_387 BUFX4_384/A gnd BUFX4_387/Y vdd BUFX4
XNOR2X1_436 INVX1_9/A BUFX4_360/Y gnd NOR2X1_436/Y vdd NOR2X1
XNOR2X1_458 NOR2X1_247/A BUFX4_357/Y gnd NOR2X1_458/Y vdd NOR2X1
XNOR2X1_447 NOR2X1_447/A BUFX4_271/Y gnd NOR2X1_447/Y vdd NOR2X1
XFILL_34_9_1 gnd vdd FILL
XFILL_26_2 gnd vdd FILL
XNOR2X1_469 NOR2X1_469/A AND2X2_47/B gnd OAI22X1_35/D vdd NOR2X1
XFILL_33_4_0 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XOAI21X1_909 INVX2_2/Y read_Write BUFX2_6/A gnd OAI21X1_910/C vdd OAI21X1
XOAI21X1_1222 BUFX4_333/Y NOR2X1_264/A BUFX4_146/Y gnd OAI22X1_82/C vdd OAI21X1
XOAI21X1_1200 OAI22X1_72/Y BUFX4_393/Y INVX8_33/Y gnd OAI22X1_81/D vdd OAI21X1
XOAI21X1_1211 AOI21X1_499/Y AOI21X1_500/Y BUFX4_40/Y gnd NAND2X1_346/B vdd OAI21X1
XOAI21X1_1244 BUFX4_341/Y NOR2X1_209/A BUFX4_156/Y gnd OAI22X1_87/C vdd OAI21X1
XMUX2X1_409 BUFX4_426/Y INVX1_329/Y MUX2X1_410/S gnd MUX2X1_409/Y vdd MUX2X1
XOAI21X1_1255 INVX1_140/Y BUFX4_250/Y NAND2X1_348/Y gnd MUX2X1_265/B vdd OAI21X1
XOAI21X1_1233 BUFX4_343/Y NOR2X1_278/A BUFX4_159/Y gnd OAI22X1_83/C vdd OAI21X1
XDFFPOSX1_812 INVX1_91/A CLKBUF1_48/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_823 NOR2X1_121/A CLKBUF1_79/Y AOI21X1_68/Y gnd vdd DFFPOSX1
XDFFPOSX1_801 NOR2X1_108/A CLKBUF1_6/Y AOI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_856 NOR2X1_137/A CLKBUF1_5/Y AOI21X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_834 NOR2X1_129/A CLKBUF1_90/Y AOI21X1_75/Y gnd vdd DFFPOSX1
XOAI21X1_1277 BUFX4_448/Y BUFX4_46/Y NOR2X1_474/B gnd OAI21X1_1277/Y vdd OAI21X1
XOAI21X1_1288 NAND2X1_32/Y MUX2X1_4/B OAI21X1_1287/Y gnd DFFPOSX1_145/D vdd OAI21X1
XDFFPOSX1_845 INVX1_394/A CLKBUF1_26/Y OAI21X1_173/Y gnd vdd DFFPOSX1
XOAI21X1_1266 NAND2X1_30/Y BUFX4_442/Y OAI21X1_1265/Y gnd OAI21X1_1266/Y vdd OAI21X1
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XDFFPOSX1_867 INVX1_105/A CLKBUF1_26/Y MUX2X1_92/Y gnd vdd DFFPOSX1
XOAI21X1_1299 BUFX4_440/Y NAND2X1_37/Y OAI21X1_1299/C gnd DFFPOSX1_206/D vdd OAI21X1
XDFFPOSX1_889 MUX2X1_245/B CLKBUF1_74/Y OAI21X1_205/Y gnd vdd DFFPOSX1
XDFFPOSX1_878 NOR2X1_585/A CLKBUF1_74/Y AOI21X1_90/Y gnd vdd DFFPOSX1
XFILL_0_9_1 gnd vdd FILL
XFILL_25_9_1 gnd vdd FILL
XFILL_24_4_0 gnd vdd FILL
XAOI21X1_561 BUFX4_65/Y NOR2X1_137/B NOR2X1_673/Y gnd AOI21X1_561/Y vdd AOI21X1
XAOI21X1_550 BUFX4_428/Y NAND2X1_50/B NOR2X1_662/Y gnd AOI21X1_550/Y vdd AOI21X1
XAOI21X1_594 MUX2X1_29/B NOR2X1_703/B NOR2X1_706/Y gnd AOI21X1_594/Y vdd AOI21X1
XAOI21X1_583 BUFX4_66/Y MUX2X1_102/S NOR2X1_695/Y gnd AOI21X1_583/Y vdd AOI21X1
XAOI21X1_572 BUFX4_422/Y NOR2X1_155/B NOR2X1_684/Y gnd AOI21X1_572/Y vdd AOI21X1
XFILL_7_5_0 gnd vdd FILL
XFILL_16_9_1 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XMUX2X1_1 INVX1_4/Y MUX2X1_1/B MUX2X1_2/S gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_119 NOR2X1_291/A CLKBUF1_88/Y AOI21X1_194/Y gnd vdd DFFPOSX1
XDFFPOSX1_108 INVX1_402/A CLKBUF1_51/Y OAI21X1_410/Y gnd vdd DFFPOSX1
XCLKBUF1_2 BUFX4_6/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XNOR2X1_200 NOR2X1_200/A NOR2X1_703/B gnd NOR2X1_200/Y vdd NOR2X1
XBUFX4_151 INVX8_32/Y gnd BUFX4_151/Y vdd BUFX4
XBUFX4_173 INVX8_13/Y gnd BUFX4_173/Y vdd BUFX4
XBUFX4_162 INVX8_24/Y gnd BUFX4_162/Y vdd BUFX4
XBUFX4_140 INVX8_22/Y gnd BUFX4_140/Y vdd BUFX4
XNOR2X1_211 NOR2X1_211/A MUX2X1_120/S gnd NOR2X1_211/Y vdd NOR2X1
XNOR2X1_233 BUFX4_455/Y BUFX4_120/Y gnd NOR2X1_233/Y vdd NOR2X1
XBUFX4_195 INVX8_27/Y gnd BUFX4_195/Y vdd BUFX4
XBUFX4_184 INVX8_19/Y gnd BUFX4_184/Y vdd BUFX4
XNOR2X1_222 BUFX4_457/Y BUFX4_56/Y gnd NOR2X1_716/B vdd NOR2X1
XNOR2X1_255 BUFX4_312/Y BUFX4_120/Y gnd MUX2X1_397/S vdd NOR2X1
XNOR2X1_266 NOR2X1_266/A NOR2X1_737/B gnd NOR2X1_266/Y vdd NOR2X1
XNOR2X1_244 AND2X2_55/A NOR2X1_727/B gnd NOR2X1_244/Y vdd NOR2X1
XNOR2X1_299 traffic_Street_1[0] traffic_Street_1[1] gnd NOR2X1_299/Y vdd NOR2X1
XNOR2X1_277 NOR2X1_277/A NOR2X1_16/Y gnd NOR2X1_277/Y vdd NOR2X1
XNOR2X1_288 NOR2X1_288/A NOR2X1_33/Y gnd NOR2X1_288/Y vdd NOR2X1
XOAI21X1_706 BUFX4_366/Y INVX1_49/A BUFX4_152/Y gnd OAI22X1_18/C vdd OAI21X1
XOAI21X1_728 INVX1_294/Y BUFX4_249/Y BUFX4_149/Y gnd OAI21X1_728/Y vdd OAI21X1
XOAI21X1_739 OAI21X1_739/A OAI21X1_739/B BUFX4_38/Y gnd NAND2X1_230/B vdd OAI21X1
XOAI21X1_717 OAI21X1_134/C BUFX4_241/Y BUFX4_97/Y gnd OAI21X1_717/Y vdd OAI21X1
XOAI21X1_1030 BUFX4_365/Y OAI21X1_113/C BUFX4_152/Y gnd AOI21X1_442/C vdd OAI21X1
XOAI21X1_1063 OAI21X1_252/C BUFX4_240/Y BUFX4_76/Y gnd OAI22X1_47/B vdd OAI21X1
XOAI21X1_1041 OAI21X1_401/C BUFX4_289/Y BUFX4_112/Y gnd OAI22X1_45/B vdd OAI21X1
XMUX2X1_217 MUX2X1_217/A MUX2X1_217/B BUFX4_411/Y gnd MUX2X1_217/Y vdd MUX2X1
XDFFPOSX1_631 INVX1_28/A CLKBUF1_81/Y MUX2X1_21/Y gnd vdd DFFPOSX1
XOAI21X1_1052 NOR2X1_510/Y AOI21X1_451/Y BUFX4_36/Y gnd OAI21X1_1055/C vdd OAI21X1
XDFFPOSX1_620 INVX1_330/A CLKBUF1_73/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XMUX2X1_228 MUX2X1_228/A MUX2X1_228/B BUFX4_85/Y gnd MUX2X1_228/Y vdd MUX2X1
XMUX2X1_206 MUX2X1_206/A MUX2X1_206/B BUFX4_96/Y gnd MUX2X1_206/Y vdd MUX2X1
XDFFPOSX1_664 INVX1_35/A CLKBUF1_4/Y MUX2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_653 NOR2X1_35/A CLKBUF1_84/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_642 NOR2X1_560/A CLKBUF1_103/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XMUX2X1_239 MUX2X1_239/A MUX2X1_239/B BUFX4_78/Y gnd MUX2X1_239/Y vdd MUX2X1
XDFFPOSX1_675 NOR2X1_45/A CLKBUF1_87/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XOAI21X1_1074 NOR2X1_517/Y NOR2X1_518/Y BUFX4_357/Y gnd NAND3X1_80/C vdd OAI21X1
XOAI21X1_1085 BUFX4_152/Y INVX1_410/Y AOI21X1_462/Y gnd AOI21X1_464/A vdd OAI21X1
XOAI21X1_1096 BUFX4_271/Y OAI21X1_1096/B BUFX4_94/Y gnd OAI21X1_1096/Y vdd OAI21X1
XDFFPOSX1_697 NOR2X1_63/A CLKBUF1_70/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_686 OAI21X1_65/C CLKBUF1_100/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XFILL_40_7_1 gnd vdd FILL
XINVX8_4 traffic_Street_0[2] gnd INVX8_4/Y vdd INVX8
XAOI21X1_380 BUFX4_153/Y OAI21X1_860/Y AOI21X1_379/Y gnd MUX2X1_221/A vdd AOI21X1
XAOI21X1_391 AOI21X1_391/A NAND3X1_75/Y BUFX4_401/Y gnd OAI21X1_907/B vdd AOI21X1
XDFFPOSX1_90 INVX1_278/A CLKBUF1_66/Y DFFPOSX1_90/D gnd vdd DFFPOSX1
XBUFX4_24 address[0] gnd BUFX4_24/Y vdd BUFX4
XBUFX4_13 address[1] gnd BUFX4_82/A vdd BUFX4
XBUFX4_35 BUFX4_33/A gnd BUFX4_35/Y vdd BUFX4
XFILL_48_8_1 gnd vdd FILL
XBUFX4_46 BUFX4_46/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_57 INVX8_6/Y gnd BUFX4_57/Y vdd BUFX4
XBUFX4_68 INVX8_4/Y gnd BUFX4_68/Y vdd BUFX4
XFILL_47_3_0 gnd vdd FILL
XBUFX4_79 BUFX4_14/Y gnd BUFX4_79/Y vdd BUFX4
XFILL_31_7_1 gnd vdd FILL
XFILL_30_2_0 gnd vdd FILL
XFILL_39_8_1 gnd vdd FILL
XFILL_38_3_0 gnd vdd FILL
XINVX8_16 INVX8_16/A gnd INVX8_16/Y vdd INVX8
XINVX8_27 INVX8_27/A gnd INVX8_27/Y vdd INVX8
XFILL_22_7_1 gnd vdd FILL
XOAI21X1_503 BUFX4_306/Y INVX4_11/Y NAND3X1_46/B gnd INVX1_206/A vdd OAI21X1
XOAI21X1_514 NOR3X1_12/Y OAI21X1_504/Y AOI22X1_6/Y gnd AOI21X1_238/B vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_525 OR2X2_6/Y NOR2X1_331/Y AOI22X1_6/B gnd INVX1_210/A vdd OAI21X1
XOAI21X1_536 XNOR2X1_6/Y OAI21X1_534/Y OAI21X1_536/C gnd OAI21X1_536/Y vdd OAI21X1
XOAI21X1_547 XNOR2X1_8/A INVX2_4/Y NOR2X1_1/B gnd OAI21X1_547/Y vdd OAI21X1
XOAI21X1_558 AOI21X1_250/Y AOI21X1_251/Y BUFX4_410/Y gnd OAI21X1_558/Y vdd OAI21X1
XOAI21X1_569 AND2X2_51/B INVX1_232/Y OAI21X1_569/C gnd OAI21X1_571/C vdd OAI21X1
XDFFPOSX1_450 INVX1_429/A CLKBUF1_82/Y MUX2X1_364/Y gnd vdd DFFPOSX1
XDFFPOSX1_483 AOI21X1_273/B CLKBUF1_68/Y OAI21X1_1474/Y gnd vdd DFFPOSX1
XDFFPOSX1_461 INVX1_382/A CLKBUF1_10/Y MUX2X1_367/Y gnd vdd DFFPOSX1
XDFFPOSX1_472 NOR2X1_712/A CLKBUF1_50/Y AOI21X1_600/Y gnd vdd DFFPOSX1
XDFFPOSX1_494 AND2X2_52/B CLKBUF1_13/Y DFFPOSX1_494/D gnd vdd DFFPOSX1
XFILL_5_8_1 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_29_3_0 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XOAI21X1_311 MUX2X1_83/B NAND2X1_77/Y OAI21X1_310/Y gnd OAI21X1_311/Y vdd OAI21X1
XOAI21X1_322 BUFX4_386/Y BUFX4_311/Y OAI21X1_889/A gnd OAI21X1_323/C vdd OAI21X1
XOAI21X1_300 BUFX4_386/Y BUFX4_458/Y NOR2X1_517/A gnd OAI21X1_301/C vdd OAI21X1
XOAI21X1_333 NAND2X1_80/Y MUX2X1_86/B OAI21X1_333/C gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_355 NAND2X1_84/Y MUX2X1_40/B OAI21X1_355/C gnd OAI21X1_355/Y vdd OAI21X1
XOAI21X1_344 INVX4_3/A BUFX4_199/Y INVX1_277/A gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_388 INVX1_179/Y AOI21X1_7/B NAND2X1_98/Y gnd OAI21X1_388/Y vdd OAI21X1
XOAI21X1_366 BUFX4_191/Y BUFX4_198/Y INVX1_443/A gnd OAI21X1_367/C vdd OAI21X1
XOAI21X1_377 BUFX4_178/Y OAI21X1_7/B NAND2X1_95/Y gnd DFFPOSX1_71/D vdd OAI21X1
XOAI21X1_399 BUFX4_121/Y NOR2X1_16/A OAI21X1_868/A gnd OAI21X1_399/Y vdd OAI21X1
XINVX1_408 INVX1_408/A gnd INVX1_408/Y vdd INVX1
XINVX1_419 INVX1_419/A gnd INVX1_419/Y vdd INVX1
XDFFPOSX1_280 INVX1_352/A CLKBUF1_69/Y MUX2X1_330/Y gnd vdd DFFPOSX1
XDFFPOSX1_291 INVX1_318/A CLKBUF1_50/Y OAI21X1_1449/Y gnd vdd DFFPOSX1
XNAND2X1_361 NAND2X1_361/A NAND2X1_2/Y gnd NAND2X1_361/Y vdd NAND2X1
XNAND2X1_350 DFFPOSX1_1/Q BUFX4_253/Y gnd NAND2X1_350/Y vdd NAND2X1
XFILL_45_6_1 gnd vdd FILL
XFILL_44_1_0 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XFILL_36_6_1 gnd vdd FILL
XFILL_35_1_0 gnd vdd FILL
XNAND3X1_1 NOR2X1_2/A INVX1_1/A NOR2X1_6/Y gnd MUX2X1_2/S vdd NAND3X1
XFILL_2_6_1 gnd vdd FILL
XFILL_27_6_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XOAI21X1_130 MUX2X1_61/B NAND2X1_44/Y OAI21X1_129/Y gnd OAI21X1_130/Y vdd OAI21X1
XAOI22X1_6 AOI22X1_6/A AOI22X1_6/B AOI22X1_6/C AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_174 BUFX4_131/Y BUFX4_297/Y NOR2X1_595/A gnd OAI21X1_174/Y vdd OAI21X1
XOAI21X1_163 NAND2X1_53/Y BUFX4_180/Y OAI21X1_163/C gnd OAI21X1_163/Y vdd OAI21X1
XOAI21X1_152 BUFX4_386/Y BUFX4_187/Y OAI21X1_678/A gnd OAI21X1_153/C vdd OAI21X1
XOAI21X1_141 NAND2X1_48/Y MUX2X1_58/A OAI21X1_140/Y gnd OAI21X1_141/Y vdd OAI21X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_216 police_Interrupt gnd AND2X2_18/B vdd INVX1
XOAI21X1_185 BUFX4_214/Y NAND2X1_58/Y OAI21X1_185/C gnd OAI21X1_185/Y vdd OAI21X1
XOAI21X1_196 BUFX4_387/Y BUFX4_406/Y INVX1_397/A gnd OAI21X1_197/C vdd OAI21X1
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XINVX1_227 INVX1_227/A gnd INVX1_227/Y vdd INVX1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_16 INVX8_5/A INVX4_2/Y gnd OAI21X1_11/A vdd NAND2X1
XNAND2X1_180 BUFX4_260/Y INVX1_455/A gnd NAND2X1_180/Y vdd NAND2X1
XNAND2X1_49 traffic_Street_1[1] NAND2X1_50/B gnd NAND2X1_49/Y vdd NAND2X1
XNAND2X1_38 INVX8_17/A INVX4_2/Y gnd MUX2X1_51/S vdd NAND2X1
XNAND2X1_27 INVX8_10/A INVX4_3/Y gnd MUX2X1_29/S vdd NAND2X1
XNAND2X1_191 BUFX4_36/Y MUX2X1_187/Y gnd AOI22X1_16/A vdd NAND2X1
XNOR2X1_607 NOR2X1_289/A BUFX4_332/Y gnd OAI22X1_84/A vdd NOR2X1
XFILL_18_6_1 gnd vdd FILL
XNOR2X1_618 NOR2X1_190/A BUFX4_340/Y gnd OAI22X1_89/A vdd NOR2X1
XNOR2X1_629 NOR2X1_629/A NOR2X1_60/Y gnd NOR2X1_629/Y vdd NOR2X1
XFILL_17_1_0 gnd vdd FILL
XAOI21X1_209 NAND3X1_14/B OR2X2_4/Y BUFX4_320/Y gnd NAND3X1_20/C vdd AOI21X1
XAOI22X1_14 AOI22X1_14/A AOI22X1_14/B BUFX4_400/Y MUX2X1_180/Y gnd AOI22X1_14/Y vdd
+ AOI22X1
XAOI22X1_25 AOI22X1_25/A AOI22X1_25/B NAND3X1_77/Y AOI22X1_25/D gnd AOI22X1_25/Y vdd
+ AOI22X1
XOAI21X1_1404 BUFX4_143/Y BUFX4_403/Y NOR2X1_534/A gnd OAI21X1_1405/C vdd OAI21X1
XOAI21X1_1426 BUFX4_383/Y BUFX4_140/Y AND2X2_39/B gnd OAI21X1_1426/Y vdd OAI21X1
XOAI21X1_1437 NAND2X1_66/Y BUFX4_317/Y OAI21X1_1437/C gnd DFFPOSX1_265/D vdd OAI21X1
XOAI21X1_1415 NAND2X1_62/Y BUFX4_445/Y OAI21X1_1415/C gnd OAI21X1_1415/Y vdd OAI21X1
XOAI21X1_1459 BUFX4_126/Y BUFX4_435/Y NAND2X1_238/A gnd OAI21X1_1460/C vdd OAI21X1
XNOR3X1_4 INVX4_8/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XOAI21X1_1448 BUFX4_384/Y BUFX4_431/Y INVX1_318/A gnd OAI21X1_1449/C vdd OAI21X1
XOAI22X1_9 OAI22X1_9/A OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XFILL_42_4_1 gnd vdd FILL
XAOI21X1_80 MUX2X1_49/A NOR2X1_137/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XAOI21X1_91 AND2X2_2/B NOR2X1_155/B AOI21X1_91/C gnd AOI21X1_91/Y vdd AOI21X1
XFILL_49_0_0 gnd vdd FILL
XBUFX4_322 INVX8_1/Y gnd BUFX4_322/Y vdd BUFX4
XBUFX4_311 INVX8_26/Y gnd BUFX4_311/Y vdd BUFX4
XBUFX4_300 BUFX4_302/A gnd BUFX4_300/Y vdd BUFX4
XBUFX4_355 BUFX4_25/Y gnd BUFX4_355/Y vdd BUFX4
XBUFX4_344 BUFX4_30/Y gnd BUFX4_344/Y vdd BUFX4
XBUFX4_333 BUFX4_26/Y gnd BUFX4_333/Y vdd BUFX4
XNOR2X1_404 NOR2X1_71/A BUFX4_334/Y gnd NOR2X1_404/Y vdd NOR2X1
XBUFX4_388 BUFX4_384/A gnd NOR2X1_77/B vdd BUFX4
XNOR2X1_415 BUFX4_364/Y INVX1_295/Y gnd NOR2X1_416/A vdd NOR2X1
XBUFX4_366 BUFX4_27/Y gnd BUFX4_366/Y vdd BUFX4
XBUFX4_377 INVX8_14/Y gnd BUFX4_377/Y vdd BUFX4
XNOR2X1_426 BUFX4_414/Y OAI22X1_21/Y gnd NOR2X1_426/Y vdd NOR2X1
XNOR2X1_437 BUFX4_49/Y NOR2X1_437/B gnd NOR2X1_437/Y vdd NOR2X1
XBUFX4_399 address[5] gnd INVX8_33/A vdd BUFX4
XNOR2X1_459 NOR2X1_459/A BUFX4_235/Y gnd NOR2X1_459/Y vdd NOR2X1
XNOR2X1_448 NOR2X1_165/A BUFX4_331/Y gnd NOR2X1_448/Y vdd NOR2X1
XFILL_26_3 gnd vdd FILL
XFILL_33_4_1 gnd vdd FILL
XFILL_19_2 gnd vdd FILL
XOAI21X1_1212 BUFX4_330/Y OAI21X1_150/C BUFX4_153/Y gnd OAI22X1_76/C vdd OAI21X1
XOAI21X1_1201 INVX1_119/A BUFX4_280/Y AOI21X1_498/Y gnd OAI21X1_1203/C vdd OAI21X1
XOAI21X1_1234 INVX1_178/A BUFX4_233/Y BUFX4_102/Y gnd OAI22X1_83/B vdd OAI21X1
XOAI21X1_1256 INVX1_144/Y BUFX4_252/Y NAND2X1_349/Y gnd MUX2X1_265/A vdd OAI21X1
XOAI21X1_1223 OAI21X1_350/C BUFX4_226/Y BUFX4_98/Y gnd OAI22X1_82/B vdd OAI21X1
XDFFPOSX1_824 NOR2X1_122/A CLKBUF1_42/Y AOI21X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_802 NOR2X1_109/A CLKBUF1_51/Y AOI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_813 INVX1_92/A CLKBUF1_44/Y OAI21X1_143/Y gnd vdd DFFPOSX1
XOAI21X1_1245 NOR2X1_212/A BUFX4_240/Y AND2X2_32/B gnd OAI22X1_87/B vdd OAI21X1
XDFFPOSX1_857 NOR2X1_138/A CLKBUF1_62/Y AOI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_846 NOR2X1_595/A CLKBUF1_53/Y OAI21X1_175/Y gnd vdd DFFPOSX1
XOAI21X1_1278 NAND2X1_31/Y BUFX4_64/Y OAI21X1_1277/Y gnd DFFPOSX1_148/D vdd OAI21X1
XOAI21X1_1267 BUFX4_301/Y BUFX4_45/Y NOR2X1_420/B gnd OAI21X1_1268/C vdd OAI21X1
XDFFPOSX1_835 INVX1_93/A CLKBUF1_2/Y MUX2X1_80/Y gnd vdd DFFPOSX1
XOAI21X1_1289 INVX1_301/Y NOR2X1_76/B NAND2X1_353/Y gnd DFFPOSX1_215/D vdd OAI21X1
XDFFPOSX1_879 NOR2X1_154/A CLKBUF1_101/Y AOI21X1_91/Y gnd vdd DFFPOSX1
XDFFPOSX1_868 NOR2X1_143/A CLKBUF1_2/Y AOI21X1_84/Y gnd vdd DFFPOSX1
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XFILL_24_4_1 gnd vdd FILL
XAOI21X1_540 MUX2X1_29/B NOR2X1_97/B NOR2X1_652/Y gnd AOI21X1_540/Y vdd AOI21X1
XAOI21X1_562 BUFX4_321/Y NOR2X1_137/B NOR2X1_674/Y gnd AOI21X1_562/Y vdd AOI21X1
XAOI21X1_551 BUFX4_318/Y NAND2X1_50/B NOR2X1_663/Y gnd AOI21X1_551/Y vdd AOI21X1
XAOI21X1_584 BUFX4_317/Y MUX2X1_102/S NOR2X1_696/Y gnd AOI21X1_584/Y vdd AOI21X1
XAOI21X1_595 BUFX4_444/Y NOR2X1_707/B NOR2X1_707/Y gnd AOI21X1_595/Y vdd AOI21X1
XAOI21X1_573 BUFX4_73/Y NOR2X1_155/B NOR2X1_685/Y gnd AOI21X1_573/Y vdd AOI21X1
XFILL_7_5_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd INVX2_22/A vdd XOR2X1
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 INVX1_5/Y MUX2X1_6/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XDFFPOSX1_109 NOR2X1_608/A CLKBUF1_63/Y OAI21X1_412/Y gnd vdd DFFPOSX1
XCLKBUF1_3 BUFX4_4/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XBUFX4_130 INVX8_20/Y gnd BUFX4_130/Y vdd BUFX4
XBUFX4_152 INVX8_32/Y gnd BUFX4_152/Y vdd BUFX4
XBUFX4_163 INVX8_24/Y gnd BUFX4_163/Y vdd BUFX4
XBUFX4_141 INVX8_22/Y gnd BUFX4_141/Y vdd BUFX4
XNOR2X1_234 BUFX4_455/Y BUFX4_193/Y gnd NOR2X1_234/Y vdd NOR2X1
XBUFX4_185 INVX8_19/Y gnd BUFX4_185/Y vdd BUFX4
XBUFX4_196 INVX8_27/Y gnd BUFX4_196/Y vdd BUFX4
XNOR2X1_201 INVX2_1/Y INVX2_12/Y gnd INVX8_24/A vdd NOR2X1
XNOR2X1_223 NOR2X1_223/A NOR2X1_716/B gnd NOR2X1_223/Y vdd NOR2X1
XBUFX4_174 INVX8_13/Y gnd BUFX4_174/Y vdd BUFX4
XNOR2X1_212 NOR2X1_212/A MUX2X1_120/S gnd NOR2X1_212/Y vdd NOR2X1
XNOR2X1_267 NOR2X1_454/A NOR2X1_737/B gnd NOR2X1_267/Y vdd NOR2X1
XNOR2X1_256 INVX2_10/Y INVX2_6/Y gnd INVX8_27/A vdd NOR2X1
XNOR2X1_245 BUFX4_311/Y BUFX4_142/Y gnd NOR2X1_729/B vdd NOR2X1
XFILL_31_1 gnd vdd FILL
XNOR2X1_289 NOR2X1_289/A NOR2X1_33/Y gnd NOR2X1_289/Y vdd NOR2X1
XNOR2X1_278 NOR2X1_278/A NOR2X1_16/Y gnd NOR2X1_278/Y vdd NOR2X1
XOAI21X1_729 INVX1_296/Y BUFX4_251/Y BUFX4_103/Y gnd NOR2X1_416/B vdd OAI21X1
XOAI21X1_707 NOR2X1_78/A BUFX4_235/Y BUFX4_95/Y gnd OAI22X1_18/B vdd OAI21X1
XOAI21X1_718 OAI21X1_718/A OAI21X1_718/B BUFX4_418/Y gnd AOI21X1_316/B vdd OAI21X1
XOAI21X1_1020 INVX1_44/Y BUFX4_268/Y NAND2X1_309/Y gnd AOI21X1_438/B vdd OAI21X1
XOAI21X1_1031 INVX1_67/Y BUFX4_277/Y NAND2X1_314/Y gnd AOI21X1_443/B vdd OAI21X1
XDFFPOSX1_610 INVX1_17/A CLKBUF1_80/Y MUX2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_632 INVX1_29/A CLKBUF1_30/Y MUX2X1_22/Y gnd vdd DFFPOSX1
XOAI21X1_1053 BUFX4_326/Y INVX1_169/A BUFX4_159/Y gnd AOI21X1_452/C vdd OAI21X1
XOAI21X1_1042 AOI21X1_447/Y BUFX4_419/Y NAND2X1_319/Y gnd NOR2X1_507/B vdd OAI21X1
XDFFPOSX1_621 NAND2X1_13/A CLKBUF1_25/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XMUX2X1_229 MUX2X1_229/A MUX2X1_229/B BUFX4_86/Y gnd MUX2X1_229/Y vdd MUX2X1
XMUX2X1_218 MUX2X1_218/A OAI22X1_25/Y BUFX4_170/Y gnd MUX2X1_218/Y vdd MUX2X1
XMUX2X1_207 MUX2X1_207/A MUX2X1_207/B INVX8_33/Y gnd MUX2X1_207/Y vdd MUX2X1
XOAI21X1_1064 AOI21X1_454/Y BUFX4_33/Y NAND2X1_327/Y gnd AOI22X1_32/B vdd OAI21X1
XDFFPOSX1_665 INVX1_36/A CLKBUF1_4/Y MUX2X1_28/Y gnd vdd DFFPOSX1
XOAI21X1_1086 BUFX4_151/Y INVX1_411/Y AOI21X1_463/Y gnd AOI21X1_464/B vdd OAI21X1
XDFFPOSX1_654 NOR2X1_36/A CLKBUF1_84/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_643 NOR2X1_28/A CLKBUF1_76/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XOAI21X1_1075 BUFX4_32/Y MUX2X1_254/Y NAND3X1_80/Y gnd NOR2X1_519/B vdd OAI21X1
XOAI21X1_1097 NOR2X1_525/Y OAI21X1_1096/Y OAI21X1_1095/Y gnd NOR2X1_526/B vdd OAI21X1
XDFFPOSX1_698 NOR2X1_64/A CLKBUF1_53/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_687 NOR2X1_55/A CLKBUF1_43/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_676 NOR2X1_46/A CLKBUF1_87/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XAOI21X1_370 BUFX4_50/Y AOI22X1_21/Y INVX8_33/A gnd AOI22X1_23/C vdd AOI21X1
XAOI21X1_381 INVX1_176/Y BUFX4_349/Y BUFX4_159/Y gnd AOI21X1_381/Y vdd AOI21X1
XAOI21X1_392 street OAI21X1_908/Y AOI21X1_392/C gnd AOI21X1_392/Y vdd AOI21X1
XDFFPOSX1_80 NOR2X1_277/A CLKBUF1_91/Y DFFPOSX1_80/D gnd vdd DFFPOSX1
XDFFPOSX1_91 NOR2X1_451/A CLKBUF1_40/Y DFFPOSX1_91/D gnd vdd DFFPOSX1
XBUFX4_14 address[1] gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 BUFX4_28/A gnd BUFX4_25/Y vdd BUFX4
XBUFX4_36 BUFX4_33/A gnd BUFX4_36/Y vdd BUFX4
XBUFX4_69 INVX8_4/Y gnd BUFX4_69/Y vdd BUFX4
XBUFX4_47 address[4] gnd INVX8_28/A vdd BUFX4
XBUFX4_58 INVX8_6/Y gnd BUFX4_58/Y vdd BUFX4
XFILL_47_3_1 gnd vdd FILL
XFILL_30_2_1 gnd vdd FILL
XFILL_38_3_1 gnd vdd FILL
XINVX8_17 INVX8_17/A gnd BUFX4_54/A vdd INVX8
XINVX8_28 INVX8_28/A gnd INVX8_28/Y vdd INVX8
XOAI21X1_504 INVX1_206/Y NAND3X1_47/Y NAND2X1_146/Y gnd OAI21X1_504/Y vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_515 OAI21X1_515/A INVX1_207/Y NAND3X1_58/A gnd OAI21X1_515/Y vdd OAI21X1
XOAI21X1_526 OAI21X1_515/Y INVX1_210/Y INVX4_9/Y gnd OAI21X1_528/A vdd OAI21X1
XOAI21X1_537 INVX4_12/Y INVX2_26/Y OAI21X1_497/A gnd AOI21X1_245/C vdd OAI21X1
XOAI21X1_548 INVX2_5/Y XNOR2X1_8/A OAI21X1_547/Y gnd OAI21X1_548/Y vdd OAI21X1
XOAI21X1_559 AOI21X1_249/Y BUFX4_411/Y OAI21X1_558/Y gnd AOI22X1_11/C vdd OAI21X1
XDFFPOSX1_440 NOR2X1_630/A CLKBUF1_24/Y AOI21X1_518/Y gnd vdd DFFPOSX1
XDFFPOSX1_451 NOR2X1_703/A CLKBUF1_37/Y AOI21X1_591/Y gnd vdd DFFPOSX1
XDFFPOSX1_473 INVX1_378/A CLKBUF1_4/Y MUX2X1_373/Y gnd vdd DFFPOSX1
XDFFPOSX1_462 INVX1_430/A CLKBUF1_50/Y MUX2X1_368/Y gnd vdd DFFPOSX1
XDFFPOSX1_495 INVX1_264/A CLKBUF1_18/Y OAI21X1_1490/Y gnd vdd DFFPOSX1
XDFFPOSX1_484 INVX1_319/A CLKBUF1_74/Y OAI21X1_1476/Y gnd vdd DFFPOSX1
XFILL_4_3_1 gnd vdd FILL
XFILL_29_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XOAI21X1_323 NAND2X1_79/Y BUFX4_176/Y OAI21X1_323/C gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_312 BUFX4_313/Y BUFX4_300/Y NOR2X1_381/A gnd OAI21X1_313/C vdd OAI21X1
XOAI21X1_301 NAND2X1_76/Y BUFX4_380/Y OAI21X1_301/C gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_334 NOR2X1_84/B BUFX4_308/Y INVX1_444/A gnd OAI21X1_335/C vdd OAI21X1
XOAI21X1_356 INVX4_5/A BUFX4_195/Y INVX1_404/A gnd OAI21X1_356/Y vdd OAI21X1
XOAI21X1_345 NAND2X1_82/Y BUFX4_214/Y OAI21X1_344/Y gnd OAI21X1_345/Y vdd OAI21X1
XOAI21X1_389 BUFX4_450/Y BUFX4_293/Y INVX1_278/A gnd OAI21X1_389/Y vdd OAI21X1
XOAI21X1_367 BUFX4_473/Y NAND2X1_85/Y OAI21X1_367/C gnd DFFPOSX1_41/D vdd OAI21X1
XOAI21X1_378 BUFX4_372/Y OAI21X1_7/B NAND2X1_96/Y gnd OAI21X1_378/Y vdd OAI21X1
XINVX1_409 BUFX2_8/A gnd INVX1_409/Y vdd INVX1
XDFFPOSX1_270 INVX1_243/A CLKBUF1_31/Y DFFPOSX1_270/D gnd vdd DFFPOSX1
XDFFPOSX1_281 INVX1_422/A CLKBUF1_69/Y MUX2X1_331/Y gnd vdd DFFPOSX1
XDFFPOSX1_292 OAI21X1_958/B CLKBUF1_10/Y DFFPOSX1_292/D gnd vdd DFFPOSX1
XNAND2X1_351 DFFPOSX1_9/Q BUFX4_255/Y gnd NAND2X1_351/Y vdd NAND2X1
XNAND2X1_362 NAND2X1_362/A NAND2X1_2/Y gnd NAND2X1_362/Y vdd NAND2X1
XNAND2X1_340 NAND2X1_340/A BUFX4_336/Y gnd NAND2X1_340/Y vdd NAND2X1
XFILL_44_1_1 gnd vdd FILL
XOAI21X1_890 NOR2X1_458/Y OAI21X1_890/B OAI21X1_888/Y gnd AOI21X1_389/B vdd OAI21X1
XFILL_7_2 gnd vdd FILL
XMUX2X1_390 BUFX4_429/Y INVX1_324/Y NOR2X1_727/B gnd MUX2X1_390/Y vdd MUX2X1
XFILL_35_1_1 gnd vdd FILL
XNAND3X1_2 NOR2X1_2/A INVX2_5/A NOR2X1_6/Y gnd MUX2X1_6/S vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XOAI21X1_120 NAND2X1_40/Y MUX2X1_64/B OAI21X1_119/Y gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_131 BUFX4_58/Y BUFX4_397/Y OAI21X1_131/C gnd OAI21X1_132/C vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AOI22X1_7/B AOI22X1_7/C AND2X2_13/Y gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_164 BUFX4_454/Y BUFX4_185/Y INVX1_396/A gnd OAI21X1_164/Y vdd OAI21X1
XOAI21X1_142 INVX1_91/Y NAND2X1_50/B NAND2X1_49/Y gnd OAI21X1_142/Y vdd OAI21X1
XOAI21X1_153 NAND2X1_52/Y BUFX4_218/Y OAI21X1_153/C gnd OAI21X1_153/Y vdd OAI21X1
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XOAI21X1_175 NAND2X1_56/Y MUX2X1_83/B OAI21X1_174/Y gnd OAI21X1_175/Y vdd OAI21X1
XOAI21X1_186 BUFX4_137/Y BUFX4_128/Y NAND2X1_257/A gnd OAI21X1_186/Y vdd OAI21X1
XOAI21X1_197 NAND2X1_59/Y MUX2X1_57/A OAI21X1_197/C gnd OAI21X1_197/Y vdd OAI21X1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XINVX1_228 INVX1_228/A gnd INVX1_228/Y vdd INVX1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_170 BUFX4_223/Y NOR2X1_629/A gnd NAND2X1_170/Y vdd NAND2X1
XNAND2X1_17 NOR2X1_2/A NOR2X1_4/Y gnd XNOR2X1_8/A vdd NAND2X1
XNAND2X1_28 INVX8_10/A INVX4_4/Y gnd OAI21X1_54/A vdd NAND2X1
XNAND2X1_39 INVX8_17/A INVX8_6/A gnd NAND2X1_39/Y vdd NAND2X1
XNAND2X1_192 NOR2X1_28/A INVX8_31/A gnd NAND2X1_192/Y vdd NAND2X1
XNAND2X1_181 BUFX4_391/Y NAND2X1_181/B gnd AOI22X1_17/A vdd NAND2X1
XFILL_46_9_0 gnd vdd FILL
XNOR2X1_608 NOR2X1_608/A BUFX4_236/Y gnd NOR2X1_608/Y vdd NOR2X1
XNOR2X1_619 NOR2X1_619/A AND2X2_52/A gnd NOR2X1_619/Y vdd NOR2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 AOI22X1_15/A AOI22X1_15/B BUFX4_165/Y AOI22X1_15/D gnd AOI22X1_15/Y vdd
+ AOI22X1
XAOI22X1_26 AOI22X1_26/A AOI22X1_26/B AOI22X1_26/C BUFX4_167/Y gnd AOI22X1_26/Y vdd
+ AOI22X1
XOAI21X1_1405 BUFX4_320/Y NAND2X1_60/Y OAI21X1_1405/C gnd DFFPOSX1_189/D vdd OAI21X1
XOAI21X1_1438 BUFX4_60/Y BUFX4_432/Y OAI21X1_599/B gnd OAI21X1_1439/C vdd OAI21X1
XOAI21X1_1427 NAND2X1_64/Y BUFX4_66/Y OAI21X1_1426/Y gnd DFFPOSX1_212/D vdd OAI21X1
XOAI21X1_1416 BUFX4_119/Y BUFX4_407/Y OAI21X1_754/B gnd OAI21X1_1417/C vdd OAI21X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_4/Y NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XOAI21X1_1449 NAND2X1_69/Y BUFX4_420/Y OAI21X1_1449/C gnd OAI21X1_1449/Y vdd OAI21X1
XFILL_37_9_0 gnd vdd FILL
XFILL_20_8_0 gnd vdd FILL
XFILL_3_9_0 gnd vdd FILL
XFILL_28_9_0 gnd vdd FILL
XFILL_11_8_0 gnd vdd FILL
XAOI21X1_70 BUFX4_381/Y MUX2X1_320/S AOI21X1_70/C gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_92 BUFX4_174/Y NOR2X1_155/B AOI21X1_92/C gnd AOI21X1_92/Y vdd AOI21X1
XAOI21X1_81 MUX2X1_86/B NOR2X1_137/B NOR2X1_138/Y gnd AOI21X1_81/Y vdd AOI21X1
XFILL_49_0_1 gnd vdd FILL
XBUFX4_301 BUFX4_302/A gnd BUFX4_301/Y vdd BUFX4
XBUFX4_312 INVX8_26/Y gnd BUFX4_312/Y vdd BUFX4
XBUFX4_334 BUFX4_28/Y gnd BUFX4_334/Y vdd BUFX4
XBUFX4_323 INVX8_1/Y gnd MUX2X1_8/B vdd BUFX4
XFILL_19_9_0 gnd vdd FILL
XBUFX4_345 BUFX4_27/Y gnd BUFX4_345/Y vdd BUFX4
XBUFX4_378 INVX8_14/Y gnd MUX2X1_82/B vdd BUFX4
XBUFX4_356 BUFX4_29/Y gnd BUFX4_356/Y vdd BUFX4
XNOR2X1_405 NOR2X1_405/A NOR2X1_405/B gnd NOR2X1_405/Y vdd NOR2X1
XNOR2X1_416 NOR2X1_416/A NOR2X1_416/B gnd NOR2X1_416/Y vdd NOR2X1
XBUFX4_389 BUFX4_384/A gnd BUFX4_389/Y vdd BUFX4
XBUFX4_367 BUFX4_30/Y gnd BUFX4_367/Y vdd BUFX4
XNOR2X1_449 NOR2X1_449/A AND2X2_41/A gnd NOR2X1_449/Y vdd NOR2X1
XNOR2X1_427 AND2X2_36/B NOR2X1_427/B gnd NOR2X1_427/Y vdd NOR2X1
XNOR2X1_438 NOR2X1_438/A AND2X2_47/B gnd NOR2X1_438/Y vdd NOR2X1
XFILL_19_3 gnd vdd FILL
XOAI21X1_1213 OAI21X1_158/C BUFX4_291/Y BUFX4_94/Y gnd OAI22X1_76/B vdd OAI21X1
XOAI21X1_1202 OAI21X1_238/C BUFX4_281/Y BUFX4_90/Y gnd OAI21X1_1203/B vdd OAI21X1
XOAI21X1_1224 BUFX4_363/Y NOR2X1_274/A BUFX4_157/Y gnd AOI21X1_501/C vdd OAI21X1
XOAI21X1_1235 BUFX4_343/Y NOR2X1_285/A BUFX4_159/Y gnd OAI22X1_84/C vdd OAI21X1
XDFFPOSX1_814 NOR2X1_591/A CLKBUF1_75/Y AOI21X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_803 OAI21X1_134/C CLKBUF1_55/Y OAI21X1_135/Y gnd vdd DFFPOSX1
XOAI21X1_1246 BUFX4_335/Y OAI21X1_278/C BUFX4_152/Y gnd OAI22X1_88/C vdd OAI21X1
XOAI21X1_1279 BUFX4_448/Y BUFX4_42/Y NOR2X1_522/B gnd OAI21X1_1279/Y vdd OAI21X1
XOAI21X1_1268 NAND2X1_30/Y BUFX4_426/Y OAI21X1_1268/C gnd DFFPOSX1_239/D vdd OAI21X1
XDFFPOSX1_847 NOR2X1_132/A CLKBUF1_69/Y AOI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_836 INVX1_94/A CLKBUF1_48/Y MUX2X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_825 NOR2X1_123/A CLKBUF1_42/Y AOI21X1_70/Y gnd vdd DFFPOSX1
XOAI21X1_1257 BUFX4_416/Y OAI22X1_92/Y AOI21X1_509/Y gnd NAND3X1_82/B vdd OAI21X1
XDFFPOSX1_858 NOR2X1_596/A CLKBUF1_62/Y AOI21X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_869 INVX1_106/A CLKBUF1_93/Y MUX2X1_93/Y gnd vdd DFFPOSX1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XAOI21X1_530 BUFX4_439/Y NOR2X1_85/B NOR2X1_642/Y gnd AOI21X1_530/Y vdd AOI21X1
XAOI21X1_552 BUFX4_428/Y MUX2X1_320/S NOR2X1_664/Y gnd AOI21X1_552/Y vdd AOI21X1
XAOI21X1_541 BUFX4_69/Y MUX2X1_75/S NOR2X1_653/Y gnd AOI21X1_541/Y vdd AOI21X1
XAOI21X1_574 BUFX4_317/Y NOR2X1_155/B NOR2X1_686/Y gnd AOI21X1_574/Y vdd AOI21X1
XAOI21X1_563 BUFX4_426/Y MUX2X1_89/S NOR2X1_675/Y gnd AOI21X1_563/Y vdd AOI21X1
XAOI21X1_585 BUFX4_420/Y MUX2X1_108/S NOR2X1_697/Y gnd AOI21X1_585/Y vdd AOI21X1
XAOI21X1_596 MUX2X1_27/B NOR2X1_707/B NOR2X1_708/Y gnd AOI21X1_596/Y vdd AOI21X1
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 INVX2_22/A XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XFILL_43_7_0 gnd vdd FILL
XMUX2X1_3 INVX1_6/Y BUFX4_71/Y MUX2X1_2/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 BUFX4_10/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XBUFX4_120 BUFX4_124/A gnd BUFX4_120/Y vdd BUFX4
XBUFX4_131 INVX8_20/Y gnd BUFX4_131/Y vdd BUFX4
XBUFX4_153 INVX8_32/Y gnd BUFX4_153/Y vdd BUFX4
XBUFX4_142 INVX8_7/Y gnd BUFX4_142/Y vdd BUFX4
XBUFX4_164 INVX8_24/Y gnd BUFX4_164/Y vdd BUFX4
XBUFX4_186 INVX8_19/Y gnd BUFX4_186/Y vdd BUFX4
XBUFX4_197 INVX8_27/Y gnd BUFX4_197/Y vdd BUFX4
XBUFX4_175 INVX8_13/Y gnd MUX2X1_40/B vdd BUFX4
XNOR2X1_224 NOR2X1_224/A NOR2X1_716/B gnd NOR2X1_224/Y vdd NOR2X1
XNOR2X1_202 INVX4_2/A BUFX4_161/Y gnd NOR2X1_707/B vdd NOR2X1
XNOR2X1_213 BUFX4_161/Y NOR2X1_39/B gnd MUX2X1_376/S vdd NOR2X1
XNOR2X1_235 NOR2X1_235/A NOR2X1_234/Y gnd NOR2X1_235/Y vdd NOR2X1
XNOR2X1_257 BUFX4_299/Y BUFX4_196/Y gnd MUX2X1_400/S vdd NOR2X1
XNOR2X1_246 NOR2X1_246/A NOR2X1_729/B gnd NOR2X1_246/Y vdd NOR2X1
XFILL_31_2 gnd vdd FILL
XFILL_34_7_0 gnd vdd FILL
XNOR2X1_279 NOR2X1_279/A AOI21X1_7/B gnd NOR2X1_279/Y vdd NOR2X1
XNOR2X1_268 NOR2X1_268/A NOR2X1_737/B gnd NOR2X1_268/Y vdd NOR2X1
XOAI21X1_708 OAI22X1_18/Y BUFX4_416/Y BUFX4_204/Y gnd AOI21X1_311/C vdd OAI21X1
XOAI21X1_719 BUFX4_358/Y OAI21X1_125/C BUFX4_158/Y gnd OAI22X1_19/C vdd OAI21X1
XOAI21X1_1021 BUFX4_363/Y NOR2X1_68/A BUFX4_157/Y gnd NOR2X1_500/B vdd OAI21X1
XOAI21X1_1010 NOR2X1_496/Y NOR2X1_497/Y BUFX4_394/Y gnd OAI21X1_1010/Y vdd OAI21X1
XDFFPOSX1_622 NAND2X1_14/A CLKBUF1_19/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_611 INVX1_18/A CLKBUF1_76/Y MUX2X1_13/Y gnd vdd DFFPOSX1
XOAI21X1_1054 INVX1_173/Y BUFX4_229/Y NAND2X1_321/Y gnd AOI21X1_453/B vdd OAI21X1
XDFFPOSX1_600 NAND2X1_6/A CLKBUF1_98/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XMUX2X1_219 MUX2X1_219/A MUX2X1_219/B BUFX4_99/Y gnd MUX2X1_219/Y vdd MUX2X1
XMUX2X1_208 MUX2X1_208/A MUX2X1_208/B BUFX4_99/Y gnd MUX2X1_208/Y vdd MUX2X1
XOAI21X1_1043 INVX1_401/Y BUFX4_291/Y AOI21X1_448/Y gnd OAI21X1_1045/C vdd OAI21X1
XOAI21X1_1032 BUFX4_353/Y NOR2X1_99/A BUFX4_158/Y gnd NOR2X1_502/B vdd OAI21X1
XDFFPOSX1_666 INVX1_37/A CLKBUF1_95/Y MUX2X1_29/Y gnd vdd DFFPOSX1
XOAI21X1_1076 INVX1_406/Y BUFX4_255/Y AOI21X1_458/Y gnd OAI21X1_1076/Y vdd OAI21X1
XOAI21X1_1087 AND2X2_23/A OAI21X1_1087/B AOI21X1_465/Y gnd OAI21X1_1087/Y vdd OAI21X1
XDFFPOSX1_644 NOR2X1_29/A CLKBUF1_103/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_633 INVX1_30/A CLKBUF1_73/Y MUX2X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_655 OAI21X1_35/C CLKBUF1_51/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XOAI21X1_1065 INVX1_405/Y BUFX4_242/Y AOI21X1_455/Y gnd OAI21X1_1065/Y vdd OAI21X1
XOAI21X1_1098 BUFX4_353/Y DFFPOSX1_185/Q BUFX4_158/Y gnd OAI22X1_51/C vdd OAI21X1
XDFFPOSX1_699 NOR2X1_403/A CLKBUF1_80/Y OAI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_688 INVX1_41/A CLKBUF1_70/Y MUX2X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_677 NOR2X1_47/A CLKBUF1_100/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XFILL_0_7_0 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XAOI21X1_360 INVX1_45/Y BUFX4_252/Y OAI21X1_824/Y gnd AOI21X1_360/Y vdd AOI21X1
XAOI21X1_393 BUFX4_31/Y MUX2X1_229/Y BUFX4_392/Y gnd AOI21X1_393/Y vdd AOI21X1
XAOI21X1_371 INVX1_335/Y BUFX4_270/Y OAI21X1_844/Y gnd AOI21X1_371/Y vdd AOI21X1
XAOI21X1_382 AOI21X1_382/A BUFX4_338/Y AND2X2_36/Y gnd OAI21X1_873/B vdd AOI21X1
XDFFPOSX1_81 NOR2X1_278/A CLKBUF1_21/Y DFFPOSX1_81/D gnd vdd DFFPOSX1
XDFFPOSX1_70 NAND2X1_94/A CLKBUF1_76/Y OAI21X1_376/Y gnd vdd DFFPOSX1
XDFFPOSX1_92 NOR2X1_505/A CLKBUF1_28/Y DFFPOSX1_92/D gnd vdd DFFPOSX1
XFILL_8_8_0 gnd vdd FILL
XBUFX4_15 address[1] gnd BUFX4_85/A vdd BUFX4
XBUFX4_26 BUFX4_28/A gnd BUFX4_26/Y vdd BUFX4
XBUFX4_59 INVX8_6/Y gnd BUFX4_59/Y vdd BUFX4
XBUFX4_48 address[4] gnd BUFX4_48/Y vdd BUFX4
XBUFX4_37 BUFX4_33/A gnd BUFX4_37/Y vdd BUFX4
XFILL_16_7_0 gnd vdd FILL
XINVX8_18 INVX8_18/A gnd INVX8_18/Y vdd INVX8
XINVX8_29 INVX8_29/A gnd INVX8_29/Y vdd INVX8
XOAI21X1_505 INVX4_12/A AOI22X1_6/B AOI22X1_6/A gnd INVX1_207/A vdd OAI21X1
XOAI21X1_538 INVX2_17/Y BUFX4_306/Y OAI21X1_538/C gnd AND2X2_15/A vdd OAI21X1
XOAI21X1_516 AND2X2_2/Y NOR2X1_301/Y INVX1_209/Y gnd OR2X2_6/A vdd OAI21X1
XOAI21X1_527 NOR2X1_336/B INVX4_10/A INVX4_12/Y gnd NAND3X1_63/C vdd OAI21X1
XOAI21X1_549 BUFX4_189/Y INVX4_1/Y INVX1_27/A gnd OAI21X1_550/C vdd OAI21X1
XDFFPOSX1_430 BUFX2_7/A CLKBUF1_96/Y OAI21X1_1084/Y gnd vdd DFFPOSX1
XDFFPOSX1_463 NOR2X1_707/A CLKBUF1_102/Y AOI21X1_595/Y gnd vdd DFFPOSX1
XDFFPOSX1_441 INVX1_361/A CLKBUF1_70/Y MUX2X1_271/Y gnd vdd DFFPOSX1
XDFFPOSX1_474 INVX1_435/A CLKBUF1_22/Y MUX2X1_374/Y gnd vdd DFFPOSX1
XDFFPOSX1_452 NOR2X1_704/A CLKBUF1_1/Y AOI21X1_592/Y gnd vdd DFFPOSX1
XDFFPOSX1_496 NOR2X1_435/B CLKBUF1_79/Y DFFPOSX1_496/D gnd vdd DFFPOSX1
XDFFPOSX1_485 AOI21X1_414/B CLKBUF1_89/Y DFFPOSX1_485/D gnd vdd DFFPOSX1
XFILL_40_5_0 gnd vdd FILL
XAOI21X1_190 BUFX4_173/Y NOR2X1_33/Y NOR2X1_287/Y gnd AOI21X1_190/Y vdd AOI21X1
XFILL_48_6_0 gnd vdd FILL
XFILL_31_5_0 gnd vdd FILL
XFILL_39_6_0 gnd vdd FILL
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_313 NAND2X1_78/Y BUFX4_218/Y OAI21X1_313/C gnd OAI21X1_313/Y vdd OAI21X1
XOAI21X1_302 NOR2X1_77/B BUFX4_457/Y OAI21X1_302/C gnd OAI21X1_303/C vdd OAI21X1
XOAI21X1_335 NAND2X1_80/Y BUFX4_467/Y OAI21X1_335/C gnd OAI21X1_335/Y vdd OAI21X1
XOAI21X1_346 INVX4_3/A BUFX4_199/Y OAI21X1_876/A gnd OAI21X1_347/C vdd OAI21X1
XOAI21X1_324 BUFX4_389/Y BUFX4_313/Y INVX1_408/A gnd OAI21X1_325/C vdd OAI21X1
XOAI21X1_357 NAND2X1_84/Y BUFX4_372/Y OAI21X1_356/Y gnd OAI21X1_357/Y vdd OAI21X1
XOAI21X1_379 BUFX4_473/Y OAI21X1_7/B NAND2X1_97/Y gnd DFFPOSX1_73/D vdd OAI21X1
XOAI21X1_368 BUFX4_209/Y NAND2X1_2/Y NAND2X1_86/Y gnd DFFPOSX1_42/D vdd OAI21X1
XDFFPOSX1_282 OAI21X1_599/B CLKBUF1_9/Y DFFPOSX1_282/D gnd vdd DFFPOSX1
XDFFPOSX1_260 INVX1_354/A CLKBUF1_93/Y MUX2X1_333/Y gnd vdd DFFPOSX1
XDFFPOSX1_271 OAI21X1_765/B CLKBUF1_5/Y OAI21X1_1377/Y gnd vdd DFFPOSX1
XDFFPOSX1_293 OAI21X1_1452/C CLKBUF1_10/Y DFFPOSX1_293/D gnd vdd DFFPOSX1
XNAND2X1_330 NOR2X1_237/A BUFX4_251/Y gnd NAND2X1_330/Y vdd NAND2X1
XNAND2X1_363 NAND2X1_363/A NAND2X1_2/Y gnd NAND2X1_363/Y vdd NAND2X1
XNAND2X1_352 NOR2X1_249/A BUFX4_257/Y gnd NAND2X1_352/Y vdd NAND2X1
XNAND2X1_341 INVX8_33/Y OAI22X1_66/Y gnd NAND2X1_341/Y vdd NAND2X1
XFILL_5_6_0 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XOAI21X1_880 INVX1_164/Y AND2X2_46/B NAND2X1_264/Y gnd MUX2X1_225/B vdd OAI21X1
XOAI21X1_891 BUFX4_32/Y MUX2X1_226/Y AOI21X1_389/Y gnd NAND3X1_75/C vdd OAI21X1
XMUX2X1_391 AND2X2_6/B INVX1_440/Y NOR2X1_727/B gnd MUX2X1_391/Y vdd MUX2X1
XMUX2X1_380 BUFX4_324/Y INVX1_432/Y NOR2X1_220/B gnd MUX2X1_380/Y vdd MUX2X1
XNAND3X1_3 NOR2X1_2/A INVX1_14/A NOR2X1_6/Y gnd MUX2X1_14/S vdd NAND3X1
XOAI21X1_121 INVX4_4/A BUFX4_52/Y NOR2X1_501/A gnd OAI21X1_122/C vdd OAI21X1
XOAI21X1_110 MUX2X1_59/B NAND2X1_39/Y OAI21X1_110/C gnd OAI21X1_110/Y vdd OAI21X1
XAOI22X1_8 AOI22X1_8/A AOI22X1_8/B AOI22X1_8/C INVX4_9/A gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_165 NAND2X1_53/Y BUFX4_381/Y OAI21X1_164/Y gnd OAI21X1_165/Y vdd OAI21X1
XOAI21X1_154 NOR2X1_77/B BUFX4_183/Y AND2X2_34/B gnd OAI21X1_155/C vdd OAI21X1
XOAI21X1_143 INVX1_92/Y NAND2X1_50/B NAND2X1_50/Y gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_132 MUX2X1_58/A NAND2X1_44/Y OAI21X1_132/C gnd OAI21X1_132/Y vdd OAI21X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XOAI21X1_176 BUFX4_385/Y BUFX4_131/Y OAI21X1_686/A gnd OAI21X1_177/C vdd OAI21X1
XOAI21X1_187 MUX2X1_49/A NAND2X1_58/Y OAI21X1_186/Y gnd OAI21X1_187/Y vdd OAI21X1
XOAI21X1_198 BUFX4_387/Y BUFX4_406/Y OAI21X1_198/C gnd OAI21X1_198/Y vdd OAI21X1
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XNAND2X1_18 NOR2X1_4/Y NOR2X1_8/Y gnd BUFX4_384/A vdd NAND2X1
XNAND2X1_171 BUFX4_393/Y AOI22X1_11/Y gnd AOI22X1_14/B vdd NAND2X1
XNAND2X1_29 INVX8_10/A INVX8_9/A gnd OAI21X1_64/B vdd NAND2X1
XNAND2X1_160 NAND2X1_160/A NOR3X1_7/Y gnd XNOR2X1_5/B vdd NAND2X1
XNAND2X1_193 NOR2X1_34/A BUFX4_223/Y gnd NAND2X1_193/Y vdd NAND2X1
XNAND2X1_182 BUFX4_101/Y NOR2X1_728/A gnd OAI21X1_605/C vdd NAND2X1
XFILL_46_9_1 gnd vdd FILL
XFILL_45_4_0 gnd vdd FILL
XNOR2X1_609 BUFX4_412/Y NOR2X1_609/B gnd OAI22X1_86/C vdd NOR2X1
XAOI22X1_27 AOI22X1_27/A NOR2X1_488/Y AOI22X1_27/C BUFX4_207/Y gnd AOI22X1_27/Y vdd
+ AOI22X1
XAOI22X1_16 AOI22X1_16/A AOI22X1_16/B AOI22X1_16/C BUFX4_204/Y gnd MUX2X1_190/B vdd
+ AOI22X1
XOAI21X1_1428 BUFX4_383/Y BUFX4_141/Y AOI21X1_472/A gnd OAI21X1_1428/Y vdd OAI21X1
XOAI21X1_1417 NAND2X1_62/Y BUFX4_422/Y OAI21X1_1417/C gnd DFFPOSX1_415/D vdd OAI21X1
XOAI21X1_1406 BUFX4_452/Y BUFX4_407/Y NOR2X1_370/B gnd OAI21X1_1407/C vdd OAI21X1
XOAI21X1_1439 BUFX4_444/Y NAND2X1_68/Y OAI21X1_1439/C gnd DFFPOSX1_282/D vdd OAI21X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XFILL_37_9_1 gnd vdd FILL
XFILL_36_4_0 gnd vdd FILL
XFILL_20_8_1 gnd vdd FILL
XFILL_3_9_1 gnd vdd FILL
XFILL_28_9_1 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XFILL_27_4_0 gnd vdd FILL
XFILL_11_8_1 gnd vdd FILL
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_71 MUX2X1_83/B MUX2X1_320/S AOI21X1_71/C gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_60 BUFX4_371/Y NOR2X1_107/B NOR2X1_108/Y gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_82 MUX2X1_83/B NOR2X1_137/B AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XAOI21X1_93 BUFX4_380/Y NOR2X1_155/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XBUFX4_313 INVX8_26/Y gnd BUFX4_313/Y vdd BUFX4
XBUFX4_302 BUFX4_302/A gnd INVX4_2/A vdd BUFX4
XBUFX4_346 BUFX4_28/Y gnd BUFX4_346/Y vdd BUFX4
XFILL_19_9_1 gnd vdd FILL
XBUFX4_324 INVX8_1/Y gnd BUFX4_324/Y vdd BUFX4
XBUFX4_335 BUFX4_27/Y gnd BUFX4_335/Y vdd BUFX4
XBUFX4_368 BUFX4_25/Y gnd BUFX4_368/Y vdd BUFX4
XBUFX4_379 INVX8_14/Y gnd MUX2X1_86/B vdd BUFX4
XFILL_18_4_0 gnd vdd FILL
XBUFX4_357 BUFX4_27/Y gnd BUFX4_357/Y vdd BUFX4
XNOR2X1_406 NOR2X1_75/A BUFX4_234/Y gnd OAI22X1_18/D vdd NOR2X1
XNOR2X1_417 BUFX4_111/Y NOR2X1_417/B gnd NOR2X1_418/A vdd NOR2X1
XNOR2X1_439 BUFX4_410/Y NOR2X1_439/B gnd OAI22X1_24/A vdd NOR2X1
XNOR2X1_428 BUFX4_220/Y NOR2X1_428/B gnd OAI22X1_22/D vdd NOR2X1
XOAI22X1_90 NOR2X1_620/Y OAI22X1_90/B OAI22X1_90/C NOR2X1_619/Y gnd MUX2X1_264/A vdd
+ OAI22X1
XOAI21X1_1203 NOR2X1_583/Y OAI21X1_1203/B OAI21X1_1203/C gnd NOR2X1_584/B vdd OAI21X1
XOAI21X1_1214 BUFX4_325/Y NOR2X1_129/A BUFX4_150/Y gnd OAI22X1_77/C vdd OAI21X1
XOAI21X1_1236 OAI21X1_403/C BUFX4_235/Y BUFX4_103/Y gnd OAI22X1_84/B vdd OAI21X1
XOAI21X1_1225 DFFPOSX1_37/Q BUFX4_227/Y BUFX4_99/Y gnd AOI21X1_502/C vdd OAI21X1
XDFFPOSX1_815 OAI21X1_677/B CLKBUF1_16/Y OAI21X1_145/Y gnd vdd DFFPOSX1
XDFFPOSX1_804 INVX1_334/A CLKBUF1_20/Y OAI21X1_137/Y gnd vdd DFFPOSX1
XOAI21X1_1247 NOR2X1_220/A BUFX4_242/Y BUFX4_106/Y gnd OAI22X1_88/B vdd OAI21X1
XDFFPOSX1_848 INVX1_101/A CLKBUF1_53/Y MUX2X1_88/Y gnd vdd DFFPOSX1
XOAI21X1_1269 BUFX4_299/Y BUFX4_42/Y OAI21X1_935/B gnd OAI21X1_1270/C vdd OAI21X1
XOAI21X1_1258 INVX1_444/Y AND2X2_27/A NAND2X1_350/Y gnd MUX2X1_266/B vdd OAI21X1
XDFFPOSX1_837 INVX1_95/A CLKBUF1_32/Y MUX2X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_826 NOR2X1_124/A CLKBUF1_75/Y AOI21X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_859 INVX1_102/A CLKBUF1_31/Y MUX2X1_89/Y gnd vdd DFFPOSX1
XAOI21X1_520 MUX2X1_1/B NOR2X1_65/Y NOR2X1_632/Y gnd AOI21X1_520/Y vdd AOI21X1
XAOI21X1_531 BUFX4_424/Y MUX2X1_50/S NOR2X1_643/Y gnd AOI21X1_531/Y vdd AOI21X1
XAOI21X1_553 BUFX4_318/Y MUX2X1_320/S NOR2X1_665/Y gnd AOI21X1_553/Y vdd AOI21X1
XAOI21X1_542 BUFX4_316/Y MUX2X1_75/S NOR2X1_654/Y gnd AOI21X1_542/Y vdd AOI21X1
XAOI21X1_586 BUFX4_437/Y INVX1_219/A NOR2X1_698/Y gnd AOI21X1_586/Y vdd AOI21X1
XAOI21X1_564 BUFX4_321/Y MUX2X1_89/S NOR2X1_676/Y gnd AOI21X1_564/Y vdd AOI21X1
XAOI21X1_575 BUFX4_422/Y MUX2X1_340/S NOR2X1_687/Y gnd AOI21X1_575/Y vdd AOI21X1
XAOI21X1_597 BUFX4_70/Y NOR2X1_707/B NOR2X1_709/Y gnd AOI21X1_597/Y vdd AOI21X1
XXOR2X1_3 XOR2X1_3/A INVX2_22/A gnd XOR2X1_3/Y vdd XOR2X1
XFILL_43_7_1 gnd vdd FILL
XMUX2X1_4 INVX1_7/Y MUX2X1_4/B MUX2X1_2/S gnd MUX2X1_4/Y vdd MUX2X1
XFILL_42_2_0 gnd vdd FILL
XCLKBUF1_5 BUFX4_1/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_110 BUFX4_14/Y gnd BUFX4_110/Y vdd BUFX4
XBUFX4_121 BUFX4_124/A gnd BUFX4_121/Y vdd BUFX4
XBUFX4_154 INVX8_32/Y gnd BUFX4_154/Y vdd BUFX4
XBUFX4_132 INVX8_8/Y gnd BUFX4_132/Y vdd BUFX4
XBUFX4_143 INVX8_7/Y gnd BUFX4_143/Y vdd BUFX4
XBUFX4_187 INVX8_19/Y gnd BUFX4_187/Y vdd BUFX4
XBUFX4_165 INVX8_29/Y gnd BUFX4_165/Y vdd BUFX4
XNOR2X1_225 NOR2X1_516/A NOR2X1_716/B gnd NOR2X1_225/Y vdd NOR2X1
XBUFX4_176 INVX8_13/Y gnd BUFX4_176/Y vdd BUFX4
XNOR2X1_203 NOR2X1_466/A NOR2X1_707/B gnd NOR2X1_203/Y vdd NOR2X1
XNOR2X1_214 NOR2X1_214/A MUX2X1_376/S gnd NOR2X1_214/Y vdd NOR2X1
XNOR2X1_236 NOR2X1_236/A NOR2X1_234/Y gnd NOR2X1_236/Y vdd NOR2X1
XBUFX4_198 INVX8_27/Y gnd BUFX4_198/Y vdd BUFX4
XNOR2X1_258 NOR2X1_453/A MUX2X1_400/S gnd NOR2X1_258/Y vdd NOR2X1
XNOR2X1_247 NOR2X1_247/A NOR2X1_729/B gnd NOR2X1_247/Y vdd NOR2X1
XFILL_31_3 gnd vdd FILL
XFILL_34_7_1 gnd vdd FILL
XNOR2X1_269 NOR2X1_269/A NOR2X1_737/B gnd NOR2X1_269/Y vdd NOR2X1
XFILL_33_2_0 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XOAI21X1_709 AOI21X1_311/Y NOR2X1_405/Y BUFX4_390/Y gnd OAI21X1_709/Y vdd OAI21X1
XOAI21X1_1022 OAI21X1_87/C BUFX4_270/Y BUFX4_104/Y gnd AOI21X1_439/C vdd OAI21X1
XOAI21X1_1000 OAI21X1_999/Y AND2X2_43/Y BUFX4_416/Y gnd OAI22X1_43/D vdd OAI21X1
XOAI21X1_1011 INVX1_397/Y BUFX4_419/Y NAND2X1_307/Y gnd AOI21X1_434/B vdd OAI21X1
XOAI21X1_1055 AOI21X1_453/Y BUFX4_36/Y OAI21X1_1055/C gnd MUX2X1_253/A vdd OAI21X1
XDFFPOSX1_623 INVX1_272/A CLKBUF1_81/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_601 NAND2X1_7/A CLKBUF1_73/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_612 INVX1_19/A CLKBUF1_98/Y MUX2X1_14/Y gnd vdd DFFPOSX1
XMUX2X1_209 MUX2X1_209/A MUX2X1_208/Y BUFX4_419/Y gnd AOI22X1_19/C vdd MUX2X1
XOAI21X1_1044 INVX1_186/Y BUFX4_220/Y BUFX4_114/Y gnd OAI21X1_1044/Y vdd OAI21X1
XOAI21X1_1033 INVX1_71/A AND2X2_41/A BUFX4_109/Y gnd AOI21X1_444/C vdd OAI21X1
XOAI21X1_1077 INVX1_147/Y BUFX4_257/Y BUFX4_84/Y gnd OAI21X1_1077/Y vdd OAI21X1
XOAI21X1_1088 BUFX4_265/Y NOR2X1_628/A BUFX4_87/Y gnd OAI21X1_1089/B vdd OAI21X1
XDFFPOSX1_634 INVX1_31/A CLKBUF1_30/Y MUX2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_645 NOR2X1_30/A CLKBUF1_66/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XOAI21X1_1066 INVX1_136/Y BUFX4_244/Y BUFX4_78/Y gnd OAI21X1_1067/A vdd OAI21X1
XDFFPOSX1_656 NOR2X1_438/A CLKBUF1_63/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_689 INVX1_42/A CLKBUF1_70/Y MUX2X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_678 NOR2X1_48/A CLKBUF1_87/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_667 NOR2X1_40/A CLKBUF1_77/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XOAI21X1_1099 BUFX4_273/Y NOR2X1_645/A BUFX4_95/Y gnd OAI22X1_51/B vdd OAI21X1
XINVX1_390 INVX1_390/A gnd INVX1_390/Y vdd INVX1
XFILL_0_7_1 gnd vdd FILL
XFILL_25_7_1 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 INVX8_7/A gnd INVX8_7/Y vdd INVX8
XAOI21X1_350 BUFX4_146/Y INVX1_329/Y OAI21X1_797/Y gnd AOI21X1_350/Y vdd AOI21X1
XAOI21X1_361 NOR2X1_81/A BUFX4_93/Y OAI21X1_827/Y gnd OAI22X1_25/B vdd AOI21X1
XAOI21X1_383 INVX1_181/Y BUFX4_355/Y BUFX4_156/Y gnd OAI21X1_872/C vdd AOI21X1
XAOI21X1_394 NOR2X1_638/A BUFX4_365/Y BUFX4_87/Y gnd OAI21X1_915/C vdd AOI21X1
XAOI21X1_372 BUFX4_152/Y AOI21X1_372/B AOI21X1_371/Y gnd OAI21X1_847/B vdd AOI21X1
XDFFPOSX1_60 INVX1_165/A CLKBUF1_30/Y MUX2X1_152/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 NAND2X1_95/A CLKBUF1_73/Y DFFPOSX1_71/D gnd vdd DFFPOSX1
XDFFPOSX1_93 NOR2X1_606/A CLKBUF1_84/Y DFFPOSX1_93/D gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_175/A CLKBUF1_66/Y MUX2X1_162/Y gnd vdd DFFPOSX1
XFILL_8_8_1 gnd vdd FILL
XFILL_7_3_0 gnd vdd FILL
XBUFX4_16 address[1] gnd BUFX4_75/A vdd BUFX4
XBUFX4_49 address[4] gnd BUFX4_49/Y vdd BUFX4
XBUFX4_27 BUFX4_28/A gnd BUFX4_27/Y vdd BUFX4
XBUFX4_38 BUFX4_33/A gnd BUFX4_38/Y vdd BUFX4
XFILL_16_7_1 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XINVX8_19 INVX8_19/A gnd INVX8_19/Y vdd INVX8
XOAI21X1_506 OAI21X1_506/A NOR2X1_334/A INVX1_207/A gnd NAND3X1_58/C vdd OAI21X1
XOAI21X1_517 INVX1_209/A INVX2_24/Y XNOR2X1_4/B gnd AND2X2_12/A vdd OAI21X1
XOAI21X1_528 OAI21X1_528/A NOR2X1_338/Y NAND3X1_63/Y gnd OAI21X1_528/Y vdd OAI21X1
XOAI21X1_539 OR2X2_4/Y traffic_Street_0[2] traffic_Street_0[3] gnd OAI21X1_539/Y vdd
+ OAI21X1
XDFFPOSX1_431 BUFX2_8/A CLKBUF1_100/Y AOI21X1_512/Y gnd vdd DFFPOSX1
XDFFPOSX1_420 INVX1_192/A CLKBUF1_71/Y OAI21X1_546/Y gnd vdd DFFPOSX1
XDFFPOSX1_453 NOR2X1_705/A CLKBUF1_82/Y AOI21X1_593/Y gnd vdd DFFPOSX1
XDFFPOSX1_464 NOR2X1_428/B CLKBUF1_1/Y AOI21X1_596/Y gnd vdd DFFPOSX1
XDFFPOSX1_442 NOR2X1_521/A CLKBUF1_43/Y AOI21X1_519/Y gnd vdd DFFPOSX1
XDFFPOSX1_475 INVX1_255/A CLKBUF1_95/Y MUX2X1_375/Y gnd vdd DFFPOSX1
XDFFPOSX1_497 NOR2X1_485/B CLKBUF1_79/Y OAI21X1_1494/Y gnd vdd DFFPOSX1
XDFFPOSX1_486 AOI21X1_487/B CLKBUF1_68/Y OAI21X1_1480/Y gnd vdd DFFPOSX1
XFILL_40_5_1 gnd vdd FILL
XAOI21X1_180 BUFX4_375/Y NOR2X1_16/Y NOR2X1_277/Y gnd DFFPOSX1_80/D vdd AOI21X1
XAOI21X1_191 BUFX4_375/Y NOR2X1_33/Y NOR2X1_288/Y gnd AOI21X1_191/Y vdd AOI21X1
XFILL_48_6_1 gnd vdd FILL
XFILL_47_1_0 gnd vdd FILL
XFILL_31_5_1 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XFILL_39_6_1 gnd vdd FILL
XFILL_38_1_0 gnd vdd FILL
XFILL_22_5_1 gnd vdd FILL
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_314 BUFX4_313/Y BUFX4_300/Y INVX1_341/A gnd OAI21X1_314/Y vdd OAI21X1
XOAI21X1_303 NAND2X1_76/Y BUFX4_469/Y OAI21X1_303/C gnd OAI21X1_303/Y vdd OAI21X1
XOAI21X1_336 BUFX4_194/Y BUFX4_309/Y DFFPOSX1_6/Q gnd OAI21X1_337/C vdd OAI21X1
XOAI21X1_347 NAND2X1_82/Y MUX2X1_40/B OAI21X1_347/C gnd DFFPOSX1_19/D vdd OAI21X1
XOAI21X1_325 NAND2X1_79/Y BUFX4_380/Y OAI21X1_325/C gnd OAI21X1_325/Y vdd OAI21X1
XOAI21X1_369 BUFX4_173/Y NAND2X1_2/Y NAND2X1_87/Y gnd DFFPOSX1_43/D vdd OAI21X1
XOAI21X1_358 INVX4_5/A BUFX4_197/Y DFFPOSX1_37/Q gnd OAI21X1_359/C vdd OAI21X1
XBUFX4_1 clock gnd BUFX4_1/Y vdd BUFX4
XDFFPOSX1_250 INVX1_239/A CLKBUF1_41/Y MUX2X1_354/Y gnd vdd DFFPOSX1
XDFFPOSX1_261 NOR2X1_676/A CLKBUF1_62/Y AOI21X1_564/Y gnd vdd DFFPOSX1
XDFFPOSX1_272 INVX1_351/A CLKBUF1_26/Y DFFPOSX1_272/D gnd vdd DFFPOSX1
XDFFPOSX1_283 NAND2X1_239/B CLKBUF1_82/Y OAI21X1_1441/Y gnd vdd DFFPOSX1
XDFFPOSX1_294 INVX1_455/A CLKBUF1_34/Y MUX2X1_325/Y gnd vdd DFFPOSX1
XNAND2X1_320 BUFX4_37/Y NOR2X1_508/Y gnd NAND2X1_320/Y vdd NAND2X1
XNAND2X1_331 BUFX4_32/Y NOR2X1_520/Y gnd NAND2X1_331/Y vdd NAND2X1
XNAND2X1_342 BUFX4_205/Y NAND2X1_342/B gnd OAI22X1_69/C vdd NAND2X1
XNAND2X1_353 traffic_Street_0[1] NOR2X1_76/B gnd NAND2X1_353/Y vdd NAND2X1
XFILL_5_6_1 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XFILL_29_1_0 gnd vdd FILL
XFILL_13_5_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XOAI21X1_892 INVX1_138/Y BUFX4_232/Y NAND2X1_268/Y gnd MUX2X1_227/B vdd OAI21X1
XOAI21X1_881 INVX1_172/Y INVX8_31/A NAND2X1_265/Y gnd MUX2X1_225/A vdd OAI21X1
XOAI21X1_870 INVX1_338/Y BUFX4_283/Y OAI21X1_870/C gnd MUX2X1_224/B vdd OAI21X1
XMUX2X1_370 BUFX4_70/Y INVX1_376/Y MUX2X1_369/S gnd MUX2X1_370/Y vdd MUX2X1
XMUX2X1_381 BUFX4_439/Y INVX1_266/Y NOR2X1_232/Y gnd MUX2X1_381/Y vdd MUX2X1
XMUX2X1_392 BUFX4_429/Y INVX1_325/Y NOR2X1_729/B gnd MUX2X1_392/Y vdd MUX2X1
XNAND3X1_4 NOR2X1_2/A INVX1_23/A NOR2X1_6/Y gnd OAI21X1_7/B vdd NAND3X1
XOAI21X1_100 NAND2X1_36/Y BUFX4_469/Y OAI21X1_99/Y gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_111 BUFX4_56/Y BUFX4_53/Y OAI21X1_111/C gnd OAI21X1_112/C vdd OAI21X1
XOAI21X1_122 NAND2X1_40/Y BUFX4_371/Y OAI21X1_122/C gnd OAI21X1_122/Y vdd OAI21X1
XAOI22X1_9 OR2X2_2/A XNOR2X1_4/A AOI22X1_9/C AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_155 NAND2X1_52/Y BUFX4_176/Y OAI21X1_155/C gnd OAI21X1_155/Y vdd OAI21X1
XOAI21X1_144 BUFX4_59/Y BUFX4_184/Y OAI21X1_677/B gnd OAI21X1_144/Y vdd OAI21X1
XOAI21X1_133 INVX1_90/Y NOR2X1_107/B NAND2X1_47/Y gnd OAI21X1_133/Y vdd OAI21X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XOAI21X1_166 BUFX4_454/Y BUFX4_186/Y NOR2X1_593/A gnd OAI21X1_167/C vdd OAI21X1
XOAI21X1_177 NAND2X1_57/Y BUFX4_214/Y OAI21X1_177/C gnd OAI21X1_177/Y vdd OAI21X1
XOAI21X1_188 BUFX4_136/Y BUFX4_127/Y NAND2X1_301/A gnd OAI21X1_188/Y vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XOAI21X1_199 NAND2X1_59/Y BUFX4_465/Y OAI21X1_198/Y gnd OAI21X1_199/Y vdd OAI21X1
XNAND2X1_150 NAND3X1_56/A XNOR2X1_4/Y gnd NOR2X1_334/B vdd NAND2X1
XNAND2X1_161 NAND2X1_161/A INVX2_26/Y gnd XNOR2X1_6/B vdd NAND2X1
XNAND2X1_19 INVX8_5/A INVX4_3/Y gnd MUX2X1_21/S vdd NAND2X1
XNAND2X1_183 BUFX4_273/Y NOR2X1_730/A gnd NAND2X1_183/Y vdd NAND2X1
XNAND2X1_194 NOR2X1_45/A BUFX4_225/Y gnd OAI21X1_629/C vdd NAND2X1
XNAND2X1_172 BUFX4_229/Y NAND2X1_172/B gnd OAI21X1_563/C vdd NAND2X1
XFILL_45_4_1 gnd vdd FILL
XAOI22X1_28 AOI22X1_28/A AOI22X1_28/B AOI22X1_28/C BUFX4_401/Y gnd OAI22X1_42/C vdd
+ AOI22X1
XAOI22X1_17 AOI22X1_17/A AOI22X1_17/B MUX2X1_190/Y BUFX4_402/Y gnd AOI22X1_17/Y vdd
+ AOI22X1
XOAI21X1_1429 NAND2X1_64/Y BUFX4_317/Y OAI21X1_1428/Y gnd DFFPOSX1_213/D vdd OAI21X1
XOAI21X1_1407 NAND2X1_61/Y AND2X2_5/B OAI21X1_1407/C gnd DFFPOSX1_174/D vdd OAI21X1
XOAI21X1_1418 BUFX4_119/Y BUFX4_406/Y MUX2X1_230/A gnd OAI21X1_1419/C vdd OAI21X1
XNOR3X1_7 NOR3X1_3/Y OR2X2_5/Y NOR3X1_6/Y gnd NOR3X1_7/Y vdd NOR3X1
XFILL_5_1 gnd vdd FILL
XFILL_47_1 gnd vdd FILL
XFILL_36_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_27_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_61 BUFX4_470/Y NOR2X1_107/B NOR2X1_109/Y gnd AOI21X1_61/Y vdd AOI21X1
XAOI21X1_50 MUX2X1_44/A NOR2X1_92/B NOR2X1_94/Y gnd AOI21X1_50/Y vdd AOI21X1
XAOI21X1_83 BUFX4_467/Y MUX2X1_89/S NOR2X1_141/Y gnd AOI21X1_83/Y vdd AOI21X1
XAOI21X1_72 BUFX4_218/Y AOI21X1_72/B NOR2X1_126/Y gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_94 BUFX4_465/Y NOR2X1_155/B AOI21X1_94/C gnd AOI21X1_94/Y vdd AOI21X1
XOAI21X1_1 MUX2X1_8/B NAND2X1_2/Y NAND2X1_3/Y gnd OAI21X1_1/Y vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XBUFX4_303 BUFX4_302/A gnd BUFX4_303/Y vdd BUFX4
XBUFX4_325 BUFX4_29/Y gnd BUFX4_325/Y vdd BUFX4
XBUFX4_314 INVX8_1/Y gnd MUX2X1_4/B vdd BUFX4
XBUFX4_336 BUFX4_27/Y gnd BUFX4_336/Y vdd BUFX4
XBUFX4_369 BUFX4_30/Y gnd BUFX4_369/Y vdd BUFX4
XFILL_18_4_1 gnd vdd FILL
XBUFX4_347 BUFX4_26/Y gnd BUFX4_347/Y vdd BUFX4
XNOR2X1_407 NOR2X1_80/A BUFX4_366/Y gnd OAI22X1_18/A vdd NOR2X1
XBUFX4_358 BUFX4_26/Y gnd BUFX4_358/Y vdd BUFX4
XNOR2X1_418 NOR2X1_418/A NOR2X1_418/B gnd NOR2X1_419/B vdd NOR2X1
XNOR2X1_429 NOR2X1_713/A BUFX4_341/Y gnd NOR2X1_429/Y vdd NOR2X1
XOAI22X1_80 OAI22X1_80/A OAI22X1_80/B OAI22X1_80/C BUFX4_202/Y gnd OAI22X1_80/Y vdd
+ OAI22X1
XOAI22X1_91 OAI22X1_91/A OAI22X1_91/B OAI22X1_91/C INVX8_29/A gnd OAI22X1_91/Y vdd
+ OAI22X1
XOAI21X1_1204 BUFX4_335/Y NOR2X1_157/A BUFX4_152/Y gnd OAI22X1_73/C vdd OAI21X1
XOAI21X1_1215 INVX1_96/A BUFX4_220/Y BUFX4_95/Y gnd OAI22X1_77/B vdd OAI21X1
XOAI21X1_1226 AOI21X1_501/Y AOI21X1_502/Y INVX8_30/A gnd AOI21X1_503/B vdd OAI21X1
XDFFPOSX1_805 INVX1_400/A CLKBUF1_20/Y OAI21X1_139/Y gnd vdd DFFPOSX1
XOAI21X1_1237 BUFX4_338/Y OAI21X1_419/C BUFX4_156/Y gnd OAI21X1_1239/B vdd OAI21X1
XOAI21X1_1259 INVX1_148/Y BUFX4_256/Y NAND2X1_351/Y gnd MUX2X1_266/A vdd OAI21X1
XDFFPOSX1_827 OAI21X1_160/C CLKBUF1_48/Y OAI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_838 INVX1_96/A CLKBUF1_85/Y MUX2X1_83/Y gnd vdd DFFPOSX1
XDFFPOSX1_816 INVX1_336/A CLKBUF1_75/Y OAI21X1_147/Y gnd vdd DFFPOSX1
XOAI21X1_1248 OAI22X1_88/Y BUFX4_35/Y BUFX4_207/Y gnd OAI22X1_91/A vdd OAI21X1
XDFFPOSX1_849 AND2X2_44/A CLKBUF1_62/Y AOI21X1_77/Y gnd vdd DFFPOSX1
XAOI21X1_510 AOI21X1_510/A BUFX4_336/Y BUFX4_155/Y gnd AOI21X1_510/Y vdd AOI21X1
XAOI21X1_521 BUFX4_421/Y NOR2X1_65/Y NOR2X1_633/Y gnd AOI21X1_521/Y vdd AOI21X1
XAOI21X1_532 BUFX4_67/Y MUX2X1_50/S NOR2X1_644/Y gnd AOI21X1_532/Y vdd AOI21X1
XAOI21X1_543 BUFX4_443/Y NOR2X1_107/B NOR2X1_655/Y gnd AOI21X1_543/Y vdd AOI21X1
XAOI21X1_554 BUFX4_439/Y AOI21X1_72/B NOR2X1_666/Y gnd AOI21X1_554/Y vdd AOI21X1
XAOI21X1_565 BUFX4_321/Y MUX2X1_92/S NOR2X1_677/Y gnd AOI21X1_565/Y vdd AOI21X1
XAOI21X1_576 BUFX4_73/Y MUX2X1_340/S NOR2X1_688/Y gnd AOI21X1_576/Y vdd AOI21X1
XAOI21X1_587 BUFX4_420/Y INVX1_219/A NOR2X1_699/Y gnd AOI21X1_587/Y vdd AOI21X1
XAOI21X1_598 BUFX4_324/Y NOR2X1_707/B NOR2X1_710/Y gnd AOI21X1_598/Y vdd AOI21X1
XXOR2X1_4 OR2X2_7/A OR2X2_7/B gnd XOR2X1_4/Y vdd XOR2X1
XMUX2X1_5 INVX1_8/Y MUX2X1_1/B MUX2X1_6/S gnd MUX2X1_5/Y vdd MUX2X1
XFILL_42_2_1 gnd vdd FILL
XCLKBUF1_6 BUFX4_2/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_100 BUFX4_87/A gnd BUFX4_100/Y vdd BUFX4
XBUFX4_111 BUFX4_82/A gnd BUFX4_111/Y vdd BUFX4
XBUFX4_133 INVX8_8/Y gnd BUFX4_133/Y vdd BUFX4
XBUFX4_122 BUFX4_124/A gnd INVX4_5/A vdd BUFX4
XBUFX4_155 INVX8_32/Y gnd BUFX4_155/Y vdd BUFX4
XBUFX4_144 INVX8_7/Y gnd BUFX4_144/Y vdd BUFX4
XNOR2X1_215 NOR2X1_467/A MUX2X1_376/S gnd NOR2X1_215/Y vdd NOR2X1
XBUFX4_188 INVX8_9/Y gnd BUFX4_188/Y vdd BUFX4
XBUFX4_166 INVX8_29/Y gnd BUFX4_166/Y vdd BUFX4
XBUFX4_177 INVX8_13/Y gnd BUFX4_177/Y vdd BUFX4
XNOR2X1_204 NOR2X1_204/A NOR2X1_707/B gnd NOR2X1_204/Y vdd NOR2X1
XNOR2X1_237 NOR2X1_237/A NOR2X1_234/Y gnd NOR2X1_237/Y vdd NOR2X1
XBUFX4_199 INVX8_27/Y gnd BUFX4_199/Y vdd BUFX4
XNOR2X1_226 NOR2X1_226/A NOR2X1_716/B gnd NOR2X1_226/Y vdd NOR2X1
XNOR2X1_248 NOR2X1_248/A NOR2X1_729/B gnd NOR2X1_248/Y vdd NOR2X1
XNOR2X1_259 NOR2X1_601/A MUX2X1_400/S gnd NOR2X1_259/Y vdd NOR2X1
XFILL_33_2_1 gnd vdd FILL
XFILL_17_2 gnd vdd FILL
XOAI21X1_1001 INVX1_393/Y BUFX4_248/Y BUFX4_97/Y gnd AOI21X1_433/C vdd OAI21X1
XOAI21X1_1012 MUX2X1_245/Y BUFX4_366/Y BUFX4_101/Y gnd AOI21X1_434/C vdd OAI21X1
XDFFPOSX1_602 NAND2X1_8/A CLKBUF1_28/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XOAI21X1_1023 NOR2X1_500/Y AOI21X1_439/Y BUFX4_412/Y gnd OAI21X1_1024/C vdd OAI21X1
XDFFPOSX1_613 INVX1_20/A CLKBUF1_78/Y MUX2X1_15/Y gnd vdd DFFPOSX1
XOAI21X1_1045 OAI21X1_1044/Y AND2X2_46/Y OAI21X1_1045/C gnd OAI21X1_1048/B vdd OAI21X1
XOAI21X1_1034 NOR2X1_502/Y AOI21X1_444/Y BUFX4_415/Y gnd OAI21X1_1035/C vdd OAI21X1
XOAI21X1_1056 INVX1_150/Y BUFX4_231/Y NAND2X1_322/Y gnd MUX2X1_250/B vdd OAI21X1
XOAI21X1_1078 OAI21X1_1077/Y AND2X2_49/Y OAI21X1_1076/Y gnd OAI21X1_1078/Y vdd OAI21X1
XOAI21X1_1089 NOR2X1_521/Y OAI21X1_1089/B OAI21X1_1087/Y gnd MUX2X1_256/A vdd OAI21X1
XDFFPOSX1_635 NOR2X1_23/A CLKBUF1_21/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_624 OAI21X1_12/C CLKBUF1_84/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_646 NOR2X1_31/A CLKBUF1_21/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XOAI21X1_1067 OAI21X1_1067/A AND2X2_47/Y OAI21X1_1065/Y gnd NAND2X1_328/B vdd OAI21X1
XDFFPOSX1_657 NOR2X1_494/A CLKBUF1_88/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_668 NOR2X1_41/A CLKBUF1_4/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_679 INVX1_38/A CLKBUF1_87/Y MUX2X1_30/Y gnd vdd DFFPOSX1
XINVX1_380 INVX1_380/A gnd INVX1_380/Y vdd INVX1
XINVX1_391 INVX1_391/A gnd INVX1_391/Y vdd INVX1
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 INVX8_8/A gnd INVX8_8/Y vdd INVX8
XAOI21X1_351 INVX1_15/Y BUFX4_347/Y AOI21X1_351/C gnd NOR3X1_14/C vdd AOI21X1
XAOI21X1_340 BUFX4_222/Y INVX1_319/Y BUFX4_78/Y gnd AOI21X1_340/Y vdd AOI21X1
XAOI21X1_373 NOR2X1_171/A BUFX4_151/Y BUFX4_337/Y gnd AOI21X1_373/Y vdd AOI21X1
XAOI21X1_395 AND2X2_27/A NOR2X1_644/A BUFX4_89/Y gnd AOI21X1_395/Y vdd AOI21X1
XAOI21X1_384 INVX1_152/Y BUFX4_350/Y OAI21X1_877/Y gnd OAI21X1_879/A vdd AOI21X1
XAOI21X1_362 AOI21X1_362/A BUFX4_96/Y OAI21X1_830/Y gnd OAI22X1_25/C vdd AOI21X1
XDFFPOSX1_61 INVX1_166/A CLKBUF1_91/Y MUX2X1_153/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 NAND2X1_96/A CLKBUF1_73/Y OAI21X1_378/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 NAND2X1_90/A CLKBUF1_81/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_176/A CLKBUF1_21/Y MUX2X1_163/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 NOR2X1_282/A CLKBUF1_98/Y DFFPOSX1_94/D gnd vdd DFFPOSX1
XFILL_7_3_1 gnd vdd FILL
XBUFX4_17 address[0] gnd BUFX4_17/Y vdd BUFX4
XBUFX4_28 BUFX4_28/A gnd BUFX4_28/Y vdd BUFX4
XBUFX4_39 BUFX4_33/A gnd BUFX4_39/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XOAI21X1_507 OAI22X1_2/C INVX4_7/A INVX2_24/A gnd OAI21X1_507/Y vdd OAI21X1
XOAI21X1_518 OAI21X1_515/Y AND2X2_12/Y INVX4_9/Y gnd OAI21X1_520/A vdd OAI21X1
XOAI21X1_529 AOI21X1_237/Y OAI21X1_510/Y AOI22X1_6/A gnd AOI22X1_8/B vdd OAI21X1
XDFFPOSX1_421 INVX2_16/A CLKBUF1_59/Y XNOR2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_410 NOR2X1_690/A CLKBUF1_71/Y AOI21X1_578/Y gnd vdd DFFPOSX1
XDFFPOSX1_454 NOR2X1_706/A CLKBUF1_95/Y AOI21X1_594/Y gnd vdd DFFPOSX1
XDFFPOSX1_465 NOR2X1_709/A CLKBUF1_4/Y AOI21X1_597/Y gnd vdd DFFPOSX1
XDFFPOSX1_432 NOR2X1_2/A CLKBUF1_11/Y XOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_443 INVX1_258/A CLKBUF1_39/Y OAI21X1_1454/Y gnd vdd DFFPOSX1
XDFFPOSX1_498 NOR2X1_567/B CLKBUF1_79/Y DFFPOSX1_498/D gnd vdd DFFPOSX1
XDFFPOSX1_487 INVX1_253/A CLKBUF1_7/Y MUX2X1_378/Y gnd vdd DFFPOSX1
XDFFPOSX1_476 NOR2X1_713/A CLKBUF1_1/Y AOI21X1_601/Y gnd vdd DFFPOSX1
XNOR2X1_590 BUFX4_394/Y NOR2X1_590/B gnd OAI22X1_81/A vdd NOR2X1
XAOI21X1_192 BUFX4_468/Y NOR2X1_33/Y NOR2X1_289/Y gnd AOI21X1_192/Y vdd AOI21X1
XAOI21X1_181 BUFX4_468/Y NOR2X1_16/Y NOR2X1_278/Y gnd DFFPOSX1_81/D vdd AOI21X1
XAOI21X1_170 BUFX4_214/Y NOR2X1_737/B NOR2X1_266/Y gnd DFFPOSX1_22/D vdd AOI21X1
XFILL_47_1_1 gnd vdd FILL
XFILL_30_0_1 gnd vdd FILL
XFILL_38_1_1 gnd vdd FILL
XFILL_50_8_0 gnd vdd FILL
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_304 BUFX4_132/Y BUFX4_459/Y INVX1_283/A gnd OAI21X1_304/Y vdd OAI21X1
XOAI21X1_337 BUFX4_217/Y NAND2X1_81/Y OAI21X1_337/C gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_326 BUFX4_389/Y BUFX4_310/Y AOI21X1_510/A gnd OAI21X1_327/C vdd OAI21X1
XOAI21X1_315 NAND2X1_78/Y BUFX4_176/Y OAI21X1_314/Y gnd OAI21X1_315/Y vdd OAI21X1
XOAI21X1_348 INVX4_3/A BUFX4_195/Y INVX1_403/A gnd OAI21X1_349/C vdd OAI21X1
XOAI21X1_359 NAND2X1_84/Y MUX2X1_83/B OAI21X1_359/C gnd OAI21X1_359/Y vdd OAI21X1
XDFFPOSX1_240 OAI21X1_935/B CLKBUF1_19/Y DFFPOSX1_240/D gnd vdd DFFPOSX1
XBUFX4_2 clock gnd BUFX4_2/Y vdd BUFX4
XDFFPOSX1_262 INVX1_237/A CLKBUF1_29/Y OAI21X1_1431/Y gnd vdd DFFPOSX1
XDFFPOSX1_273 INVX1_423/A CLKBUF1_26/Y DFFPOSX1_273/D gnd vdd DFFPOSX1
XDFFPOSX1_251 NOR2X1_697/A CLKBUF1_39/Y AOI21X1_585/Y gnd vdd DFFPOSX1
XDFFPOSX1_284 OAI21X1_957/B CLKBUF1_82/Y DFFPOSX1_284/D gnd vdd DFFPOSX1
XDFFPOSX1_295 INVX1_456/A CLKBUF1_56/Y MUX2X1_326/Y gnd vdd DFFPOSX1
XNAND2X1_310 BUFX4_393/Y AOI22X1_29/Y gnd AOI22X1_31/A vdd NAND2X1
XNAND2X1_321 NAND2X1_96/A AND2X2_37/B gnd NAND2X1_321/Y vdd NAND2X1
XNAND2X1_332 BUFX4_205/Y NAND2X1_332/B gnd OAI22X1_50/C vdd NAND2X1
XNAND2X1_343 OAI21X1_115/C BUFX4_271/Y gnd NAND2X1_343/Y vdd NAND2X1
XNAND2X1_354 traffic_Street_0[2] NOR2X1_97/B gnd NAND2X1_354/Y vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_29_1_1 gnd vdd FILL
XFILL_41_8_0 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XOAI21X1_860 INVX1_103/Y BUFX4_276/Y OAI21X1_860/C gnd OAI21X1_860/Y vdd OAI21X1
XOAI21X1_893 INVX1_142/Y BUFX4_234/Y OAI21X1_893/C gnd MUX2X1_227/A vdd OAI21X1
XOAI21X1_882 BUFX4_360/Y INVX1_156/A BUFX4_149/Y gnd OAI22X1_30/C vdd OAI21X1
XOAI21X1_871 INVX1_185/Y BUFX4_285/Y OAI21X1_871/C gnd MUX2X1_224/A vdd OAI21X1
XMUX2X1_360 INVX1_427/Y MUX2X1_29/B MUX2X1_360/S gnd MUX2X1_360/Y vdd MUX2X1
XMUX2X1_382 BUFX4_428/Y INVX1_320/Y NOR2X1_232/Y gnd MUX2X1_382/Y vdd MUX2X1
XMUX2X1_393 AND2X2_6/B INVX1_441/Y NOR2X1_729/B gnd MUX2X1_393/Y vdd MUX2X1
XMUX2X1_371 BUFX4_324/Y INVX1_433/Y MUX2X1_369/S gnd MUX2X1_371/Y vdd MUX2X1
XFILL_49_9_0 gnd vdd FILL
XFILL_32_8_0 gnd vdd FILL
XNAND3X1_5 NAND3X1_5/A NAND3X1_5/B NAND3X1_5/C gnd AOI22X1_1/D vdd NAND3X1
XFILL_23_8_0 gnd vdd FILL
XOAI21X1_101 BUFX4_189/Y BUFX4_478/Y OAI21X1_101/C gnd OAI21X1_101/Y vdd OAI21X1
XOAI21X1_112 MUX2X1_64/B NAND2X1_39/Y OAI21X1_112/C gnd OAI21X1_112/Y vdd OAI21X1
XOAI21X1_156 BUFX4_386/Y BUFX4_187/Y INVX1_395/A gnd OAI21X1_156/Y vdd OAI21X1
XOAI21X1_145 MUX2X1_39/B NAND2X1_51/Y OAI21X1_144/Y gnd OAI21X1_145/Y vdd OAI21X1
XOAI21X1_134 BUFX4_121/Y BUFX4_397/Y OAI21X1_134/C gnd OAI21X1_134/Y vdd OAI21X1
XOAI21X1_123 BUFX4_449/Y BUFX4_54/Y NOR2X1_579/A gnd OAI21X1_123/Y vdd OAI21X1
XOAI21X1_167 NAND2X1_53/Y BUFX4_467/Y OAI21X1_167/C gnd OAI21X1_167/Y vdd OAI21X1
XOAI21X1_189 MUX2X1_82/B NAND2X1_58/Y OAI21X1_188/Y gnd OAI21X1_189/Y vdd OAI21X1
XOAI21X1_178 INVX4_3/A BUFX4_128/Y NAND2X1_259/A gnd OAI21X1_179/C vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XNAND2X1_162 INVX2_16/A police_Interrupt gnd NOR2X1_349/A vdd NAND2X1
XNAND2X1_151 NAND3X1_44/Y NAND3X1_51/Y gnd NAND2X1_151/Y vdd NAND2X1
XNAND2X1_140 NAND3X1_10/Y NAND3X1_11/C gnd OR2X2_6/B vdd NAND2X1
XFILL_6_9_0 gnd vdd FILL
XNAND2X1_184 BUFX4_275/Y NAND2X1_184/B gnd OAI21X1_608/C vdd NAND2X1
XNAND2X1_195 OAI21X1_59/C BUFX4_227/Y gnd OAI21X1_630/C vdd NAND2X1
XNAND2X1_173 BUFX4_231/Y NOR2X1_646/A gnd OAI21X1_564/C vdd NAND2X1
XFILL_14_8_0 gnd vdd FILL
XAOI22X1_29 AOI22X1_29/A AOI22X1_29/B AOI22X1_29/C BUFX4_167/Y gnd AOI22X1_29/Y vdd
+ AOI22X1
XAOI22X1_18 INVX4_13/Y MUX2X1_191/Y AOI22X1_18/C AOI22X1_18/D gnd AOI22X1_18/Y vdd
+ AOI22X1
XOAI21X1_1408 BUFX4_452/Y BUFX4_405/Y INVX1_309/A gnd OAI21X1_1408/Y vdd OAI21X1
XOAI21X1_1419 NAND2X1_62/Y BUFX4_73/Y OAI21X1_1419/C gnd OAI21X1_1419/Y vdd OAI21X1
XOAI21X1_690 INVX1_286/Y BUFX4_288/Y NAND2X1_217/Y gnd MUX2X1_201/A vdd OAI21X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XMUX2X1_190 MUX2X1_190/A MUX2X1_190/B BUFX4_390/Y gnd MUX2X1_190/Y vdd MUX2X1
XFILL_5_2 gnd vdd FILL
XAOI21X1_40 BUFX4_216/Y MUX2X1_45/S NOR2X1_78/Y gnd AOI21X1_40/Y vdd AOI21X1
XAOI21X1_62 MUX2X1_71/B AOI21X1_62/B NOR2X1_111/Y gnd AOI21X1_62/Y vdd AOI21X1
XAOI21X1_51 MUX2X1_58/A NOR2X1_92/B NOR2X1_95/Y gnd AOI21X1_51/Y vdd AOI21X1
XAOI21X1_84 MUX2X1_49/A MUX2X1_92/S NOR2X1_143/Y gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_73 BUFX4_180/Y AOI21X1_72/B NOR2X1_127/Y gnd AOI21X1_73/Y vdd AOI21X1
XAOI21X1_95 BUFX4_216/Y MUX2X1_340/S AOI21X1_95/C gnd AOI21X1_95/Y vdd AOI21X1
XOAI21X1_2 MUX2X1_1/B NAND2X1_6/B OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XBUFX4_304 BUFX4_306/A gnd OAI22X1_2/C vdd BUFX4
XBUFX4_337 BUFX4_30/Y gnd BUFX4_337/Y vdd BUFX4
XBUFX4_326 BUFX4_28/Y gnd BUFX4_326/Y vdd BUFX4
XBUFX4_315 INVX8_1/Y gnd MUX2X1_29/B vdd BUFX4
XBUFX4_348 BUFX4_25/Y gnd BUFX4_348/Y vdd BUFX4
XFILL_46_7_0 gnd vdd FILL
XBUFX4_359 BUFX4_30/Y gnd BUFX4_359/Y vdd BUFX4
XNOR2X1_408 NOR2X1_408/A BUFX4_240/Y gnd NOR2X1_408/Y vdd NOR2X1
XNOR2X1_419 BUFX4_41/Y NOR2X1_419/B gnd NOR2X1_419/Y vdd NOR2X1
XOAI22X1_70 OAI22X1_70/A OAI22X1_70/B OAI22X1_70/C NOR2X1_579/Y gnd OAI22X1_70/Y vdd
+ OAI22X1
XOAI22X1_81 OAI22X1_81/A OAI22X1_81/B NOR2X1_576/Y OAI22X1_81/D gnd OAI22X1_81/Y vdd
+ OAI22X1
XOAI22X1_92 OAI22X1_92/A OAI22X1_92/B OAI22X1_92/C NOR2X1_621/Y gnd OAI22X1_92/Y vdd
+ OAI22X1
XOAI21X1_1238 NOR2X1_293/A BUFX4_368/Y AOI21X1_508/Y gnd OAI21X1_1239/C vdd OAI21X1
XOAI21X1_1216 BUFX4_361/Y NOR2X1_134/A BUFX4_154/Y gnd OAI22X1_78/C vdd OAI21X1
XOAI21X1_1227 INVX1_174/Y BUFX4_229/Y BUFX4_100/Y gnd AOI21X1_504/C vdd OAI21X1
XDFFPOSX1_806 OAI21X1_140/C CLKBUF1_63/Y OAI21X1_141/Y gnd vdd DFFPOSX1
XOAI21X1_1205 OAI21X1_198/C BUFX4_283/Y BUFX4_91/Y gnd OAI22X1_73/B vdd OAI21X1
XOAI21X1_1249 BUFX4_359/Y OAI21X1_246/C BUFX4_147/Y gnd OAI22X1_89/C vdd OAI21X1
XDFFPOSX1_828 AOI21X1_378/A CLKBUF1_2/Y OAI21X1_163/Y gnd vdd DFFPOSX1
XDFFPOSX1_839 INVX1_97/A CLKBUF1_85/Y MUX2X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_817 NAND2X1_303/A CLKBUF1_17/Y OAI21X1_149/Y gnd vdd DFFPOSX1
XFILL_37_7_0 gnd vdd FILL
XAOI21X1_500 NOR2X1_176/A BUFX4_289/Y AOI21X1_500/C gnd AOI21X1_500/Y vdd AOI21X1
XAOI21X1_522 BUFX4_64/Y NOR2X1_65/Y NOR2X1_634/Y gnd AOI21X1_522/Y vdd AOI21X1
XFILL_20_6_0 gnd vdd FILL
XAOI21X1_511 NAND2X1_352/Y AOI21X1_510/Y AOI21X1_511/C gnd AOI21X1_511/Y vdd AOI21X1
XAOI21X1_544 MUX2X1_6/B NOR2X1_107/B NOR2X1_656/Y gnd AOI21X1_544/Y vdd AOI21X1
XAOI21X1_533 BUFX4_324/Y MUX2X1_55/S NOR2X1_645/Y gnd AOI21X1_533/Y vdd AOI21X1
XAOI21X1_577 BUFX4_320/Y MUX2X1_340/S NOR2X1_689/Y gnd AOI21X1_577/Y vdd AOI21X1
XAOI21X1_555 BUFX4_424/Y AOI21X1_72/B NOR2X1_667/Y gnd AOI21X1_555/Y vdd AOI21X1
XAOI21X1_566 BUFX4_441/Y MUX2X1_94/S NOR2X1_678/Y gnd AOI21X1_566/Y vdd AOI21X1
XAOI21X1_599 BUFX4_420/Y MUX2X1_369/S NOR2X1_711/Y gnd AOI21X1_599/Y vdd AOI21X1
XAOI21X1_588 BUFX4_66/Y INVX1_219/A NOR2X1_700/Y gnd AOI21X1_588/Y vdd AOI21X1
XFILL_3_7_0 gnd vdd FILL
XXOR2X1_5 NOR2X1_4/Y NOR2X1_2/A gnd XOR2X1_5/Y vdd XOR2X1
XFILL_28_7_0 gnd vdd FILL
XMUX2X1_6 INVX1_9/Y MUX2X1_6/B MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XFILL_11_6_0 gnd vdd FILL
XCLKBUF1_7 BUFX4_4/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XBUFX4_101 BUFX4_87/A gnd BUFX4_101/Y vdd BUFX4
XBUFX4_112 BUFX4_85/A gnd BUFX4_112/Y vdd BUFX4
XFILL_19_7_0 gnd vdd FILL
XBUFX4_134 INVX8_8/Y gnd NOR2X1_96/B vdd BUFX4
XBUFX4_123 BUFX4_124/A gnd BUFX4_123/Y vdd BUFX4
XBUFX4_145 INVX8_7/Y gnd NOR2X1_39/B vdd BUFX4
XBUFX4_156 INVX8_32/Y gnd BUFX4_156/Y vdd BUFX4
XBUFX4_178 INVX8_13/Y gnd BUFX4_178/Y vdd BUFX4
XBUFX4_167 INVX8_29/Y gnd BUFX4_167/Y vdd BUFX4
XNOR2X1_205 BUFX4_161/Y BUFX4_61/Y gnd MUX2X1_369/S vdd NOR2X1
XNOR2X1_216 NOR2X1_216/A MUX2X1_376/S gnd NOR2X1_216/Y vdd NOR2X1
XNOR2X1_238 NOR2X1_238/A NOR2X1_234/Y gnd NOR2X1_238/Y vdd NOR2X1
XBUFX4_189 INVX8_9/Y gnd BUFX4_189/Y vdd BUFX4
XNOR2X1_249 NOR2X1_249/A NOR2X1_729/B gnd NOR2X1_249/Y vdd NOR2X1
XNOR2X1_227 BUFX4_457/Y BUFX4_142/Y gnd NOR2X1_231/B vdd NOR2X1
XFILL_17_3 gnd vdd FILL
XOAI21X1_1002 INVX1_394/Y BUFX4_251/Y BUFX4_150/Y gnd OAI21X1_1002/Y vdd OAI21X1
XOAI21X1_1013 MUX2X1_247/Y BUFX4_357/Y BUFX4_155/Y gnd OAI21X1_1014/A vdd OAI21X1
XDFFPOSX1_603 INVX1_8/A CLKBUF1_91/Y MUX2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_614 INVX1_21/A CLKBUF1_28/Y MUX2X1_16/Y gnd vdd DFFPOSX1
XOAI21X1_1024 AOI21X1_438/Y BUFX4_413/Y OAI21X1_1024/C gnd AOI22X1_29/C vdd OAI21X1
XOAI21X1_1035 AOI21X1_443/Y BUFX4_416/Y OAI21X1_1035/C gnd AOI22X1_30/C vdd OAI21X1
XOAI21X1_1046 INVX1_402/Y INVX8_31/A BUFX4_158/Y gnd AOI21X1_449/C vdd OAI21X1
XDFFPOSX1_647 INVX1_274/A CLKBUF1_84/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_636 NOR2X1_24/A CLKBUF1_30/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_625 OAI21X1_14/C CLKBUF1_40/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XOAI21X1_1057 INVX1_403/Y BUFX4_233/Y NAND2X1_323/Y gnd MUX2X1_250/A vdd OAI21X1
XOAI21X1_1079 INVX1_407/Y BUFX4_258/Y BUFX4_155/Y gnd AOI21X1_459/C vdd OAI21X1
XOAI21X1_1068 INVX1_132/Y AND2X2_52/A BUFX4_147/Y gnd AOI21X1_456/C vdd OAI21X1
XDFFPOSX1_669 NOR2X1_42/A CLKBUF1_4/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XDFFPOSX1_658 OAI21X1_41/C CLKBUF1_63/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XINVX1_381 INVX1_381/A gnd INVX1_381/Y vdd INVX1
XINVX1_392 INVX1_392/A gnd INVX1_392/Y vdd INVX1
XINVX8_9 INVX8_9/A gnd INVX8_9/Y vdd INVX8
XAOI21X1_352 INVX1_330/Y AND2X2_22/A AOI21X1_352/C gnd NOR3X1_14/B vdd AOI21X1
XAOI21X1_341 AOI21X1_341/A AOI21X1_341/B BUFX4_417/Y gnd AOI21X1_342/C vdd AOI21X1
XAOI21X1_330 BUFX4_272/Y INVX1_308/Y AOI21X1_330/C gnd AOI21X1_331/C vdd AOI21X1
XAOI21X1_374 NOR2X1_179/A BUFX4_151/Y BUFX4_337/Y gnd OAI21X1_852/C vdd AOI21X1
XAOI21X1_385 INVX1_339/Y BUFX4_290/Y OAI21X1_878/Y gnd AOI21X1_385/Y vdd AOI21X1
XAOI21X1_363 INVX1_74/Y BUFX4_262/Y OAI21X1_836/Y gnd AOI21X1_364/C vdd AOI21X1
XAOI21X1_396 BUFX4_411/Y OAI21X1_920/Y BUFX4_49/Y gnd AOI21X1_396/Y vdd AOI21X1
XDFFPOSX1_62 INVX1_167/A CLKBUF1_98/Y MUX2X1_154/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 NAND2X1_325/A CLKBUF1_72/Y OAI21X1_365/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 NAND2X1_91/A CLKBUF1_73/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XDFFPOSX1_84 INVX1_177/A CLKBUF1_66/Y MUX2X1_164/Y gnd vdd DFFPOSX1
XDFFPOSX1_73 NAND2X1_97/A CLKBUF1_72/Y DFFPOSX1_73/D gnd vdd DFFPOSX1
XDFFPOSX1_95 NOR2X1_283/A CLKBUF1_47/Y AOI21X1_186/Y gnd vdd DFFPOSX1
XBUFX4_29 BUFX4_28/A gnd BUFX4_29/Y vdd BUFX4
XBUFX4_18 address[0] gnd BUFX4_18/Y vdd BUFX4
XFILL_43_5_0 gnd vdd FILL
XFILL_34_5_0 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XOAI21X1_508 OAI22X1_2/C INVX2_20/Y INVX2_25/Y gnd AOI21X1_234/B vdd OAI21X1
XOAI21X1_519 INVX2_19/A INVX2_18/A INVX2_21/Y gnd AND2X2_13/A vdd OAI21X1
XDFFPOSX1_422 INVX2_17/A CLKBUF1_59/Y AND2X2_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_400 INVX4_7/A CLKBUF1_3/Y NAND2X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_411 INVX1_310/A CLKBUF1_33/Y MUX2X1_341/Y gnd vdd DFFPOSX1
XDFFPOSX1_433 INVX2_4/A CLKBUF1_11/Y XNOR2X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_455 OAI21X1_603/B CLKBUF1_10/Y OAI21X1_1458/Y gnd vdd DFFPOSX1
XDFFPOSX1_444 NOR2X1_702/A CLKBUF1_10/Y AOI21X1_590/Y gnd vdd DFFPOSX1
XDFFPOSX1_477 INVX1_377/A CLKBUF1_95/Y MUX2X1_376/Y gnd vdd DFFPOSX1
XDFFPOSX1_499 NOR2X1_715/A CLKBUF1_18/Y AOI21X1_603/Y gnd vdd DFFPOSX1
XDFFPOSX1_488 NOR2X1_714/A CLKBUF1_44/Y AOI21X1_602/Y gnd vdd DFFPOSX1
XDFFPOSX1_466 NOR2X1_710/A CLKBUF1_22/Y AOI21X1_598/Y gnd vdd DFFPOSX1
XFILL_0_5_0 gnd vdd FILL
XFILL_25_5_0 gnd vdd FILL
XNOR2X1_580 INVX1_76/A BUFX4_355/Y gnd OAI22X1_70/A vdd NOR2X1
XNOR2X1_591 NOR2X1_591/A BUFX4_290/Y gnd OAI22X1_76/D vdd NOR2X1
XAOI21X1_160 BUFX4_217/Y NOR2X1_733/B NOR2X1_251/Y gnd AOI21X1_160/Y vdd AOI21X1
XAOI21X1_182 BUFX4_213/Y AOI21X1_7/B NOR2X1_279/Y gnd AOI21X1_182/Y vdd AOI21X1
XAOI21X1_171 MUX2X1_40/B NOR2X1_737/B NOR2X1_267/Y gnd AOI21X1_171/Y vdd AOI21X1
XAOI21X1_193 MUX2X1_71/B NOR2X1_43/B NOR2X1_290/Y gnd AOI21X1_193/Y vdd AOI21X1
XFILL_8_6_0 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XFILL_50_8_1 gnd vdd FILL
XOAI21X1_305 MUX2X1_39/B NAND2X1_77/Y OAI21X1_304/Y gnd OAI21X1_305/Y vdd OAI21X1
XOAI21X1_338 BUFX4_194/Y BUFX4_308/Y DFFPOSX1_7/Q gnd OAI21X1_339/C vdd OAI21X1
XOAI21X1_316 BUFX4_310/Y BUFX4_300/Y INVX1_407/A gnd OAI21X1_317/C vdd OAI21X1
XOAI21X1_327 NAND2X1_79/Y BUFX4_469/Y OAI21X1_327/C gnd OAI21X1_327/Y vdd OAI21X1
XOAI21X1_349 NAND2X1_82/Y MUX2X1_86/B OAI21X1_349/C gnd OAI21X1_349/Y vdd OAI21X1
XDFFPOSX1_230 INVX1_225/A CLKBUF1_92/Y DFFPOSX1_230/D gnd vdd DFFPOSX1
XBUFX4_3 clock gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_241 OAI21X1_1087/B CLKBUF1_94/Y DFFPOSX1_241/D gnd vdd DFFPOSX1
XDFFPOSX1_252 INVX1_358/A CLKBUF1_13/Y MUX2X1_355/Y gnd vdd DFFPOSX1
XDFFPOSX1_263 INVX1_306/A CLKBUF1_39/Y OAI21X1_1433/Y gnd vdd DFFPOSX1
XDFFPOSX1_274 INVX1_257/A CLKBUF1_37/Y MUX2X1_357/Y gnd vdd DFFPOSX1
XDFFPOSX1_285 OAI21X1_1153/B CLKBUF1_82/Y OAI21X1_1445/Y gnd vdd DFFPOSX1
XDFFPOSX1_296 INVX1_457/A CLKBUF1_34/Y MUX2X1_327/Y gnd vdd DFFPOSX1
XNAND2X1_300 BUFX4_48/Y OAI21X1_993/Y gnd NAND2X1_300/Y vdd NAND2X1
XNAND2X1_311 NAND2X1_311/A BUFX4_272/Y gnd NAND2X1_311/Y vdd NAND2X1
XNAND2X1_322 NOR2X1_263/A BUFX4_230/Y gnd NAND2X1_322/Y vdd NAND2X1
XNAND2X1_333 BUFX4_207/Y NAND2X1_333/B gnd OAI22X1_52/C vdd NAND2X1
XNAND2X1_344 NOR2X1_95/A BUFX4_273/Y gnd NAND2X1_344/Y vdd NAND2X1
XNAND2X1_355 traffic_Street_0[3] NOR2X1_107/B gnd NAND2X1_355/Y vdd NAND2X1
XFILL_41_8_1 gnd vdd FILL
XFILL_40_3_0 gnd vdd FILL
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XOAI21X1_850 AND2X2_32/Y OAI21X1_850/B OAI21X1_850/C gnd NAND2X1_256/B vdd OAI21X1
XOAI21X1_872 NOR2X1_291/A BUFX4_355/Y OAI21X1_872/C gnd OAI21X1_873/C vdd OAI21X1
XOAI21X1_861 NOR2X1_143/A BUFX4_277/Y BUFX4_110/Y gnd AOI21X1_379/C vdd OAI21X1
XOAI21X1_883 NAND2X1_91/A BUFX4_223/Y BUFX4_76/Y gnd OAI22X1_30/B vdd OAI21X1
XOAI21X1_894 BUFX4_331/Y NOR2X1_224/A BUFX4_155/Y gnd OAI22X1_31/C vdd OAI21X1
XMUX2X1_350 INVX1_238/Y BUFX4_437/Y MUX2X1_353/S gnd MUX2X1_350/Y vdd MUX2X1
XMUX2X1_361 BUFX4_444/Y INVX1_259/Y MUX2X1_364/S gnd MUX2X1_361/Y vdd MUX2X1
XMUX2X1_383 BUFX4_63/Y INVX1_383/Y NOR2X1_232/Y gnd MUX2X1_383/Y vdd MUX2X1
XMUX2X1_372 BUFX4_444/Y INVX1_256/Y MUX2X1_120/S gnd MUX2X1_372/Y vdd MUX2X1
XMUX2X1_394 BUFX4_439/Y INVX1_263/Y MUX2X1_397/S gnd MUX2X1_394/Y vdd MUX2X1
XFILL_49_9_1 gnd vdd FILL
XFILL_48_4_0 gnd vdd FILL
XFILL_32_8_1 gnd vdd FILL
XFILL_31_3_0 gnd vdd FILL
XNAND3X1_6 AND2X2_2/B NAND3X1_5/A NAND3X1_6/C gnd NAND3X1_8/B vdd NAND3X1
XFILL_39_4_0 gnd vdd FILL
XFILL_23_8_1 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 BUFX4_218/Y NAND2X1_37/Y OAI21X1_101/Y gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_113 BUFX4_56/Y BUFX4_53/Y OAI21X1_113/C gnd OAI21X1_114/C vdd OAI21X1
XOAI21X1_146 BUFX4_59/Y BUFX4_183/Y INVX1_336/A gnd OAI21X1_147/C vdd OAI21X1
XOAI21X1_135 NAND2X1_48/Y MUX2X1_71/B OAI21X1_134/Y gnd OAI21X1_135/Y vdd OAI21X1
XOAI21X1_124 NAND2X1_40/Y MUX2X1_58/A OAI21X1_123/Y gnd OAI21X1_124/Y vdd OAI21X1
XOAI21X1_168 BUFX4_129/Y BUFX4_301/Y NOR2X1_396/A gnd OAI21X1_169/C vdd OAI21X1
XOAI21X1_179 NAND2X1_57/Y MUX2X1_49/A OAI21X1_179/C gnd OAI21X1_179/Y vdd OAI21X1
XOAI21X1_157 NAND2X1_52/Y BUFX4_381/Y OAI21X1_156/Y gnd OAI21X1_157/Y vdd OAI21X1
XNAND2X1_141 NAND2X1_141/A OAI21X1_497/Y gnd NOR2X1_334/A vdd NAND2X1
XNAND2X1_152 NAND3X1_55/Y NAND3X1_53/Y gnd NAND2X1_152/Y vdd NAND2X1
XNAND2X1_130 NAND3X1_19/B NAND3X1_19/C gnd INVX1_196/A vdd NAND2X1
XNAND2X1_163 NAND3X1_68/B AND2X2_18/A gnd OAI21X1_538/C vdd NAND2X1
XFILL_6_9_1 gnd vdd FILL
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_185 BUFX4_277/Y NOR2X1_715/A gnd OAI21X1_609/C vdd NAND2X1
XNAND2X1_196 BUFX4_31/Y OAI22X1_6/Y gnd OAI21X1_633/C vdd NAND2X1
XNAND2X1_174 BUFX4_38/Y MUX2X1_177/Y gnd AOI22X1_12/D vdd NAND2X1
XFILL_14_8_1 gnd vdd FILL
XFILL_13_3_0 gnd vdd FILL
XAOI22X1_19 AOI22X1_19/A AOI22X1_19/B AOI22X1_19/C BUFX4_171/Y gnd AOI22X1_19/Y vdd
+ AOI22X1
XOAI21X1_1409 NAND2X1_61/Y BUFX4_422/Y OAI21X1_1408/Y gnd OAI21X1_1409/Y vdd OAI21X1
XNOR3X1_9 NOR3X1_3/Y INVX4_11/Y NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XOAI21X1_691 MUX2X1_95/B BUFX4_290/Y NAND2X1_218/Y gnd MUX2X1_202/B vdd OAI21X1
XOAI21X1_680 BUFX4_153/Y INVX1_97/A BUFX4_278/Y gnd OAI21X1_681/B vdd OAI21X1
XMUX2X1_180 AOI22X1_13/Y MUX2X1_180/B BUFX4_394/Y gnd MUX2X1_180/Y vdd MUX2X1
XMUX2X1_191 AOI22X1_14/Y AOI22X1_17/Y INVX4_14/Y gnd MUX2X1_191/Y vdd MUX2X1
XAOI21X1_52 MUX2X1_59/B NOR2X1_97/B NOR2X1_97/Y gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_30 MUX2X1_82/B NOR2X1_60/Y NOR2X1_63/Y gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_41 BUFX4_216/Y NOR2X1_83/B NOR2X1_80/Y gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_85 BUFX4_467/Y MUX2X1_92/S AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XAOI21X1_74 BUFX4_381/Y AOI21X1_72/B AOI21X1_74/C gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_63 MUX2X1_40/B AOI21X1_62/B AOI21X1_63/C gnd AOI21X1_63/Y vdd AOI21X1
XOAI21X1_3 MUX2X1_6/B NAND2X1_6/B OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XAOI21X1_96 BUFX4_174/Y MUX2X1_340/S NOR2X1_160/Y gnd AOI21X1_96/Y vdd AOI21X1
XBUFX4_305 BUFX4_306/A gnd BUFX4_305/Y vdd BUFX4
XBUFX4_327 BUFX4_27/Y gnd BUFX4_327/Y vdd BUFX4
XBUFX4_316 INVX8_1/Y gnd BUFX4_316/Y vdd BUFX4
XFILL_46_7_1 gnd vdd FILL
XBUFX4_349 BUFX4_28/Y gnd BUFX4_349/Y vdd BUFX4
XBUFX4_338 BUFX4_25/Y gnd BUFX4_338/Y vdd BUFX4
XFILL_45_2_0 gnd vdd FILL
XNOR2X1_409 INVX1_77/A AND2X2_47/B gnd OAI22X1_19/D vdd NOR2X1
XOAI22X1_60 NOR2X1_524/Y OAI22X1_60/B OAI22X1_60/C OAI22X1_60/D gnd OAI22X1_60/Y vdd
+ OAI22X1
XOAI22X1_82 NOR2X1_602/Y OAI22X1_82/B OAI22X1_82/C NOR2X1_601/Y gnd OAI22X1_82/Y vdd
+ OAI22X1
XOAI22X1_93 BUFX4_400/Y OAI22X1_93/B AND2X2_54/Y OAI22X1_93/D gnd OAI22X1_93/Y vdd
+ OAI22X1
XOAI22X1_71 OAI22X1_71/A OAI22X1_71/B OAI22X1_71/C NOR2X1_581/Y gnd OAI22X1_71/Y vdd
+ OAI22X1
XOAI21X1_1206 BUFX4_342/Y NOR2X1_162/A BUFX4_148/Y gnd OAI22X1_74/C vdd OAI21X1
XOAI21X1_1228 INVX1_170/Y BUFX4_346/Y BUFX4_149/Y gnd OAI21X1_1229/A vdd OAI21X1
XOAI21X1_1217 OAI21X1_182/C BUFX4_222/Y BUFX4_96/Y gnd OAI22X1_78/B vdd OAI21X1
XDFFPOSX1_829 INVX1_396/A CLKBUF1_2/Y OAI21X1_165/Y gnd vdd DFFPOSX1
XDFFPOSX1_818 OAI21X1_150/C CLKBUF1_75/Y OAI21X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_807 INVX1_290/A CLKBUF1_77/Y AOI21X1_62/Y gnd vdd DFFPOSX1
XOAI21X1_1239 NOR2X1_608/Y OAI21X1_1239/B OAI21X1_1239/C gnd NOR2X1_609/B vdd OAI21X1
XFILL_37_7_1 gnd vdd FILL
XFILL_36_2_0 gnd vdd FILL
XAOI21X1_501 INVX1_154/Y BUFX4_363/Y AOI21X1_501/C gnd AOI21X1_501/Y vdd AOI21X1
XAOI21X1_523 MUX2X1_8/B NOR2X1_65/Y NOR2X1_635/Y gnd AOI21X1_523/Y vdd AOI21X1
XFILL_20_6_1 gnd vdd FILL
XAOI21X1_512 INVX1_409/Y NOR2X1_624/A NOR2X1_624/Y gnd AOI21X1_512/Y vdd AOI21X1
XAOI21X1_534 BUFX4_443/Y NOR2X1_92/B NOR2X1_646/Y gnd AOI21X1_534/Y vdd AOI21X1
XAOI21X1_556 BUFX4_67/Y AOI21X1_72/B NOR2X1_668/Y gnd AOI21X1_556/Y vdd AOI21X1
XAOI21X1_567 BUFX4_426/Y MUX2X1_94/S NOR2X1_679/Y gnd AOI21X1_567/Y vdd AOI21X1
XAOI21X1_545 BUFX4_69/Y NOR2X1_107/B NOR2X1_657/Y gnd AOI21X1_545/Y vdd AOI21X1
XAOI21X1_578 AND2X2_5/B NOR2X1_167/B NOR2X1_690/Y gnd AOI21X1_578/Y vdd AOI21X1
XAOI21X1_589 BUFX4_317/Y INVX1_219/A NOR2X1_701/Y gnd AOI21X1_589/Y vdd AOI21X1
XFILL_3_7_1 gnd vdd FILL
XFILL_28_7_1 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XMUX2X1_7 INVX1_10/Y BUFX4_71/Y MUX2X1_6/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_11_6_1 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XCLKBUF1_8 BUFX4_8/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XBUFX4_102 BUFX4_82/A gnd BUFX4_102/Y vdd BUFX4
XBUFX4_124 BUFX4_124/A gnd BUFX4_124/Y vdd BUFX4
XBUFX4_146 INVX8_32/Y gnd BUFX4_146/Y vdd BUFX4
XFILL_19_7_1 gnd vdd FILL
XBUFX4_113 BUFX4_85/A gnd BUFX4_113/Y vdd BUFX4
XBUFX4_135 INVX8_8/Y gnd BUFX4_135/Y vdd BUFX4
XBUFX4_157 INVX8_32/Y gnd BUFX4_157/Y vdd BUFX4
XBUFX4_179 INVX8_13/Y gnd MUX2X1_49/A vdd BUFX4
XFILL_18_2_0 gnd vdd FILL
XBUFX4_168 INVX8_29/Y gnd BUFX4_168/Y vdd BUFX4
XNOR2X1_206 NOR2X1_206/A MUX2X1_369/S gnd NOR2X1_206/Y vdd NOR2X1
XNOR2X1_217 NOR2X1_613/A MUX2X1_376/S gnd NOR2X1_217/Y vdd NOR2X1
XNOR2X1_239 INVX2_12/Y INVX2_8/Y gnd INVX8_26/A vdd NOR2X1
XNOR2X1_228 NOR2X1_384/A NOR2X1_231/B gnd NOR2X1_228/Y vdd NOR2X1
XOAI21X1_1003 OAI21X1_1002/Y AND2X2_44/Y BUFX4_39/Y gnd OAI22X1_44/A vdd OAI21X1
XOAI21X1_1025 INVX1_58/Y BUFX4_106/Y BUFX4_330/Y gnd OAI21X1_1025/Y vdd OAI21X1
XDFFPOSX1_604 INVX1_9/A CLKBUF1_98/Y MUX2X1_6/Y gnd vdd DFFPOSX1
XOAI21X1_1014 OAI21X1_1014/A NOR2X1_498/Y BUFX4_50/Y gnd OAI21X1_1015/B vdd OAI21X1
XOAI21X1_1036 INVX1_88/Y BUFX4_282/Y NAND2X1_315/Y gnd MUX2X1_249/B vdd OAI21X1
XDFFPOSX1_637 NOR2X1_25/A CLKBUF1_103/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XOAI21X1_1058 INVX1_153/Y BUFX4_235/Y NAND2X1_324/Y gnd MUX2X1_251/B vdd OAI21X1
XDFFPOSX1_626 OAI21X1_16/C CLKBUF1_91/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_648 INVX1_331/A CLKBUF1_84/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_615 INVX1_22/A CLKBUF1_76/Y MUX2X1_17/Y gnd vdd DFFPOSX1
XOAI21X1_1069 INVX1_134/Y BUFX4_247/Y BUFX4_79/Y gnd AOI21X1_457/C vdd OAI21X1
XOAI21X1_1047 INVX1_182/Y BUFX4_223/Y BUFX4_115/Y gnd AOI21X1_450/C vdd OAI21X1
XINVX1_360 INVX1_360/A gnd INVX1_360/Y vdd INVX1
XINVX1_371 INVX1_371/A gnd INVX1_371/Y vdd INVX1
XDFFPOSX1_659 OAI21X1_43/C CLKBUF1_63/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XINVX1_393 INVX1_393/A gnd INVX1_393/Y vdd INVX1
XINVX1_382 INVX1_382/A gnd INVX1_382/Y vdd INVX1
XAOI21X1_342 BUFX4_418/Y MUX2X1_214/Y AOI21X1_342/C gnd MUX2X1_216/A vdd AOI21X1
XAOI21X1_320 BUFX4_252/Y NOR2X1_656/A BUFX4_104/Y gnd OAI21X1_731/C vdd AOI21X1
XAOI21X1_331 BUFX4_147/Y AOI21X1_331/B AOI21X1_331/C gnd AOI21X1_332/B vdd AOI21X1
XAOI21X1_386 NAND2X1_263/Y OAI21X1_879/Y BUFX4_207/Y gnd AOI21X1_386/Y vdd AOI21X1
XAOI21X1_353 BUFX4_240/Y INVX1_5/Y BUFX4_87/Y gnd OAI21X1_801/C vdd AOI21X1
XAOI21X1_364 BUFX4_152/Y OAI21X1_835/Y AOI21X1_364/C gnd AOI21X1_364/Y vdd AOI21X1
XAOI21X1_375 BUFX4_418/Y AOI21X1_375/B BUFX4_168/Y gnd AOI22X1_22/D vdd AOI21X1
XAOI21X1_397 AOI21X1_396/Y AOI21X1_397/B BUFX4_402/Y gnd AOI22X1_24/B vdd AOI21X1
XDFFPOSX1_41 INVX1_443/A CLKBUF1_25/Y DFFPOSX1_41/D gnd vdd DFFPOSX1
XDFFPOSX1_52 NAND2X1_92/A CLKBUF1_47/Y DFFPOSX1_52/D gnd vdd DFFPOSX1
XDFFPOSX1_63 INVX1_168/A CLKBUF1_73/Y MUX2X1_155/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 NOR2X1_271/A CLKBUF1_11/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_178/A CLKBUF1_103/Y MUX2X1_165/Y gnd vdd DFFPOSX1
XDFFPOSX1_96 NOR2X1_284/A CLKBUF1_21/Y AOI21X1_187/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX1_280/A CLKBUF1_66/Y OAI21X1_381/Y gnd vdd DFFPOSX1
XOAI21X1_1570 MUX2X1_6/B NAND2X1_2/Y NAND2X1_362/Y gnd DFFPOSX1_592/D vdd OAI21X1
XBUFX4_19 address[0] gnd BUFX4_19/Y vdd BUFX4
XFILL_43_5_1 gnd vdd FILL
XFILL_42_0_0 gnd vdd FILL
XFILL_34_5_1 gnd vdd FILL
XFILL_22_2 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XOAI21X1_509 NOR2X1_334/B NOR3X1_12/A AOI21X1_236/Y gnd AOI21X1_237/B vdd OAI21X1
XFILL_15_1 gnd vdd FILL
XDFFPOSX1_401 INVX4_6/A CLKBUF1_3/Y NAND2X1_152/Y gnd vdd DFFPOSX1
XDFFPOSX1_412 NOR2X1_691/A CLKBUF1_44/Y AOI21X1_579/Y gnd vdd DFFPOSX1
XDFFPOSX1_456 NAND2X1_238/A CLKBUF1_49/Y OAI21X1_1460/Y gnd vdd DFFPOSX1
XDFFPOSX1_423 MUX2X1_176/B CLKBUF1_59/Y MUX2X1_176/Y gnd vdd DFFPOSX1
XDFFPOSX1_434 NOR2X1_1/B CLKBUF1_14/Y OAI21X1_548/Y gnd vdd DFFPOSX1
XDFFPOSX1_445 INVX1_380/A CLKBUF1_39/Y DFFPOSX1_445/D gnd vdd DFFPOSX1
XDFFPOSX1_467 INVX1_254/A CLKBUF1_82/Y MUX2X1_369/Y gnd vdd DFFPOSX1
XDFFPOSX1_478 INVX1_434/A CLKBUF1_61/Y MUX2X1_377/Y gnd vdd DFFPOSX1
XDFFPOSX1_489 INVX1_375/A CLKBUF1_65/Y MUX2X1_379/Y gnd vdd DFFPOSX1
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XFILL_0_5_1 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XNOR2X1_570 BUFX4_39/Y NOR2X1_570/B gnd NOR2X1_570/Y vdd NOR2X1
XFILL_24_0_0 gnd vdd FILL
XNOR2X1_592 NOR2X1_124/A BUFX4_330/Y gnd NOR2X1_592/Y vdd NOR2X1
XNOR2X1_581 INVX1_89/A BUFX4_277/Y gnd NOR2X1_581/Y vdd NOR2X1
XAOI21X1_150 MUX2X1_86/B NOR2X1_234/Y NOR2X1_237/Y gnd AOI21X1_150/Y vdd AOI21X1
XAOI21X1_194 BUFX4_177/Y NOR2X1_43/B NOR2X1_291/Y gnd AOI21X1_194/Y vdd AOI21X1
XAOI21X1_183 BUFX4_375/Y AOI21X1_7/B NOR2X1_280/Y gnd AOI21X1_183/Y vdd AOI21X1
XAOI21X1_161 BUFX4_180/Y NOR2X1_733/B NOR2X1_252/Y gnd AOI21X1_161/Y vdd AOI21X1
XAOI21X1_172 MUX2X1_86/B NOR2X1_737/B NOR2X1_268/Y gnd AOI21X1_172/Y vdd AOI21X1
XFILL_8_6_1 gnd vdd FILL
XDFFPOSX1_990 NOR2X1_615/A CLKBUF1_74/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XFILL_7_1_0 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XOAI21X1_306 BUFX4_137/Y BUFX4_455/Y OAI21X1_306/C gnd OAI21X1_307/C vdd OAI21X1
XOAI21X1_328 NOR2X1_84/B BUFX4_308/Y INVX1_282/A gnd OAI21X1_329/C vdd OAI21X1
XOAI21X1_317 NAND2X1_78/Y BUFX4_380/Y OAI21X1_317/C gnd OAI21X1_317/Y vdd OAI21X1
XOAI21X1_339 BUFX4_180/Y NAND2X1_81/Y OAI21X1_339/C gnd DFFPOSX1_7/D vdd OAI21X1
XDFFPOSX1_220 INVX1_360/A CLKBUF1_40/Y MUX2X1_274/Y gnd vdd DFFPOSX1
XDFFPOSX1_231 INVX1_300/A CLKBUF1_92/Y DFFPOSX1_231/D gnd vdd DFFPOSX1
XBUFX4_4 clock gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_242 INVX1_238/A CLKBUF1_61/Y MUX2X1_350/Y gnd vdd DFFPOSX1
XDFFPOSX1_264 AND2X2_40/B CLKBUF1_13/Y DFFPOSX1_264/D gnd vdd DFFPOSX1
XDFFPOSX1_253 INVX1_421/A CLKBUF1_86/Y MUX2X1_356/Y gnd vdd DFFPOSX1
XDFFPOSX1_275 INVX1_317/A CLKBUF1_50/Y MUX2X1_358/Y gnd vdd DFFPOSX1
XDFFPOSX1_286 INVX1_245/A CLKBUF1_32/Y DFFPOSX1_286/D gnd vdd DFFPOSX1
XDFFPOSX1_297 INVX1_458/A CLKBUF1_32/Y MUX2X1_328/Y gnd vdd DFFPOSX1
XNAND2X1_301 NAND2X1_301/A BUFX4_252/Y gnd NAND2X1_301/Y vdd NAND2X1
XNAND2X1_323 NOR2X1_268/A BUFX4_232/Y gnd NAND2X1_323/Y vdd NAND2X1
XNAND2X1_312 NOR2X1_104/A BUFX4_274/Y gnd NAND2X1_312/Y vdd NAND2X1
XNAND2X1_345 BUFX4_33/Y MUX2X1_261/Y gnd NAND2X1_345/Y vdd NAND2X1
XNAND2X1_334 AND2X2_41/A NOR2X1_696/A gnd AOI21X1_473/A vdd NAND2X1
XNAND2X1_356 traffic_Street_0[0] NAND2X1_50/B gnd NAND2X1_356/Y vdd NAND2X1
XFILL_40_3_1 gnd vdd FILL
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XOAI21X1_851 INVX1_117/Y BUFX4_108/Y BUFX4_344/Y gnd OAI21X1_853/B vdd OAI21X1
XOAI21X1_840 INVX1_82/A BUFX4_265/Y BUFX4_102/Y gnd AOI21X1_369/C vdd OAI21X1
XOAI21X1_862 MUX2X1_88/B BUFX4_112/Y NAND2X1_258/Y gnd MUX2X1_220/B vdd OAI21X1
XOAI21X1_884 OAI22X1_30/Y BUFX4_417/Y INVX8_29/A gnd AOI21X1_387/C vdd OAI21X1
XOAI21X1_873 BUFX4_117/Y OAI21X1_873/B OAI21X1_873/C gnd OAI21X1_874/A vdd OAI21X1
XOAI21X1_895 OAI21X1_895/A BUFX4_236/Y BUFX4_80/Y gnd OAI22X1_31/B vdd OAI21X1
XMUX2X1_340 BUFX4_437/Y INVX1_240/Y MUX2X1_340/S gnd MUX2X1_340/Y vdd MUX2X1
XMUX2X1_362 MUX2X1_27/B INVX1_315/Y MUX2X1_364/S gnd MUX2X1_362/Y vdd MUX2X1
XMUX2X1_373 BUFX4_70/Y INVX1_378/Y MUX2X1_120/S gnd MUX2X1_373/Y vdd MUX2X1
XMUX2X1_384 BUFX4_322/Y INVX1_436/Y NOR2X1_232/Y gnd MUX2X1_384/Y vdd MUX2X1
XMUX2X1_351 INVX1_305/Y BUFX4_420/Y MUX2X1_353/S gnd MUX2X1_351/Y vdd MUX2X1
XMUX2X1_395 BUFX4_428/Y INVX1_323/Y MUX2X1_397/S gnd MUX2X1_395/Y vdd MUX2X1
XFILL_48_4_1 gnd vdd FILL
XFILL_31_3_1 gnd vdd FILL
XNAND3X1_7 INVX4_6/Y INVX1_187/Y NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XFILL_39_4_1 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_103 BUFX4_193/Y NOR2X1_74/B AOI21X1_362/A gnd OAI21X1_104/C vdd OAI21X1
XOAI21X1_147 BUFX4_176/Y NAND2X1_51/Y OAI21X1_147/C gnd OAI21X1_147/Y vdd OAI21X1
XOAI21X1_136 BUFX4_121/Y BUFX4_396/Y INVX1_334/A gnd OAI21X1_136/Y vdd OAI21X1
XOAI21X1_114 MUX2X1_44/A NAND2X1_39/Y OAI21X1_114/C gnd OAI21X1_114/Y vdd OAI21X1
XOAI21X1_125 BUFX4_58/Y BUFX4_397/Y OAI21X1_125/C gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_169 NAND2X1_56/Y BUFX4_214/Y OAI21X1_169/C gnd OAI21X1_169/Y vdd OAI21X1
XOAI21X1_158 NOR2X1_77/B BUFX4_183/Y OAI21X1_158/C gnd OAI21X1_159/C vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd north_South[0] vdd BUFX2
XNAND2X1_153 INVX1_206/A NAND2X1_146/Y gnd NOR3X1_12/C vdd NAND2X1
XNAND2X1_142 AND2X2_10/B AND2X2_10/A gnd NAND3X1_46/B vdd NAND2X1
XNAND2X1_120 OAI21X1_467/Y NOR2X1_349/B gnd INVX4_9/A vdd NAND2X1
XNAND2X1_131 INVX1_196/A INVX1_201/A gnd NAND2X1_132/B vdd NAND2X1
XNAND2X1_164 MUX2X1_176/B NOR3X1_7/Y gnd MUX2X1_176/A vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_175 BUFX4_233/Y NAND2X1_175/B gnd NAND2X1_175/Y vdd NAND2X1
XNAND2X1_186 AND2X2_41/A NOR2X1_719/A gnd OAI21X1_610/C vdd NAND2X1
XNAND2X1_197 NOR2X1_271/A BUFX4_232/Y gnd OAI21X1_640/C vdd NAND2X1
XFILL_13_3_1 gnd vdd FILL
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 MUX2X1_1/B NOR2X1_16/Y NOR2X1_17/Y gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_681 NOR2X1_394/Y OAI21X1_681/B OAI21X1_679/Y gnd OAI21X1_681/Y vdd OAI21X1
XOAI21X1_670 INVX1_284/Y BUFX4_268/Y OAI21X1_670/C gnd OAI21X1_672/C vdd OAI21X1
XOAI21X1_692 INVX1_287/Y AND2X2_46/B NAND2X1_219/Y gnd MUX2X1_202/A vdd OAI21X1
XMUX2X1_192 MUX2X1_192/A MUX2X1_192/B BUFX4_112/Y gnd MUX2X1_192/Y vdd MUX2X1
XMUX2X1_170 BUFX4_209/Y INVX1_184/Y MUX2X1_31/S gnd MUX2X1_170/Y vdd MUX2X1
XMUX2X1_181 MUX2X1_181/A MUX2X1_181/B BUFX4_38/Y gnd MUX2X1_181/Y vdd MUX2X1
XAOI21X1_31 BUFX4_473/Y NOR2X1_60/Y NOR2X1_64/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_20 MUX2X1_6/B NOR2X1_47/B NOR2X1_46/Y gnd AOI21X1_20/Y vdd AOI21X1
XAOI21X1_42 MUX2X1_40/B NOR2X1_83/B NOR2X1_81/Y gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_53 MUX2X1_64/B NOR2X1_97/B NOR2X1_98/Y gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_75 BUFX4_467/Y AOI21X1_72/B AOI21X1_75/C gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_86 BUFX4_217/Y MUX2X1_94/S AOI21X1_86/C gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_64 BUFX4_371/Y AOI21X1_62/B NOR2X1_113/Y gnd AOI21X1_64/Y vdd AOI21X1
XOAI21X1_4 BUFX4_71/Y NAND2X1_6/B NAND2X1_7/Y gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_97 BUFX4_380/Y MUX2X1_340/S AOI21X1_97/C gnd AOI21X1_97/Y vdd AOI21X1
XBUFX4_306 BUFX4_306/A gnd BUFX4_306/Y vdd BUFX4
XBUFX4_328 BUFX4_30/Y gnd BUFX4_328/Y vdd BUFX4
XBUFX4_317 INVX8_1/Y gnd BUFX4_317/Y vdd BUFX4
XBUFX4_339 BUFX4_26/Y gnd BUFX4_339/Y vdd BUFX4
XFILL_45_2_1 gnd vdd FILL
XOAI22X1_61 OAI22X1_61/A OAI22X1_61/B OAI22X1_61/C OAI22X1_61/D gnd NOR2X1_554/B vdd
+ OAI22X1
XOAI22X1_50 MUX2X1_256/Y BUFX4_206/Y OAI22X1_50/C OAI22X1_50/D gnd OAI22X1_50/Y vdd
+ OAI22X1
XOAI22X1_83 NOR2X1_605/Y OAI22X1_83/B OAI22X1_83/C NOR2X1_604/Y gnd OAI22X1_83/Y vdd
+ OAI22X1
XOAI22X1_94 OAI22X1_94/A OAI22X1_94/B OAI22X1_94/C NOR2X1_548/Y gnd OAI22X1_94/Y vdd
+ OAI22X1
XOAI22X1_72 OAI22X1_72/A NOR2X1_578/Y OAI22X1_72/C BUFX4_207/Y gnd OAI22X1_72/Y vdd
+ OAI22X1
XOAI21X1_1229 OAI21X1_1229/A NOR2X1_603/Y BUFX4_410/Y gnd OAI21X1_1229/Y vdd OAI21X1
XOAI21X1_1218 BUFX4_329/Y OAI21X1_190/C BUFX4_150/Y gnd OAI22X1_79/C vdd OAI21X1
XOAI21X1_1207 OAI21X1_222/C BUFX4_285/Y BUFX4_92/Y gnd OAI22X1_74/B vdd OAI21X1
XDFFPOSX1_819 OAI21X1_678/A CLKBUF1_17/Y OAI21X1_153/Y gnd vdd DFFPOSX1
XDFFPOSX1_808 NOR2X1_112/A CLKBUF1_20/Y AOI21X1_63/Y gnd vdd DFFPOSX1
XFILL_3_1 gnd vdd FILL
XFILL_45_1 gnd vdd FILL
XFILL_36_2_1 gnd vdd FILL
XAOI21X1_524 MUX2X1_4/B NOR2X1_70/Y NOR2X1_636/Y gnd AOI21X1_524/Y vdd AOI21X1
XAOI21X1_513 BUFX4_442/Y NOR2X1_54/Y NOR2X1_625/Y gnd AOI21X1_513/Y vdd AOI21X1
XAOI21X1_502 INVX1_443/Y AND2X2_37/B AOI21X1_502/C gnd AOI21X1_502/Y vdd AOI21X1
XAOI21X1_557 BUFX4_322/Y AOI21X1_72/B NOR2X1_669/Y gnd AOI21X1_557/Y vdd AOI21X1
XAOI21X1_568 BUFX4_65/Y MUX2X1_94/S NOR2X1_680/Y gnd AOI21X1_568/Y vdd AOI21X1
XAOI21X1_546 MUX2X1_9/B AOI21X1_62/B NOR2X1_658/Y gnd AOI21X1_546/Y vdd AOI21X1
XAOI21X1_535 BUFX4_430/Y NOR2X1_92/B NOR2X1_647/Y gnd AOI21X1_535/Y vdd AOI21X1
XAOI21X1_579 BUFX4_73/Y NOR2X1_167/B NOR2X1_691/Y gnd AOI21X1_579/Y vdd AOI21X1
XFILL_2_2_1 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B MUX2X1_6/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 BUFX4_9/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XBUFX4_103 BUFX4_82/A gnd BUFX4_103/Y vdd BUFX4
XBUFX4_125 BUFX4_124/A gnd BUFX4_125/Y vdd BUFX4
XBUFX4_136 INVX8_8/Y gnd BUFX4_136/Y vdd BUFX4
XBUFX4_114 BUFX4_85/A gnd BUFX4_114/Y vdd BUFX4
XNOR2X1_207 NOR2X1_207/A MUX2X1_369/S gnd NOR2X1_207/Y vdd NOR2X1
XFILL_18_2_1 gnd vdd FILL
XBUFX4_169 INVX8_29/Y gnd BUFX4_169/Y vdd BUFX4
XBUFX4_158 INVX8_32/Y gnd BUFX4_158/Y vdd BUFX4
XBUFX4_147 INVX8_32/Y gnd BUFX4_147/Y vdd BUFX4
XNOR2X1_229 NOR2X1_460/A NOR2X1_231/B gnd NOR2X1_229/Y vdd NOR2X1
XNOR2X1_218 BUFX4_163/Y BUFX4_119/Y gnd NOR2X1_220/B vdd NOR2X1
XFILL_30_9_0 gnd vdd FILL
XOAI21X1_1004 MUX2X1_91/B BUFX4_253/Y NAND2X1_301/Y gnd MUX2X1_241/B vdd OAI21X1
XOAI21X1_1026 INVX1_399/Y BUFX4_150/Y AOI21X1_440/Y gnd OAI21X1_1026/Y vdd OAI21X1
XDFFPOSX1_605 INVX1_10/A CLKBUF1_78/Y MUX2X1_7/Y gnd vdd DFFPOSX1
XOAI21X1_1015 AOI21X1_434/Y OAI21X1_1015/B OAI21X1_1010/Y gnd NAND2X1_308/B vdd OAI21X1
XOAI21X1_1037 INVX1_400/Y BUFX4_284/Y NAND2X1_316/Y gnd MUX2X1_249/A vdd OAI21X1
XDFFPOSX1_638 INVX1_32/A CLKBUF1_91/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_627 NOR2X1_17/A CLKBUF1_103/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XOAI21X1_1059 INVX1_404/Y BUFX4_237/Y NAND2X1_325/Y gnd MUX2X1_251/A vdd OAI21X1
XDFFPOSX1_616 INVX1_24/A CLKBUF1_47/Y MUX2X1_18/Y gnd vdd DFFPOSX1
XOAI21X1_1048 BUFX4_37/Y OAI21X1_1048/B NAND2X1_320/Y gnd OAI21X1_1049/A vdd OAI21X1
XINVX1_361 INVX1_361/A gnd INVX1_361/Y vdd INVX1
XDFFPOSX1_649 OAI21X1_31/C CLKBUF1_103/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XINVX1_350 INVX1_350/A gnd INVX1_350/Y vdd INVX1
XINVX1_372 INVX1_372/A gnd INVX1_372/Y vdd INVX1
XINVX1_394 INVX1_394/A gnd INVX1_394/Y vdd INVX1
XINVX1_383 INVX1_383/A gnd INVX1_383/Y vdd INVX1
XNOR2X1_730 NOR2X1_730/A NOR2X1_733/B gnd NOR2X1_730/Y vdd NOR2X1
XFILL_21_9_0 gnd vdd FILL
XAOI21X1_343 BUFX4_230/Y NOR2X1_731/A BUFX4_83/Y gnd AOI21X1_343/Y vdd AOI21X1
XAOI21X1_321 INVX8_30/A OAI21X1_733/Y BUFX4_171/Y gnd AOI22X1_19/B vdd AOI21X1
XAOI21X1_332 BUFX4_35/Y AOI21X1_332/B BUFX4_166/Y gnd AOI22X1_20/A vdd AOI21X1
XAOI21X1_310 BUFX4_168/Y MUX2X1_203/Y AOI21X1_310/C gnd OAI21X1_698/B vdd AOI21X1
XAOI21X1_354 INVX1_35/Y BUFX4_368/Y BUFX4_156/Y gnd OAI21X1_807/C vdd AOI21X1
XAOI21X1_376 NOR2X1_122/A BUFX4_34/Y OAI21X1_854/Y gnd AOI21X1_376/Y vdd AOI21X1
XAOI21X1_365 BUFX4_415/Y AOI21X1_364/Y BUFX4_204/Y gnd AOI22X1_21/B vdd AOI21X1
XAOI21X1_398 BUFX4_259/Y NOR2X1_673/A AOI21X1_398/C gnd OAI22X1_37/B vdd AOI21X1
XDFFPOSX1_20 INVX1_403/A CLKBUF1_14/Y OAI21X1_349/Y gnd vdd DFFPOSX1
XAOI21X1_387 BUFX4_418/Y MUX2X1_225/Y AOI21X1_387/C gnd OAI21X1_885/A vdd AOI21X1
XDFFPOSX1_53 NAND2X1_93/A CLKBUF1_21/Y DFFPOSX1_53/D gnd vdd DFFPOSX1
XDFFPOSX1_31 NOR2X1_272/A CLKBUF1_25/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_42 AND2X2_24/B CLKBUF1_81/Y DFFPOSX1_42/D gnd vdd DFFPOSX1
XDFFPOSX1_86 NOR2X1_279/A CLKBUF1_84/Y AOI21X1_182/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 NOR2X1_449/A CLKBUF1_91/Y OAI21X1_383/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 INVX1_169/A CLKBUF1_30/Y MUX2X1_156/Y gnd vdd DFFPOSX1
XOAI21X1_1560 NAND2X1_84/Y BUFX4_324/Y OAI21X1_1560/C gnd OAI21X1_1560/Y vdd OAI21X1
XOAI21X1_1571 BUFX4_69/Y NAND2X1_2/Y NAND2X1_363/Y gnd DFFPOSX1_593/D vdd OAI21X1
XDFFPOSX1_97 NOR2X1_285/A CLKBUF1_21/Y DFFPOSX1_97/D gnd vdd DFFPOSX1
XFILL_42_0_1 gnd vdd FILL
XFILL_12_9_0 gnd vdd FILL
XFILL_33_0_1 gnd vdd FILL
XDFFPOSX1_413 NOR2X1_692/A CLKBUF1_45/Y AOI21X1_580/Y gnd vdd DFFPOSX1
XDFFPOSX1_402 INVX2_14/A CLKBUF1_3/Y OAI21X1_520/Y gnd vdd DFFPOSX1
XDFFPOSX1_435 INVX4_1/A CLKBUF1_42/Y XNOR2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_424 NAND2X1_160/A CLKBUF1_3/Y XNOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_446 INVX1_428/A CLKBUF1_10/Y OAI21X1_1456/Y gnd vdd DFFPOSX1
XDFFPOSX1_468 NOR2X1_711/A CLKBUF1_50/Y AOI21X1_599/Y gnd vdd DFFPOSX1
XDFFPOSX1_479 INVX1_252/A CLKBUF1_89/Y OAI21X1_1466/Y gnd vdd DFFPOSX1
XDFFPOSX1_457 OAI21X1_961/B CLKBUF1_10/Y DFFPOSX1_457/D gnd vdd DFFPOSX1
XINVX1_191 XNOR2X1_1/B gnd INVX1_191/Y vdd INVX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XNOR2X1_571 OAI21X1_73/C BUFX4_262/Y gnd NOR2X1_571/Y vdd NOR2X1
XNOR2X1_560 NOR2X1_560/A BUFX4_232/Y gnd OAI22X1_64/D vdd NOR2X1
XFILL_24_0_1 gnd vdd FILL
XNOR2X1_593 NOR2X1_593/A AND2X2_46/B gnd NOR2X1_593/Y vdd NOR2X1
XNOR2X1_582 NOR2X1_582/A BUFX4_339/Y gnd OAI22X1_71/A vdd NOR2X1
XAOI21X1_151 BUFX4_467/Y NOR2X1_234/Y NOR2X1_238/Y gnd AOI21X1_151/Y vdd AOI21X1
XAOI21X1_140 BUFX4_218/Y NOR2X1_716/B NOR2X1_223/Y gnd AOI21X1_140/Y vdd AOI21X1
XAOI21X1_184 BUFX4_468/Y AOI21X1_7/B NOR2X1_281/Y gnd AOI21X1_184/Y vdd AOI21X1
XAOI21X1_162 MUX2X1_86/B NOR2X1_733/B NOR2X1_253/Y gnd AOI21X1_162/Y vdd AOI21X1
XAOI21X1_173 BUFX4_473/Y NOR2X1_737/B NOR2X1_269/Y gnd DFFPOSX1_25/D vdd AOI21X1
XAOI21X1_195 BUFX4_371/Y NOR2X1_43/B NOR2X1_292/Y gnd AOI21X1_195/Y vdd AOI21X1
XOAI21X1_1390 BUFX4_387/Y BUFX4_403/Y OAI21X1_581/B gnd OAI21X1_1390/Y vdd OAI21X1
XDFFPOSX1_980 NOR2X1_211/A CLKBUF1_1/Y AOI21X1_132/Y gnd vdd DFFPOSX1
XDFFPOSX1_991 AOI21X1_304/A CLKBUF1_89/Y OAI21X1_273/Y gnd vdd DFFPOSX1
XFILL_7_1_1 gnd vdd FILL
XFILL_44_8_0 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_35_8_0 gnd vdd FILL
XOAI21X1_307 BUFX4_180/Y NAND2X1_77/Y OAI21X1_307/C gnd OAI21X1_307/Y vdd OAI21X1
XOAI21X1_329 NAND2X1_80/Y BUFX4_217/Y OAI21X1_329/C gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_318 BUFX4_310/Y BUFX4_300/Y INVX1_445/A gnd OAI21X1_319/C vdd OAI21X1
XDFFPOSX1_221 NOR2X1_523/A CLKBUF1_94/Y AOI21X1_524/Y gnd vdd DFFPOSX1
XBUFX4_5 clock gnd BUFX4_5/Y vdd BUFX4
XDFFPOSX1_210 INVX1_234/A CLKBUF1_29/Y DFFPOSX1_210/D gnd vdd DFFPOSX1
XDFFPOSX1_254 NOR2X1_671/A CLKBUF1_69/Y AOI21X1_559/Y gnd vdd DFFPOSX1
XDFFPOSX1_232 INVX1_350/A CLKBUF1_85/Y OAI21X1_1295/Y gnd vdd DFFPOSX1
XDFFPOSX1_243 INVX1_305/A CLKBUF1_39/Y MUX2X1_351/Y gnd vdd DFFPOSX1
XDFFPOSX1_276 INVX1_379/A CLKBUF1_102/Y MUX2X1_359/Y gnd vdd DFFPOSX1
XNAND2X1_302 NOR2X1_147/A AND2X2_27/A gnd NAND2X1_302/Y vdd NAND2X1
XDFFPOSX1_298 INVX1_251/A CLKBUF1_34/Y MUX2X1_321/Y gnd vdd DFFPOSX1
XDFFPOSX1_287 NOR2X1_424/B CLKBUF1_5/Y DFFPOSX1_287/D gnd vdd DFFPOSX1
XDFFPOSX1_265 OAI21X1_1436/C CLKBUF1_12/Y DFFPOSX1_265/D gnd vdd DFFPOSX1
XNAND2X1_324 NOR2X1_273/A BUFX4_234/Y gnd NAND2X1_324/Y vdd NAND2X1
XNAND2X1_313 BUFX4_31/Y MUX2X1_248/Y gnd AOI22X1_30/A vdd NAND2X1
XNAND2X1_335 NOR2X1_48/A BUFX4_234/Y gnd NAND2X1_335/Y vdd NAND2X1
XNAND2X1_357 traffic_Street_0[2] NAND2X1_50/B gnd NAND2X1_357/Y vdd NAND2X1
XNAND2X1_346 INVX8_29/A NAND2X1_346/B gnd OAI22X1_75/C vdd NAND2X1
XFILL_26_8_0 gnd vdd FILL
XFILL_1_8_0 gnd vdd FILL
XNOR2X1_390 BUFX4_201/Y NOR2X1_390/B gnd OAI22X1_12/A vdd NOR2X1
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XOAI21X1_830 INVX1_59/Y BUFX4_95/Y AND2X2_27/A gnd OAI21X1_830/Y vdd OAI21X1
XOAI21X1_841 OAI21X1_841/A AOI21X1_369/Y BUFX4_37/Y gnd OAI21X1_842/C vdd OAI21X1
XOAI21X1_852 INVX1_122/Y BUFX4_151/Y OAI21X1_852/C gnd OAI21X1_853/C vdd OAI21X1
XOAI21X1_863 INVX1_337/Y BUFX4_114/Y OAI21X1_863/C gnd MUX2X1_220/A vdd OAI21X1
XOAI21X1_885 OAI21X1_885/A AOI21X1_386/Y BUFX4_390/Y gnd OAI21X1_885/Y vdd OAI21X1
XOAI21X1_874 OAI21X1_874/A BUFX4_415/Y BUFX4_206/Y gnd OAI22X1_28/C vdd OAI21X1
XOAI21X1_896 BUFX4_32/Y MUX2X1_227/Y OAI21X1_896/C gnd NAND3X1_75/B vdd OAI21X1
XMUX2X1_330 BUFX4_65/Y INVX1_352/Y MUX2X1_88/S gnd MUX2X1_330/Y vdd MUX2X1
XMUX2X1_341 BUFX4_422/Y INVX1_310/Y NOR2X1_167/B gnd MUX2X1_341/Y vdd MUX2X1
XMUX2X1_363 BUFX4_68/Y INVX1_381/Y MUX2X1_364/S gnd MUX2X1_363/Y vdd MUX2X1
XMUX2X1_352 INVX1_359/Y BUFX4_66/Y MUX2X1_353/S gnd MUX2X1_352/Y vdd MUX2X1
XMUX2X1_374 BUFX4_324/Y INVX1_435/Y MUX2X1_120/S gnd MUX2X1_374/Y vdd MUX2X1
XFILL_9_9_0 gnd vdd FILL
XMUX2X1_385 BUFX4_439/Y INVX1_267/Y NOR2X1_233/Y gnd MUX2X1_385/Y vdd MUX2X1
XMUX2X1_396 BUFX4_67/Y INVX1_388/Y MUX2X1_397/S gnd MUX2X1_396/Y vdd MUX2X1
XFILL_17_8_0 gnd vdd FILL
XNAND3X1_8 INVX4_7/Y NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_9/B vdd NAND3X1
XFILL_50_6_0 gnd vdd FILL
XOAI21X1_104 MUX2X1_49/A NAND2X1_37/Y OAI21X1_104/C gnd OAI21X1_104/Y vdd OAI21X1
XOAI21X1_137 NAND2X1_48/Y MUX2X1_77/B OAI21X1_136/Y gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_126 MUX2X1_71/B NAND2X1_44/Y OAI21X1_125/Y gnd OAI21X1_126/Y vdd OAI21X1
XOAI21X1_115 BUFX4_61/Y BUFX4_54/Y OAI21X1_115/C gnd OAI21X1_116/C vdd OAI21X1
XOAI21X1_159 NAND2X1_52/Y BUFX4_469/Y OAI21X1_159/C gnd OAI21X1_159/Y vdd OAI21X1
XOAI21X1_148 BUFX4_59/Y BUFX4_187/Y NAND2X1_303/A gnd OAI21X1_148/Y vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd north_South[1] vdd BUFX2
XNAND2X1_110 traffic_Street_0[0] BUFX4_422/Y gnd NAND2X1_110/Y vdd NAND2X1
XNAND2X1_143 OAI22X1_2/Y NAND3X1_47/Y gnd NOR3X1_12/B vdd NAND2X1
XNAND2X1_121 NAND2X1_121/A NOR3X1_7/Y gnd NAND2X1_122/B vdd NAND2X1
XNAND2X1_132 XOR2X1_1/A NAND2X1_132/B gnd INVX2_21/A vdd NAND2X1
XNAND2X1_165 OAI21X1_539/Y INVX1_213/Y gnd NOR2X1_352/A vdd NAND2X1
XNAND2X1_154 INVX4_10/Y NAND3X1_54/C gnd AOI22X1_7/A vdd NAND2X1
XNAND2X1_187 BUFX4_281/Y NAND2X1_187/B gnd OAI21X1_611/C vdd NAND2X1
XNAND2X1_176 BUFX4_252/Y NOR2X1_678/A gnd NAND2X1_176/Y vdd NAND2X1
XNAND2X1_198 NAND2X1_198/A BUFX4_234/Y gnd NAND2X1_198/Y vdd NAND2X1
XFILL_41_6_0 gnd vdd FILL
XINVX2_2 enable gnd INVX2_2/Y vdd INVX2
XOAI21X1_660 BUFX4_331/Y NOR2X1_223/A BUFX4_155/Y gnd OAI22X1_10/C vdd OAI21X1
XAOI21X1_2 BUFX4_421/Y NOR2X1_16/Y AOI21X1_2/C gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_682 OAI21X1_681/Y BUFX4_34/Y BUFX4_165/Y gnd NOR2X1_395/B vdd OAI21X1
XOAI21X1_671 INVX1_135/Y BUFX4_270/Y BUFX4_80/Y gnd OAI21X1_671/Y vdd OAI21X1
XOAI21X1_693 INVX1_116/Y INVX8_31/A NAND2X1_220/Y gnd MUX2X1_204/B vdd OAI21X1
XMUX2X1_160 INVX1_173/Y BUFX4_375/Y MUX2X1_18/S gnd MUX2X1_160/Y vdd MUX2X1
XMUX2X1_182 MUX2X1_182/A MUX2X1_182/B BUFX4_100/Y gnd MUX2X1_182/Y vdd MUX2X1
XMUX2X1_171 MUX2X1_77/B INVX1_185/Y MUX2X1_31/S gnd MUX2X1_171/Y vdd MUX2X1
XMUX2X1_193 MUX2X1_193/A MUX2X1_193/B BUFX4_113/Y gnd MUX2X1_193/Y vdd MUX2X1
XFILL_49_7_0 gnd vdd FILL
XFILL_32_6_0 gnd vdd FILL
XFILL_23_6_0 gnd vdd FILL
XAOI21X1_10 BUFX4_64/Y NOR2X1_30/B NOR2X1_30/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_32 BUFX4_213/Y NOR2X1_65/Y NOR2X1_66/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_21 BUFX4_69/Y NOR2X1_47/B NOR2X1_47/Y gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_43 MUX2X1_44/A NOR2X1_83/B NOR2X1_82/Y gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_76 BUFX4_214/Y MUX2X1_88/S NOR2X1_132/Y gnd AOI21X1_76/Y vdd AOI21X1
XAOI21X1_54 BUFX4_371/Y NOR2X1_97/B NOR2X1_99/Y gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_65 BUFX4_470/Y AOI21X1_62/B NOR2X1_114/Y gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_98 AND2X2_3/B MUX2X1_340/S NOR2X1_162/Y gnd AOI21X1_98/Y vdd AOI21X1
XOAI21X1_5 MUX2X1_4/B NAND2X1_6/B NAND2X1_8/Y gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_87 MUX2X1_82/B MUX2X1_94/S AOI21X1_87/C gnd AOI21X1_87/Y vdd AOI21X1
XFILL_6_7_0 gnd vdd FILL
XBUFX4_307 BUFX4_306/A gnd BUFX4_307/Y vdd BUFX4
XBUFX4_318 INVX8_1/Y gnd BUFX4_318/Y vdd BUFX4
XBUFX4_329 BUFX4_29/Y gnd BUFX4_329/Y vdd BUFX4
XFILL_14_6_0 gnd vdd FILL
XOAI22X1_40 NOR2X1_493/Y OAI22X1_40/B OAI22X1_40/C OAI22X1_40/D gnd OAI22X1_40/Y vdd
+ OAI22X1
XOAI22X1_51 NOR2X1_528/Y OAI22X1_51/B OAI22X1_51/C NOR2X1_527/Y gnd OAI22X1_51/Y vdd
+ OAI22X1
XOAI22X1_84 OAI22X1_84/A OAI22X1_84/B OAI22X1_84/C OAI22X1_84/D gnd MUX2X1_263/A vdd
+ OAI22X1
XOAI22X1_62 OAI22X1_62/A OAI22X1_62/B OAI22X1_62/C OAI22X1_62/D gnd OAI22X1_62/Y vdd
+ OAI22X1
XOAI22X1_73 OAI22X1_73/A OAI22X1_73/B OAI22X1_73/C NOR2X1_585/Y gnd OAI22X1_73/Y vdd
+ OAI22X1
XOAI21X1_1219 NOR2X1_144/A BUFX4_224/Y BUFX4_97/Y gnd OAI22X1_79/B vdd OAI21X1
XOAI21X1_1208 OAI22X1_74/Y BUFX4_40/Y BUFX4_168/Y gnd OAI22X1_75/B vdd OAI21X1
XOAI21X1_490 NOR3X1_9/Y INVX2_22/Y NAND3X1_39/A gnd NOR2X1_327/B vdd OAI21X1
XDFFPOSX1_809 NOR2X1_113/A CLKBUF1_20/Y AOI21X1_64/Y gnd vdd DFFPOSX1
XFILL_3_2 gnd vdd FILL
XFILL_45_2 gnd vdd FILL
XAOI21X1_525 BUFX4_445/Y NOR2X1_76/B NOR2X1_637/Y gnd AOI21X1_525/Y vdd AOI21X1
XAOI21X1_514 BUFX4_65/Y NOR2X1_54/Y NOR2X1_626/Y gnd AOI21X1_514/Y vdd AOI21X1
XAOI21X1_503 NAND2X1_347/Y AOI21X1_503/B AND2X2_48/B gnd AOI21X1_503/Y vdd AOI21X1
XAOI21X1_558 BUFX4_426/Y MUX2X1_88/S NOR2X1_670/Y gnd AOI21X1_558/Y vdd AOI21X1
XAOI21X1_547 MUX2X1_18/B AOI21X1_62/B NOR2X1_659/Y gnd AOI21X1_547/Y vdd AOI21X1
XAOI21X1_536 BUFX4_68/Y NOR2X1_92/B NOR2X1_648/Y gnd AOI21X1_536/Y vdd AOI21X1
XAOI21X1_569 BUFX4_321/Y MUX2X1_94/S NOR2X1_681/Y gnd AOI21X1_569/Y vdd AOI21X1
XMUX2X1_9 INVX1_12/Y MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XBUFX4_137 INVX8_8/Y gnd BUFX4_137/Y vdd BUFX4
XBUFX4_104 BUFX4_75/A gnd BUFX4_104/Y vdd BUFX4
XBUFX4_115 BUFX4_85/A gnd BUFX4_115/Y vdd BUFX4
XBUFX4_126 BUFX4_124/A gnd BUFX4_126/Y vdd BUFX4
XFILL_46_5_0 gnd vdd FILL
XBUFX4_159 INVX8_32/Y gnd BUFX4_159/Y vdd BUFX4
XBUFX4_148 INVX8_32/Y gnd BUFX4_148/Y vdd BUFX4
XNOR2X1_219 NOR2X1_219/A NOR2X1_220/B gnd NOR2X1_219/Y vdd NOR2X1
XNOR2X1_208 NOR2X1_208/A MUX2X1_369/S gnd NOR2X1_208/Y vdd NOR2X1
XFILL_30_9_1 gnd vdd FILL
XOAI21X1_1005 INVX1_106/Y BUFX4_255/Y NAND2X1_302/Y gnd MUX2X1_241/A vdd OAI21X1
XOAI21X1_1027 AND2X2_45/Y OAI21X1_1025/Y OAI21X1_1026/Y gnd AOI21X1_441/B vdd OAI21X1
XOAI21X1_1016 BUFX4_167/Y MUX2X1_242/Y NAND2X1_308/Y gnd AOI22X1_31/C vdd OAI21X1
XDFFPOSX1_628 NOR2X1_18/A CLKBUF1_30/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_639 INVX1_273/A CLKBUF1_103/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XOAI21X1_1038 BUFX4_346/Y NOR2X1_277/A BUFX4_149/Y gnd NOR2X1_504/B vdd OAI21X1
XDFFPOSX1_606 INVX1_11/A CLKBUF1_28/Y MUX2X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_617 INVX1_25/A CLKBUF1_78/Y MUX2X1_19/Y gnd vdd DFFPOSX1
XOAI21X1_1049 OAI21X1_1049/A BUFX4_171/Y INVX8_28/A gnd OAI22X1_46/C vdd OAI21X1
XINVX1_351 INVX1_351/A gnd INVX1_351/Y vdd INVX1
XINVX1_340 INVX1_340/A gnd INVX1_340/Y vdd INVX1
XINVX1_362 INVX1_362/A gnd INVX1_362/Y vdd INVX1
XINVX1_384 INVX1_384/A gnd INVX1_384/Y vdd INVX1
XINVX1_373 INVX1_373/A gnd INVX1_373/Y vdd INVX1
XINVX1_395 INVX1_395/A gnd INVX1_395/Y vdd INVX1
XFILL_37_5_0 gnd vdd FILL
XNOR2X1_720 NOR2X1_720/A NOR2X1_231/B gnd NOR2X1_720/Y vdd NOR2X1
XNOR2X1_731 NOR2X1_731/A NOR2X1_733/B gnd NOR2X1_731/Y vdd NOR2X1
XAOI21X1_300 BUFX4_262/Y INVX1_283/Y BUFX4_76/Y gnd OAI21X1_662/C vdd AOI21X1
XAOI21X1_322 BUFX4_256/Y NOR2X1_643/A BUFX4_106/Y gnd AOI21X1_322/Y vdd AOI21X1
XFILL_20_4_0 gnd vdd FILL
XAOI21X1_311 BUFX4_417/Y MUX2X1_205/Y AOI21X1_311/C gnd AOI21X1_311/Y vdd AOI21X1
XFILL_21_9_1 gnd vdd FILL
XAOI21X1_333 BUFX4_276/Y INVX1_310/Y AOI21X1_333/C gnd AOI21X1_333/Y vdd AOI21X1
XAOI21X1_355 INVX1_29/Y BUFX4_326/Y BUFX4_159/Y gnd AOI21X1_355/Y vdd AOI21X1
XAOI21X1_344 BUFX4_235/Y INVX1_325/Y AOI21X1_344/C gnd AOI21X1_344/Y vdd AOI21X1
XAOI21X1_366 INVX1_87/Y BUFX4_353/Y AOI21X1_366/C gnd AOI21X1_367/C vdd AOI21X1
XAOI21X1_399 BUFX4_356/Y INVX1_354/Y AOI21X1_399/C gnd AOI21X1_399/Y vdd AOI21X1
XAOI21X1_377 NOR2X1_127/A BUFX4_419/Y BUFX4_330/Y gnd AOI21X1_377/Y vdd AOI21X1
XDFFPOSX1_10 INVX1_149/A CLKBUF1_25/Y MUX2X1_136/Y gnd vdd DFFPOSX1
XAOI21X1_388 OAI21X1_885/Y AOI21X1_388/B INVX8_33/Y gnd OAI21X1_907/A vdd AOI21X1
XDFFPOSX1_32 NOR2X1_273/A CLKBUF1_35/Y AOI21X1_176/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 NAND2X1_87/A CLKBUF1_40/Y DFFPOSX1_43/D gnd vdd DFFPOSX1
XOAI21X1_1550 NAND2X1_82/Y BUFX4_63/Y OAI21X1_1549/Y gnd OAI21X1_1550/Y vdd OAI21X1
XDFFPOSX1_54 INVX1_159/A CLKBUF1_40/Y MUX2X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 OAI21X1_350/C CLKBUF1_14/Y OAI21X1_351/Y gnd vdd DFFPOSX1
XOAI21X1_1561 BUFX4_188/Y BUFX4_195/Y OAI21X1_617/B gnd OAI21X1_1561/Y vdd OAI21X1
XDFFPOSX1_76 NOR2X1_503/A CLKBUF1_28/Y DFFPOSX1_76/D gnd vdd DFFPOSX1
XDFFPOSX1_65 INVX1_170/A CLKBUF1_21/Y MUX2X1_157/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX1_179/A CLKBUF1_21/Y OAI21X1_388/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_279/A CLKBUF1_103/Y OAI21X1_398/Y gnd vdd DFFPOSX1
XFILL_3_5_0 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XFILL_11_4_0 gnd vdd FILL
XFILL_12_9_1 gnd vdd FILL
XFILL_19_5_0 gnd vdd FILL
XDFFPOSX1_403 INVX4_8/A CLKBUF1_3/Y NAND2X1_156/Y gnd vdd DFFPOSX1
XDFFPOSX1_447 INVX1_259/A CLKBUF1_37/Y MUX2X1_361/Y gnd vdd DFFPOSX1
XDFFPOSX1_414 OAI21X1_578/B CLKBUF1_8/Y OAI21X1_1415/Y gnd vdd DFFPOSX1
XDFFPOSX1_436 INVX1_27/A CLKBUF1_42/Y OAI21X1_550/Y gnd vdd DFFPOSX1
XDFFPOSX1_425 NAND2X1_121/A CLKBUF1_3/Y OAI21X1_531/Y gnd vdd DFFPOSX1
XDFFPOSX1_458 OAI21X1_1157/B CLKBUF1_49/Y OAI21X1_1464/Y gnd vdd DFFPOSX1
XDFFPOSX1_469 INVX1_376/A CLKBUF1_102/Y MUX2X1_370/Y gnd vdd DFFPOSX1
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNOR2X1_561 NOR2X1_36/A BUFX4_332/Y gnd OAI22X1_64/A vdd NOR2X1
XNOR2X1_550 BUFX4_418/Y NOR2X1_550/B gnd OAI22X1_63/D vdd NOR2X1
XNOR2X1_583 NOR2X1_183/A BUFX4_337/Y gnd NOR2X1_583/Y vdd NOR2X1
XNOR2X1_594 INVX1_100/A BUFX4_325/Y gnd OAI22X1_77/A vdd NOR2X1
XNOR2X1_572 NOR2X1_64/A BUFX4_361/Y gnd OAI22X1_67/A vdd NOR2X1
XAOI21X1_141 BUFX4_176/Y NOR2X1_716/B NOR2X1_224/Y gnd AOI21X1_141/Y vdd AOI21X1
XAOI21X1_130 BUFX4_371/Y MUX2X1_369/S NOR2X1_208/Y gnd AOI21X1_130/Y vdd AOI21X1
XAOI21X1_163 BUFX4_467/Y NOR2X1_733/B NOR2X1_254/Y gnd DFFPOSX1_1/D vdd AOI21X1
XAOI21X1_185 BUFX4_209/Y NOR2X1_30/B NOR2X1_282/Y gnd DFFPOSX1_94/D vdd AOI21X1
XAOI21X1_174 MUX2X1_39/B MUX2X1_410/S NOR2X1_271/Y gnd DFFPOSX1_30/D vdd AOI21X1
XAOI21X1_152 BUFX4_218/Y NOR2X1_727/B NOR2X1_241/Y gnd AOI21X1_152/Y vdd AOI21X1
XAOI21X1_196 MUX2X1_66/B NOR2X1_43/B NOR2X1_293/Y gnd AOI21X1_196/Y vdd AOI21X1
XOAI21X1_1380 BUFX4_385/Y BUFX4_130/Y INVX1_423/A gnd OAI21X1_1380/Y vdd OAI21X1
XOAI21X1_1391 NAND2X1_59/Y AND2X2_5/B OAI21X1_1390/Y gnd OAI21X1_1391/Y vdd OAI21X1
XDFFPOSX1_970 INVX1_130/A CLKBUF1_61/Y MUX2X1_117/Y gnd vdd DFFPOSX1
XDFFPOSX1_992 OAI21X1_274/C CLKBUF1_7/Y OAI21X1_275/Y gnd vdd DFFPOSX1
XDFFPOSX1_981 INVX1_134/A CLKBUF1_15/Y MUX2X1_121/Y gnd vdd DFFPOSX1
XFILL_44_8_1 gnd vdd FILL
XFILL_43_3_0 gnd vdd FILL
XFILL_35_8_1 gnd vdd FILL
XFILL_34_3_0 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XOAI21X1_308 BUFX4_132/Y BUFX4_459/Y NAND2X1_329/A gnd OAI21X1_309/C vdd OAI21X1
XOAI21X1_319 NAND2X1_78/Y BUFX4_469/Y OAI21X1_319/C gnd OAI21X1_319/Y vdd OAI21X1
XBUFX4_6 clock gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_222 NOR2X1_646/A CLKBUF1_20/Y AOI21X1_534/Y gnd vdd DFFPOSX1
XDFFPOSX1_211 OAI21X1_752/B CLKBUF1_22/Y OAI21X1_1425/Y gnd vdd DFFPOSX1
XDFFPOSX1_200 NOR2X1_685/A CLKBUF1_71/Y AOI21X1_573/Y gnd vdd DFFPOSX1
XDFFPOSX1_255 NOR2X1_425/A CLKBUF1_5/Y AOI21X1_560/Y gnd vdd DFFPOSX1
XDFFPOSX1_233 AOI21X1_466/B CLKBUF1_85/Y OAI21X1_1297/Y gnd vdd DFFPOSX1
XDFFPOSX1_244 INVX1_359/A CLKBUF1_13/Y MUX2X1_352/Y gnd vdd DFFPOSX1
XDFFPOSX1_277 INVX1_427/A CLKBUF1_49/Y MUX2X1_360/Y gnd vdd DFFPOSX1
XDFFPOSX1_266 NOR2X1_698/A CLKBUF1_27/Y AOI21X1_586/Y gnd vdd DFFPOSX1
XDFFPOSX1_288 INVX1_353/A CLKBUF1_26/Y OAI21X1_1371/Y gnd vdd DFFPOSX1
XDFFPOSX1_299 INVX1_313/A CLKBUF1_34/Y MUX2X1_322/Y gnd vdd DFFPOSX1
XNAND2X1_325 NAND2X1_325/A BUFX4_236/Y gnd NAND2X1_325/Y vdd NAND2X1
XNAND2X1_303 NAND2X1_303/A BUFX4_256/Y gnd NAND2X1_303/Y vdd NAND2X1
XNAND2X1_336 OAI21X1_65/C BUFX4_236/Y gnd NAND2X1_336/Y vdd NAND2X1
XNAND2X1_314 NOR2X1_94/A BUFX4_276/Y gnd NAND2X1_314/Y vdd NAND2X1
XNAND2X1_347 BUFX4_41/Y OAI22X1_82/Y gnd NAND2X1_347/Y vdd NAND2X1
XNAND2X1_358 traffic_Street_0[0] NOR2X1_188/B gnd NAND2X1_358/Y vdd NAND2X1
XNOR3X1_10 NOR3X1_3/Y OAI22X1_2/D NOR3X1_9/C gnd NOR3X1_10/Y vdd NOR3X1
XFILL_26_8_1 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XFILL_1_8_1 gnd vdd FILL
XFILL_25_3_0 gnd vdd FILL
XNOR2X1_391 NOR2X1_118/A BUFX4_275/Y gnd OAI22X1_13/D vdd NOR2X1
XNOR2X1_380 NOR2X1_290/A BUFX4_339/Y gnd OAI22X1_7/A vdd NOR2X1
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XOAI21X1_831 INVX1_57/Y BUFX4_98/Y BUFX4_325/Y gnd OAI21X1_831/Y vdd OAI21X1
XOAI21X1_820 OAI21X1_820/A INVX4_14/Y INVX4_13/Y gnd AOI21X1_357/C vdd OAI21X1
XOAI21X1_842 AOI21X1_367/Y BUFX4_37/Y OAI21X1_842/C gnd AOI22X1_21/C vdd OAI21X1
XOAI21X1_853 AND2X2_33/Y OAI21X1_853/B OAI21X1_853/C gnd AOI21X1_375/B vdd OAI21X1
XOAI21X1_864 BUFX4_349/Y NOR2X1_276/A BUFX4_159/Y gnd OAI21X1_864/Y vdd OAI21X1
XOAI21X1_875 BUFX4_350/Y NOR2X1_262/A BUFX4_146/Y gnd OAI22X1_29/C vdd OAI21X1
XOAI21X1_897 BUFX4_359/Y OAI21X1_242/C BUFX4_147/Y gnd OAI22X1_32/C vdd OAI21X1
XOAI21X1_886 INVX1_340/Y BUFX4_225/Y NAND2X1_266/Y gnd MUX2X1_226/B vdd OAI21X1
XMUX2X1_331 BUFX4_321/Y INVX1_422/Y MUX2X1_88/S gnd MUX2X1_331/Y vdd MUX2X1
XMUX2X1_320 BUFX4_72/Y INVX1_371/Y MUX2X1_320/S gnd MUX2X1_320/Y vdd MUX2X1
XMUX2X1_364 MUX2X1_29/B INVX1_429/Y MUX2X1_364/S gnd MUX2X1_364/Y vdd MUX2X1
XMUX2X1_375 BUFX4_444/Y INVX1_255/Y MUX2X1_376/S gnd MUX2X1_375/Y vdd MUX2X1
XMUX2X1_353 INVX1_459/Y BUFX4_317/Y MUX2X1_353/S gnd MUX2X1_353/Y vdd MUX2X1
XMUX2X1_342 INVX1_236/Y BUFX4_437/Y MUX2X1_97/S gnd MUX2X1_342/Y vdd MUX2X1
XFILL_9_9_1 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XMUX2X1_386 BUFX4_424/Y INVX1_321/Y NOR2X1_233/Y gnd MUX2X1_386/Y vdd MUX2X1
XMUX2X1_397 AND2X2_6/B INVX1_439/Y MUX2X1_397/S gnd MUX2X1_397/Y vdd MUX2X1
XFILL_16_3_0 gnd vdd FILL
XFILL_17_8_1 gnd vdd FILL
XNAND3X1_9 INVX2_13/Y NAND3X1_9/B NAND3X1_9/C gnd NOR3X1_3/B vdd NAND3X1
XFILL_50_6_1 gnd vdd FILL
XOAI21X1_105 BUFX4_193/Y BUFX4_478/Y INVX1_399/A gnd OAI21X1_106/C vdd OAI21X1
XOAI21X1_138 BUFX4_121/Y BUFX4_395/Y INVX1_400/A gnd OAI21X1_139/C vdd OAI21X1
XOAI21X1_127 BUFX4_58/Y BUFX4_397/Y OAI21X1_839/B gnd OAI21X1_127/Y vdd OAI21X1
XOAI21X1_116 MUX2X1_58/A NAND2X1_39/Y OAI21X1_116/C gnd OAI21X1_116/Y vdd OAI21X1
XOAI21X1_149 BUFX4_381/Y NAND2X1_51/Y OAI21X1_148/Y gnd OAI21X1_149/Y vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd pedestrian_Hori_Street vdd BUFX2
XNAND2X1_100 AND2X2_2/B BUFX4_174/Y gnd NAND3X1_5/C vdd NAND2X1
XNAND2X1_144 NAND2X1_144/A INVX1_205/Y gnd INVX2_25/A vdd NAND2X1
XNAND2X1_133 INVX4_8/Y NOR2X1_321/B gnd INVX1_197/A vdd NAND2X1
XNAND2X1_122 ped_Hori_Interrupt NAND2X1_122/B gnd INVX4_10/A vdd NAND2X1
XNAND2X1_111 traffic_Street_0[1] AND2X2_5/B gnd NAND2X1_111/Y vdd NAND2X1
XNAND2X1_155 INVX4_9/A INVX4_10/Y gnd NOR2X1_336/A vdd NAND2X1
XNAND2X1_177 AND2X2_27/A NAND2X1_177/B gnd OAI21X1_589/C vdd NAND2X1
XNAND2X1_166 INVX1_215/Y AND2X2_16/A gnd NOR2X1_357/B vdd NAND2X1
XNAND2X1_188 BUFX4_283/Y NOR2X1_723/A gnd NAND2X1_188/Y vdd NAND2X1
XNAND2X1_199 NOR2X1_261/A BUFX4_236/Y gnd OAI21X1_642/C vdd NAND2X1
XFILL_41_6_1 gnd vdd FILL
XFILL_40_1_0 gnd vdd FILL
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_650 INVX1_281/Y BUFX4_249/Y OAI21X1_650/C gnd MUX2X1_197/B vdd OAI21X1
XAOI21X1_3 BUFX4_64/Y NOR2X1_16/Y AOI21X1_3/C gnd AOI21X1_3/Y vdd AOI21X1
XOAI21X1_683 MUX2X1_89/B BUFX4_280/Y NAND2X1_214/Y gnd MUX2X1_200/B vdd OAI21X1
XOAI21X1_661 OAI21X1_661/A BUFX4_261/Y INVX8_32/A gnd OAI22X1_10/B vdd OAI21X1
XOAI21X1_672 OAI21X1_671/Y AND2X2_25/Y OAI21X1_672/C gnd OAI21X1_672/Y vdd OAI21X1
XOAI21X1_694 INVX1_288/Y BUFX4_223/Y NAND2X1_221/Y gnd MUX2X1_204/A vdd OAI21X1
XMUX2X1_150 INVX1_163/Y BUFX4_209/Y MUX2X1_9/S gnd MUX2X1_150/Y vdd MUX2X1
XMUX2X1_161 INVX1_174/Y BUFX4_473/Y MUX2X1_18/S gnd MUX2X1_161/Y vdd MUX2X1
XMUX2X1_183 MUX2X1_183/A MUX2X1_183/B BUFX4_103/Y gnd MUX2X1_183/Y vdd MUX2X1
XMUX2X1_172 MUX2X1_61/B INVX1_186/Y MUX2X1_31/S gnd MUX2X1_172/Y vdd MUX2X1
XMUX2X1_194 MUX2X1_194/A MUX2X1_194/B BUFX4_114/Y gnd MUX2X1_194/Y vdd MUX2X1
XFILL_49_7_1 gnd vdd FILL
XFILL_48_2_0 gnd vdd FILL
XBUFX2_10 BUFX2_10/A gnd west_East[1] vdd BUFX2
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XFILL_32_6_1 gnd vdd FILL
XFILL_31_1_0 gnd vdd FILL
XNOR2X1_1 INVX2_4/A NOR2X1_1/B gnd INVX1_1/A vdd NOR2X1
XFILL_39_2_0 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_44 BUFX4_466/Y NOR2X1_83/B NOR2X1_83/Y gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_33 BUFX4_173/Y NOR2X1_65/Y NOR2X1_67/Y gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_11 MUX2X1_8/B NOR2X1_30/B NOR2X1_31/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_22 BUFX4_316/Y NOR2X1_47/B NOR2X1_48/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_55 MUX2X1_66/B NOR2X1_97/B NOR2X1_100/Y gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_77 MUX2X1_86/B MUX2X1_88/S NOR2X1_133/Y gnd AOI21X1_77/Y vdd AOI21X1
XAOI21X1_66 BUFX4_216/Y NAND2X1_50/B NOR2X1_118/Y gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_99 AND2X2_2/B NOR2X1_167/B AOI21X1_99/C gnd AOI21X1_99/Y vdd AOI21X1
XAOI21X1_88 BUFX4_467/Y MUX2X1_94/S AOI21X1_88/C gnd AOI21X1_88/Y vdd AOI21X1
XOAI21X1_6 BUFX4_442/Y OAI21X1_7/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XBUFX4_308 INVX8_26/Y gnd BUFX4_308/Y vdd BUFX4
XFILL_6_7_1 gnd vdd FILL
XFILL_5_2_0 gnd vdd FILL
XBUFX4_319 INVX8_1/Y gnd AND2X2_6/B vdd BUFX4
XFILL_13_1_0 gnd vdd FILL
XFILL_14_6_1 gnd vdd FILL
XOAI22X1_30 NOR2X1_456/Y OAI22X1_30/B OAI22X1_30/C NOR2X1_455/Y gnd OAI22X1_30/Y vdd
+ OAI22X1
XOAI22X1_52 NOR2X1_529/Y OAI22X1_52/B OAI22X1_52/C NOR2X1_526/Y gnd OAI22X1_52/Y vdd
+ OAI22X1
XOAI22X1_41 OAI22X1_41/A OAI22X1_41/B OAI22X1_41/C NOR2X1_494/Y gnd OAI22X1_41/Y vdd
+ OAI22X1
XOAI22X1_63 OAI22X1_63/A OAI22X1_63/B OAI22X1_63/C OAI22X1_63/D gnd OAI22X1_63/Y vdd
+ OAI22X1
XOAI22X1_85 OAI22X1_85/A OAI22X1_85/B OAI22X1_85/C OAI22X1_85/D gnd OAI22X1_85/Y vdd
+ OAI22X1
XOAI22X1_74 OAI22X1_74/A OAI22X1_74/B OAI22X1_74/C OAI22X1_74/D gnd OAI22X1_74/Y vdd
+ OAI22X1
XOAI21X1_1209 INVX1_113/Y AND2X2_36/B BUFX4_151/Y gnd AOI21X1_499/C vdd OAI21X1
XOAI21X1_480 BUFX4_305/Y OAI22X1_2/D INVX2_21/A gnd NAND3X1_39/A vdd OAI21X1
XOAI21X1_491 NOR2X1_328/Y NAND3X1_39/A INVX1_198/A gnd AOI21X1_227/C vdd OAI21X1
XAOI21X1_515 BUFX4_426/Y NOR2X1_57/Y NOR2X1_627/Y gnd AOI21X1_515/Y vdd AOI21X1
XAOI21X1_504 NAND2X1_97/A BUFX4_230/Y AOI21X1_504/C gnd AOI21X1_504/Y vdd AOI21X1
XAOI21X1_559 BUFX4_441/Y NOR2X1_137/B NOR2X1_671/Y gnd AOI21X1_559/Y vdd AOI21X1
XAOI21X1_548 BUFX4_69/Y AOI21X1_62/B NOR2X1_660/Y gnd AOI21X1_548/Y vdd AOI21X1
XAOI21X1_526 BUFX4_66/Y NOR2X1_76/B NOR2X1_638/Y gnd AOI21X1_526/Y vdd AOI21X1
XAOI21X1_537 BUFX4_324/Y NOR2X1_92/B NOR2X1_649/Y gnd AOI21X1_537/Y vdd AOI21X1
XBUFX4_127 INVX8_20/Y gnd BUFX4_127/Y vdd BUFX4
XBUFX4_116 BUFX4_87/A gnd BUFX4_116/Y vdd BUFX4
XBUFX4_105 BUFX4_87/A gnd AND2X2_32/B vdd BUFX4
XFILL_46_5_1 gnd vdd FILL
XBUFX4_149 INVX8_32/Y gnd BUFX4_149/Y vdd BUFX4
XBUFX4_138 INVX8_22/Y gnd BUFX4_138/Y vdd BUFX4
XNOR2X1_209 NOR2X1_209/A MUX2X1_369/S gnd NOR2X1_209/Y vdd NOR2X1
XFILL_45_0_0 gnd vdd FILL
XOAI21X1_1006 INVX1_92/Y BUFX4_257/Y NAND2X1_303/Y gnd MUX2X1_243/B vdd OAI21X1
XOAI21X1_1028 INVX1_79/Y BUFX4_273/Y NAND2X1_311/Y gnd MUX2X1_248/B vdd OAI21X1
XOAI21X1_1017 NOR2X1_76/A BUFX4_266/Y AOI21X1_435/Y gnd NAND3X1_79/B vdd OAI21X1
XOAI21X1_1039 INVX1_177/Y BUFX4_287/Y NAND2X1_318/Y gnd AOI21X1_447/B vdd OAI21X1
XDFFPOSX1_629 NOR2X1_19/A CLKBUF1_91/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_618 INVX1_26/A CLKBUF1_76/Y MUX2X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_607 INVX1_12/A CLKBUF1_81/Y MUX2X1_9/Y gnd vdd DFFPOSX1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XINVX1_330 INVX1_330/A gnd INVX1_330/Y vdd INVX1
XINVX1_341 INVX1_341/A gnd INVX1_341/Y vdd INVX1
XINVX1_396 INVX1_396/A gnd INVX1_396/Y vdd INVX1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XINVX1_374 INVX1_374/A gnd INVX1_374/Y vdd INVX1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XFILL_37_5_1 gnd vdd FILL
XFILL_36_0_0 gnd vdd FILL
XNOR2X1_710 NOR2X1_710/A NOR2X1_707/B gnd NOR2X1_710/Y vdd NOR2X1
XNOR2X1_732 NOR2X1_732/A NOR2X1_733/B gnd NOR2X1_732/Y vdd NOR2X1
XNOR2X1_721 NOR2X1_721/A NOR2X1_231/B gnd NOR2X1_721/Y vdd NOR2X1
XAOI21X1_312 INVX1_69/Y BUFX4_362/Y BUFX4_156/Y gnd OAI21X1_713/C vdd AOI21X1
XAOI21X1_301 INVX1_141/Y BUFX4_329/Y BUFX4_150/Y gnd AOI21X1_301/Y vdd AOI21X1
XFILL_20_4_1 gnd vdd FILL
XAOI21X1_323 BUFX4_261/Y INVX1_446/A OAI21X1_737/Y gnd OAI21X1_739/A vdd AOI21X1
XAOI21X1_334 BUFX4_148/Y OAI21X1_753/Y AOI21X1_333/Y gnd AOI21X1_334/Y vdd AOI21X1
XAOI21X1_356 INVX1_331/Y BUFX4_343/Y BUFX4_159/Y gnd OAI21X1_816/C vdd AOI21X1
XAOI21X1_345 BUFX4_155/Y OAI21X1_790/Y AOI21X1_344/Y gnd MUX2X1_215/A vdd AOI21X1
XAOI21X1_367 BUFX4_101/Y OAI21X1_838/Y AOI21X1_367/C gnd AOI21X1_367/Y vdd AOI21X1
XAOI21X1_378 AOI21X1_378/A BUFX4_410/Y BUFX4_274/Y gnd OAI21X1_858/C vdd AOI21X1
XDFFPOSX1_11 NOR2X1_453/A CLKBUF1_14/Y AOI21X1_164/Y gnd vdd DFFPOSX1
XAOI21X1_389 BUFX4_32/Y AOI21X1_389/B BUFX4_165/Y gnd AOI21X1_389/Y vdd AOI21X1
XDFFPOSX1_33 NOR2X1_274/A CLKBUF1_19/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_22 NOR2X1_266/A CLKBUF1_72/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XOAI21X1_1540 BUFX4_424/Y NAND2X1_81/Y OAI21X1_1540/C gnd OAI21X1_1540/Y vdd OAI21X1
XDFFPOSX1_44 NOR2X1_509/A CLKBUF1_98/Y OAI21X1_370/Y gnd vdd DFFPOSX1
XOAI21X1_1562 BUFX4_442/Y NAND2X1_85/Y OAI21X1_1561/Y gnd DFFPOSX1_587/D vdd OAI21X1
XDFFPOSX1_77 NOR2X1_604/A CLKBUF1_21/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_171/A CLKBUF1_96/Y MUX2X1_158/Y gnd vdd DFFPOSX1
XOAI21X1_1551 BUFX4_385/Y BUFX4_195/Y DFFPOSX1_570/Q gnd OAI21X1_1552/C vdd OAI21X1
XDFFPOSX1_55 INVX1_160/A CLKBUF1_40/Y MUX2X1_147/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 NOR2X1_280/A CLKBUF1_91/Y AOI21X1_183/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 OAI21X1_868/A CLKBUF1_47/Y OAI21X1_400/Y gnd vdd DFFPOSX1
XFILL_28_5_1 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_404 INVX1_188/A CLKBUF1_3/Y OAI21X1_528/Y gnd vdd DFFPOSX1
XDFFPOSX1_426 NAND2X1_158/A CLKBUF1_3/Y AND2X2_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_437 INVX1_3/A CLKBUF1_17/Y NOR2X1_362/Y gnd vdd DFFPOSX1
XDFFPOSX1_415 OAI21X1_754/B CLKBUF1_33/Y DFFPOSX1_415/D gnd vdd DFFPOSX1
XDFFPOSX1_448 INVX1_315/A CLKBUF1_102/Y MUX2X1_362/Y gnd vdd DFFPOSX1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XDFFPOSX1_459 INVX1_260/A CLKBUF1_83/Y MUX2X1_365/Y gnd vdd DFFPOSX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XNOR2X1_551 NOR2X1_551/A BUFX4_363/Y gnd NOR2X1_551/Y vdd NOR2X1
XNOR2X1_540 NOR2X1_665/A BUFX4_327/Y gnd NOR2X1_540/Y vdd NOR2X1
XNOR2X1_562 AND2X2_48/B NOR2X1_562/B gnd OAI22X1_66/B vdd NOR2X1
XNOR2X1_595 NOR2X1_595/A INVX8_31/A gnd NOR2X1_595/Y vdd NOR2X1
XNOR2X1_573 BUFX4_415/Y OAI22X1_67/Y gnd NOR2X1_573/Y vdd NOR2X1
XNOR2X1_584 BUFX4_40/Y NOR2X1_584/B gnd OAI22X1_75/D vdd NOR2X1
XAOI21X1_131 MUX2X1_66/B MUX2X1_369/S NOR2X1_209/Y gnd AOI21X1_131/Y vdd AOI21X1
XAOI21X1_120 BUFX4_377/Y MUX2X1_364/S NOR2X1_194/Y gnd AOI21X1_120/Y vdd AOI21X1
XAOI21X1_142 BUFX4_380/Y NOR2X1_716/B NOR2X1_225/Y gnd AOI21X1_142/Y vdd AOI21X1
XAOI21X1_164 MUX2X1_40/B MUX2X1_400/S NOR2X1_258/Y gnd AOI21X1_164/Y vdd AOI21X1
XAOI21X1_175 BUFX4_178/Y MUX2X1_410/S NOR2X1_272/Y gnd DFFPOSX1_31/D vdd AOI21X1
XAOI21X1_153 BUFX4_176/Y NOR2X1_727/B NOR2X1_242/Y gnd AOI21X1_153/Y vdd AOI21X1
XAOI21X1_186 BUFX4_178/Y NOR2X1_30/B NOR2X1_283/Y gnd AOI21X1_186/Y vdd AOI21X1
XAOI21X1_197 BUFX4_209/Y NOR2X1_47/B NOR2X1_294/Y gnd AOI21X1_197/Y vdd AOI21X1
XDFFPOSX1_960 NOR2X1_198/A CLKBUF1_4/Y AOI21X1_123/Y gnd vdd DFFPOSX1
XOAI21X1_1381 NAND2X1_57/Y BUFX4_321/Y OAI21X1_1380/Y gnd DFFPOSX1_273/D vdd OAI21X1
XOAI21X1_1370 BUFX4_130/Y BUFX4_297/Y INVX1_353/A gnd OAI21X1_1370/Y vdd OAI21X1
XOAI21X1_1392 BUFX4_387/Y BUFX4_403/Y INVX1_311/A gnd OAI21X1_1392/Y vdd OAI21X1
XDFFPOSX1_993 AOI21X1_455/A CLKBUF1_7/Y OAI21X1_277/Y gnd vdd DFFPOSX1
XDFFPOSX1_971 INVX1_131/A CLKBUF1_46/Y MUX2X1_118/Y gnd vdd DFFPOSX1
XDFFPOSX1_982 NOR2X1_212/A CLKBUF1_1/Y AOI21X1_133/Y gnd vdd DFFPOSX1
XFILL_43_3_1 gnd vdd FILL
XFILL_34_3_1 gnd vdd FILL
XFILL_20_2 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XOAI21X1_309 BUFX4_381/Y NAND2X1_77/Y OAI21X1_309/C gnd OAI21X1_309/Y vdd OAI21X1
XDFFPOSX1_201 NOR2X1_686/A CLKBUF1_101/Y AOI21X1_574/Y gnd vdd DFFPOSX1
XBUFX4_7 clock gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_212 AND2X2_39/B CLKBUF1_22/Y DFFPOSX1_212/D gnd vdd DFFPOSX1
XDFFPOSX1_245 INVX1_459/A CLKBUF1_41/Y MUX2X1_353/Y gnd vdd DFFPOSX1
XDFFPOSX1_223 NOR2X1_647/A CLKBUF1_65/Y AOI21X1_535/Y gnd vdd DFFPOSX1
XDFFPOSX1_234 INVX1_228/A CLKBUF1_20/Y MUX2X1_294/Y gnd vdd DFFPOSX1
XDFFPOSX1_267 AND2X2_29/B CLKBUF1_61/Y AOI21X1_587/Y gnd vdd DFFPOSX1
XDFFPOSX1_289 AOI21X1_476/B CLKBUF1_31/Y OAI21X1_1373/Y gnd vdd DFFPOSX1
XDFFPOSX1_278 INVX1_244/A CLKBUF1_69/Y MUX2X1_329/Y gnd vdd DFFPOSX1
XDFFPOSX1_256 NOR2X1_673/A CLKBUF1_93/Y AOI21X1_561/Y gnd vdd DFFPOSX1
XNAND2X1_326 OAI21X1_260/C BUFX4_359/Y gnd NAND2X1_326/Y vdd NAND2X1
XNAND2X1_304 NOR2X1_123/A BUFX4_258/Y gnd NAND2X1_304/Y vdd NAND2X1
XNAND2X1_315 NOR2X1_108/A BUFX4_281/Y gnd NAND2X1_315/Y vdd NAND2X1
XNAND2X1_348 OAI21X1_310/C BUFX4_249/Y gnd NAND2X1_348/Y vdd NAND2X1
XNAND2X1_359 traffic_Street_0[2] NOR2X1_188/B gnd NAND2X1_359/Y vdd NAND2X1
XNAND2X1_337 NAND2X1_337/A NAND2X1_337/B gnd NOR2X1_562/B vdd NAND2X1
XNOR3X1_11 INVX2_20/Y INVX2_25/Y OAI22X1_2/C gnd NOR3X1_11/Y vdd NOR3X1
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XNOR2X1_370 BUFX4_89/Y NOR2X1_370/B gnd NOR2X1_371/A vdd NOR2X1
XNOR2X1_392 NOR2X1_121/A BUFX4_327/Y gnd OAI22X1_13/A vdd NOR2X1
XNOR2X1_381 NOR2X1_381/A BUFX4_258/Y gnd OAI22X1_9/D vdd NOR2X1
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XOAI21X1_821 BUFX4_351/Y INVX1_41/A BUFX4_154/Y gnd OAI21X1_821/Y vdd OAI21X1
XOAI21X1_832 OAI21X1_831/Y AND2X2_31/Y BUFX4_414/Y gnd OAI22X1_25/D vdd OAI21X1
XOAI21X1_810 NOR2X1_50/A AND2X2_52/A BUFX4_89/Y gnd OAI22X1_23/B vdd OAI21X1
XOAI21X1_865 INVX1_179/A BUFX4_349/Y AOI21X1_381/Y gnd OAI21X1_866/C vdd OAI21X1
XOAI21X1_876 OAI21X1_876/A BUFX4_288/Y BUFX4_118/Y gnd OAI22X1_29/B vdd OAI21X1
XOAI21X1_854 INVX1_98/Y BUFX4_34/Y BUFX4_273/Y gnd OAI21X1_854/Y vdd OAI21X1
XOAI21X1_843 INVX1_109/Y BUFX4_268/Y OAI21X1_843/C gnd AOI21X1_372/B vdd OAI21X1
XOAI21X1_898 OAI21X1_898/A AND2X2_51/B BUFX4_81/Y gnd OAI22X1_32/B vdd OAI21X1
XOAI21X1_887 INVX1_146/Y BUFX4_227/Y OAI21X1_887/C gnd MUX2X1_226/A vdd OAI21X1
XMUX2X1_321 INVX1_251/Y BUFX4_439/Y MUX2X1_81/S gnd MUX2X1_321/Y vdd MUX2X1
XMUX2X1_332 BUFX4_441/Y INVX1_246/Y MUX2X1_89/S gnd MUX2X1_332/Y vdd MUX2X1
XMUX2X1_310 INVX1_296/Y MUX2X1_18/B MUX2X1_71/S gnd MUX2X1_310/Y vdd MUX2X1
XMUX2X1_354 BUFX4_437/Y INVX1_239/Y MUX2X1_108/S gnd MUX2X1_354/Y vdd MUX2X1
XMUX2X1_343 INVX1_307/Y BUFX4_430/Y MUX2X1_97/S gnd MUX2X1_343/Y vdd MUX2X1
XMUX2X1_365 INVX1_260/Y BUFX4_444/Y MUX2X1_366/S gnd MUX2X1_365/Y vdd MUX2X1
XMUX2X1_376 BUFX4_70/Y INVX1_377/Y MUX2X1_376/S gnd MUX2X1_376/Y vdd MUX2X1
XMUX2X1_398 BUFX4_441/Y INVX1_268/Y MUX2X1_400/S gnd MUX2X1_398/Y vdd MUX2X1
XMUX2X1_387 BUFX4_67/Y INVX1_384/Y NOR2X1_233/Y gnd MUX2X1_387/Y vdd MUX2X1
XDFFPOSX1_790 INVX1_84/A CLKBUF1_63/Y MUX2X1_74/Y gnd vdd DFFPOSX1
XFILL_8_4_1 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_106 BUFX4_381/Y NAND2X1_37/Y OAI21X1_106/C gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_128 MUX2X1_77/B NAND2X1_44/Y OAI21X1_127/Y gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_117 BUFX4_449/Y BUFX4_54/Y NOR2X1_408/A gnd OAI21X1_117/Y vdd OAI21X1
XOAI21X1_139 NAND2X1_48/Y BUFX4_371/Y OAI21X1_139/C gnd OAI21X1_139/Y vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd pedestrian_Vert_Street vdd BUFX2
XNAND2X1_101 traffic_Street_1[0] traffic_Street_1[1] gnd NAND3X1_5/B vdd NAND2X1
XNAND2X1_134 INVX2_22/Y NOR3X1_9/Y gnd AOI21X1_225/A vdd NAND2X1
XNAND2X1_112 OAI21X1_451/Y NAND3X1_16/Y gnd NOR3X1_6/A vdd NAND2X1
XNAND2X1_123 NOR3X1_1/B INVX1_189/Y gnd NAND2X1_123/Y vdd NAND2X1
XNAND2X1_156 NAND3X1_61/Y NAND3X1_59/Y gnd NAND2X1_156/Y vdd NAND2X1
XNAND2X1_145 INVX2_25/A AOI22X1_9/C gnd OAI21X1_502/C vdd NAND2X1
XNAND2X1_167 NAND2X1_167/A NAND3X1_69/Y gnd NAND2X1_167/Y vdd NAND2X1
XNAND2X1_178 BUFX4_34/Y AOI21X1_271/Y gnd AOI22X1_13/B vdd NAND2X1
XNAND2X1_189 NOR2X1_17/A BUFX4_290/Y gnd NAND2X1_189/Y vdd NAND2X1
XFILL_40_1_1 gnd vdd FILL
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XOAI21X1_640 INVX1_151/Y BUFX4_233/Y OAI21X1_640/C gnd MUX2X1_192/B vdd OAI21X1
XOAI21X1_651 INVX1_184/Y BUFX4_251/Y OAI21X1_651/C gnd MUX2X1_197/A vdd OAI21X1
XOAI21X1_684 MUX2X1_92/B BUFX4_282/Y OAI21X1_684/C gnd MUX2X1_200/A vdd OAI21X1
XAOI21X1_4 MUX2X1_8/B NOR2X1_16/Y AOI21X1_4/C gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_662 INVX1_137/A BUFX4_263/Y OAI21X1_662/C gnd NAND3X1_73/B vdd OAI21X1
XOAI21X1_673 INVX1_131/Y BUFX4_271/Y BUFX4_147/Y gnd AOI21X1_305/C vdd OAI21X1
XOAI21X1_695 BUFX4_345/Y NOR2X1_170/A BUFX4_152/Y gnd OAI22X1_15/C vdd OAI21X1
XMUX2X1_140 INVX1_153/Y BUFX4_372/Y MUX2X1_406/S gnd MUX2X1_140/Y vdd MUX2X1
XMUX2X1_173 OR2X2_1/Y AND2X2_3/A traffic_Street_1[3] gnd AND2X2_2/A vdd MUX2X1
XMUX2X1_162 INVX1_175/Y BUFX4_209/Y MUX2X1_21/S gnd MUX2X1_162/Y vdd MUX2X1
XMUX2X1_151 INVX1_164/Y BUFX4_178/Y MUX2X1_9/S gnd MUX2X1_151/Y vdd MUX2X1
XMUX2X1_195 MUX2X1_195/A MUX2X1_195/B BUFX4_115/Y gnd MUX2X1_195/Y vdd MUX2X1
XMUX2X1_184 MUX2X1_184/A MUX2X1_184/B BUFX4_104/Y gnd MUX2X1_186/B vdd MUX2X1
XFILL_48_2_1 gnd vdd FILL
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XFILL_31_1_1 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A INVX1_1/Y gnd NOR2X1_2/Y vdd NOR2X1
XFILL_39_2_1 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_34 BUFX4_372/Y NOR2X1_65/Y NOR2X1_68/Y gnd AOI21X1_34/Y vdd AOI21X1
XAOI21X1_12 MUX2X1_1/B NOR2X1_33/Y NOR2X1_34/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_23 MUX2X1_6/B MUX2X1_31/S NOR2X1_50/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_45 BUFX4_469/Y NOR2X1_85/B NOR2X1_85/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_67 MUX2X1_83/B NAND2X1_50/B NOR2X1_119/Y gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_56 MUX2X1_71/B MUX2X1_75/S NOR2X1_103/Y gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_78 MUX2X1_83/B MUX2X1_88/S AOI21X1_78/C gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_89 MUX2X1_44/A MUX2X1_96/S NOR2X1_151/Y gnd AOI21X1_89/Y vdd AOI21X1
XOAI21X1_7 MUX2X1_18/B OAI21X1_7/B OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XFILL_5_2_1 gnd vdd FILL
XBUFX4_309 INVX8_26/Y gnd BUFX4_309/Y vdd BUFX4
XFILL_42_9_0 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XOAI22X1_20 NOR2X1_423/Y OAI22X1_20/B OAI22X1_20/C NOR2X1_422/Y gnd OAI22X1_20/Y vdd
+ OAI22X1
XOAI22X1_42 OAI22X1_42/A OAI22X1_42/B OAI22X1_42/C INVX4_14/Y gnd OAI22X1_42/Y vdd
+ OAI22X1
XOAI22X1_31 NOR2X1_460/Y OAI22X1_31/B OAI22X1_31/C NOR2X1_459/Y gnd OAI22X1_31/Y vdd
+ OAI22X1
XOAI22X1_64 OAI22X1_64/A OAI22X1_64/B OAI22X1_64/C OAI22X1_64/D gnd OAI22X1_64/Y vdd
+ OAI22X1
XOAI22X1_75 NOR2X1_587/Y OAI22X1_75/B OAI22X1_75/C OAI22X1_75/D gnd NOR2X1_590/B vdd
+ OAI22X1
XOAI22X1_53 NOR2X1_534/Y OAI22X1_53/B OAI22X1_53/C NOR2X1_533/Y gnd OAI22X1_53/Y vdd
+ OAI22X1
XOAI22X1_86 BUFX4_206/Y MUX2X1_263/Y OAI22X1_86/C OAI22X1_86/D gnd OAI22X1_86/Y vdd
+ OAI22X1
XOAI21X1_492 OAI21X1_492/A AOI21X1_241/C INVX1_199/A gnd NOR2X1_336/B vdd OAI21X1
XOAI21X1_470 NOR3X1_1/B NAND2X1_116/Y NAND2X1_123/Y gnd NAND3X1_29/C vdd OAI21X1
XOAI21X1_481 AND2X2_6/B NOR2X1_308/B NAND3X1_15/C gnd XOR2X1_1/B vdd OAI21X1
XFILL_33_9_0 gnd vdd FILL
XAOI21X1_516 MUX2X1_4/B NOR2X1_57/Y NOR2X1_628/Y gnd AOI21X1_516/Y vdd AOI21X1
XAOI21X1_505 NAND2X1_93/A BUFX4_343/Y BUFX4_159/Y gnd AOI21X1_505/Y vdd AOI21X1
XAOI21X1_538 BUFX4_444/Y NOR2X1_97/B NOR2X1_650/Y gnd AOI21X1_538/Y vdd AOI21X1
XAOI21X1_527 BUFX4_324/Y NOR2X1_76/B NOR2X1_639/Y gnd AOI21X1_527/Y vdd AOI21X1
XAOI21X1_549 BUFX4_316/Y AOI21X1_62/B NOR2X1_661/Y gnd AOI21X1_549/Y vdd AOI21X1
XFILL_24_9_0 gnd vdd FILL
XBUFX4_128 INVX8_20/Y gnd BUFX4_128/Y vdd BUFX4
XBUFX4_117 BUFX4_87/A gnd BUFX4_117/Y vdd BUFX4
XBUFX4_106 BUFX4_82/A gnd BUFX4_106/Y vdd BUFX4
XBUFX4_139 INVX8_22/Y gnd BUFX4_139/Y vdd BUFX4
XFILL_45_0_1 gnd vdd FILL
XFILL_15_9_0 gnd vdd FILL
XOAI21X1_1007 INVX1_395/Y BUFX4_259/Y NAND2X1_304/Y gnd MUX2X1_243/A vdd OAI21X1
XOAI21X1_1018 NOR2X1_82/A BUFX4_345/Y AOI21X1_436/Y gnd NAND3X1_79/C vdd OAI21X1
XDFFPOSX1_619 NAND2X1_11/A CLKBUF1_76/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_608 INVX1_15/A CLKBUF1_47/Y MUX2X1_10/Y gnd vdd DFFPOSX1
XOAI21X1_1029 INVX1_83/Y BUFX4_275/Y NAND2X1_312/Y gnd MUX2X1_248/A vdd OAI21X1
XINVX1_331 INVX1_331/A gnd INVX1_331/Y vdd INVX1
XINVX1_353 INVX1_353/A gnd INVX1_353/Y vdd INVX1
XINVX1_342 INVX1_342/A gnd INVX1_342/Y vdd INVX1
XINVX1_320 INVX1_320/A gnd INVX1_320/Y vdd INVX1
XINVX1_386 INVX1_386/A gnd INVX1_386/Y vdd INVX1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XINVX1_397 INVX1_397/A gnd INVX1_397/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XNOR2X1_711 NOR2X1_711/A MUX2X1_369/S gnd NOR2X1_711/Y vdd NOR2X1
XFILL_43_1 gnd vdd FILL
XNOR2X1_700 NOR2X1_700/A INVX1_219/A gnd NOR2X1_700/Y vdd NOR2X1
XFILL_36_0_1 gnd vdd FILL
XNOR2X1_733 NOR2X1_733/A NOR2X1_733/B gnd NOR2X1_733/Y vdd NOR2X1
XNOR2X1_722 NOR2X1_564/A NOR2X1_231/B gnd NOR2X1_722/Y vdd NOR2X1
XAOI21X1_302 INVX8_29/A OAI21X1_659/Y NOR2X1_385/Y gnd OAI22X1_12/C vdd AOI21X1
XAOI21X1_324 BUFX4_263/Y NOR2X1_641/A AOI21X1_324/C gnd OAI21X1_739/B vdd AOI21X1
XAOI21X1_313 BUFX4_33/Y MUX2X1_206/Y AOI21X1_313/C gnd NOR2X1_411/B vdd AOI21X1
XAOI21X1_346 INVX8_28/A MUX2X1_216/Y BUFX4_401/Y gnd AOI21X1_346/Y vdd AOI21X1
XAOI21X1_357 INVX4_14/Y AOI21X1_339/Y AOI21X1_357/C gnd AOI21X1_392/C vdd AOI21X1
XAOI21X1_335 BUFX4_367/Y INVX1_311/Y BUFX4_148/Y gnd OAI21X1_756/C vdd AOI21X1
XAOI21X1_379 MUX2X1_94/B BUFX4_278/Y AOI21X1_379/C gnd AOI21X1_379/Y vdd AOI21X1
XAOI21X1_368 INVX1_78/Y BUFX4_358/Y AOI21X1_368/C gnd OAI21X1_841/A vdd AOI21X1
XDFFPOSX1_45 NAND2X1_89/A CLKBUF1_40/Y DFFPOSX1_45/D gnd vdd DFFPOSX1
XOAI21X1_1541 BUFX4_194/Y BUFX4_308/Y NAND2X1_292/B gnd OAI21X1_1542/C vdd OAI21X1
XDFFPOSX1_12 INVX1_150/A CLKBUF1_31/Y MUX2X1_137/Y gnd vdd DFFPOSX1
XOAI21X1_1530 NAND2X1_80/Y BUFX4_440/Y OAI21X1_1530/C gnd DFFPOSX1_543/D vdd OAI21X1
XDFFPOSX1_23 NOR2X1_454/A CLKBUF1_14/Y AOI21X1_171/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX1_276/A CLKBUF1_11/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XOAI21X1_1563 BUFX4_188/Y BUFX4_195/Y OAI21X1_797/B gnd OAI21X1_1563/Y vdd OAI21X1
XOAI21X1_1552 NAND2X1_82/Y BUFX4_321/Y OAI21X1_1552/C gnd DFFPOSX1_570/D vdd OAI21X1
XDFFPOSX1_78 NOR2X1_275/A CLKBUF1_66/Y AOI21X1_178/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 INVX1_161/A CLKBUF1_73/Y MUX2X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_172/A CLKBUF1_78/Y MUX2X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 NOR2X1_281/A CLKBUF1_30/Y AOI21X1_184/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_47_8_0 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XDFFPOSX1_427 NAND2X1_147/A CLKBUF1_3/Y NAND2X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_405 XNOR2X1_1/B CLKBUF1_3/Y AOI22X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_438 INVX2_3/A CLKBUF1_79/Y OAI21X1_551/Y gnd vdd DFFPOSX1
XDFFPOSX1_416 MUX2X1_230/A CLKBUF1_12/Y OAI21X1_1419/Y gnd vdd DFFPOSX1
XDFFPOSX1_449 INVX1_381/A CLKBUF1_9/Y MUX2X1_363/Y gnd vdd DFFPOSX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XINVX1_194 NOR3X1_5/A gnd INVX1_194/Y vdd INVX1
XFILL_38_8_0 gnd vdd FILL
XBUFX4_470 INVX8_15/Y gnd BUFX4_470/Y vdd BUFX4
XNOR2X1_552 NAND2X1_3/A BUFX4_227/Y gnd OAI22X1_61/D vdd NOR2X1
XNOR2X1_541 BUFX4_416/Y NOR2X1_541/B gnd NOR2X1_541/Y vdd NOR2X1
XNOR2X1_530 BUFX4_274/Y NOR2X1_530/B gnd NOR2X1_530/Y vdd NOR2X1
XNOR2X1_563 BUFX4_344/Y INVX1_434/Y gnd NOR2X1_563/Y vdd NOR2X1
XNOR2X1_574 NOR2X1_574/A AND2X2_23/A gnd OAI22X1_68/D vdd NOR2X1
XNOR2X1_585 NOR2X1_585/A BUFX4_282/Y gnd NOR2X1_585/Y vdd NOR2X1
XNOR2X1_596 NOR2X1_596/A BUFX4_325/Y gnd NOR2X1_596/Y vdd NOR2X1
XFILL_21_7_0 gnd vdd FILL
XAOI21X1_121 BUFX4_466/Y MUX2X1_364/S NOR2X1_195/Y gnd AOI21X1_121/Y vdd AOI21X1
XAOI21X1_110 MUX2X1_96/A MUX2X1_108/S NOR2X1_179/Y gnd AOI21X1_110/Y vdd AOI21X1
XAOI21X1_132 BUFX4_177/Y MUX2X1_120/S NOR2X1_211/Y gnd AOI21X1_132/Y vdd AOI21X1
XAOI21X1_176 BUFX4_372/Y MUX2X1_410/S NOR2X1_273/Y gnd AOI21X1_176/Y vdd AOI21X1
XAOI21X1_165 BUFX4_473/Y MUX2X1_400/S NOR2X1_259/Y gnd AOI21X1_165/Y vdd AOI21X1
XAOI21X1_154 BUFX4_381/Y NOR2X1_727/B NOR2X1_243/Y gnd AOI21X1_154/Y vdd AOI21X1
XAOI21X1_143 BUFX4_469/Y NOR2X1_716/B NOR2X1_226/Y gnd AOI21X1_143/Y vdd AOI21X1
XAOI21X1_187 BUFX4_375/Y NOR2X1_30/B NOR2X1_284/Y gnd AOI21X1_187/Y vdd AOI21X1
XAOI21X1_198 MUX2X1_77/B NOR2X1_47/B NOR2X1_295/Y gnd AOI21X1_198/Y vdd AOI21X1
XDFFPOSX1_950 OAI21X1_254/C CLKBUF1_10/Y OAI21X1_255/Y gnd vdd DFFPOSX1
XOAI21X1_1360 BUFX4_454/Y BUFX4_185/Y INVX1_312/A gnd OAI21X1_1361/C vdd OAI21X1
XOAI21X1_1371 NAND2X1_56/Y BUFX4_65/Y OAI21X1_1370/Y gnd OAI21X1_1371/Y vdd OAI21X1
XOAI21X1_1382 BUFX4_133/Y BUFX4_129/Y OAI21X1_587/B gnd OAI21X1_1383/C vdd OAI21X1
XDFFPOSX1_961 NOR2X1_199/A CLKBUF1_82/Y AOI21X1_124/Y gnd vdd DFFPOSX1
XDFFPOSX1_994 OAI21X1_278/C CLKBUF1_7/Y OAI21X1_279/Y gnd vdd DFFPOSX1
XOAI21X1_1393 NAND2X1_59/Y BUFX4_422/Y OAI21X1_1392/Y gnd OAI21X1_1393/Y vdd OAI21X1
XDFFPOSX1_983 NOR2X1_214/A CLKBUF1_83/Y AOI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_972 NOR2X1_466/A CLKBUF1_50/Y AOI21X1_126/Y gnd vdd DFFPOSX1
XFILL_29_8_0 gnd vdd FILL
XFILL_4_8_0 gnd vdd FILL
XFILL_12_7_0 gnd vdd FILL
XDFFPOSX1_202 INVX1_241/A CLKBUF1_59/Y MUX2X1_337/Y gnd vdd DFFPOSX1
XDFFPOSX1_213 AOI21X1_472/A CLKBUF1_29/Y DFFPOSX1_213/D gnd vdd DFFPOSX1
XBUFX4_8 clock gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_246 OAI21X1_587/B CLKBUF1_31/Y DFFPOSX1_246/D gnd vdd DFFPOSX1
XDFFPOSX1_235 INVX1_292/A CLKBUF1_65/Y MUX2X1_295/Y gnd vdd DFFPOSX1
XDFFPOSX1_224 NOR2X1_648/A CLKBUF1_83/Y AOI21X1_536/Y gnd vdd DFFPOSX1
XDFFPOSX1_279 NOR2X1_670/A CLKBUF1_70/Y AOI21X1_558/Y gnd vdd DFFPOSX1
XDFFPOSX1_257 NOR2X1_674/A CLKBUF1_69/Y AOI21X1_562/Y gnd vdd DFFPOSX1
XDFFPOSX1_268 NOR2X1_700/A CLKBUF1_13/Y AOI21X1_588/Y gnd vdd DFFPOSX1
XNAND2X1_327 BUFX4_33/Y OAI22X1_47/Y gnd NAND2X1_327/Y vdd NAND2X1
XNAND2X1_305 NOR2X1_128/A BUFX4_260/Y gnd NAND2X1_305/Y vdd NAND2X1
XNAND2X1_316 NOR2X1_113/A BUFX4_283/Y gnd NAND2X1_316/Y vdd NAND2X1
XNAND2X1_338 BUFX4_248/Y NAND2X1_338/B gnd NAND2X1_338/Y vdd NAND2X1
XNAND2X1_349 NOR2X1_238/A BUFX4_251/Y gnd NAND2X1_349/Y vdd NAND2X1
XNOR3X1_12 NOR3X1_12/A NOR3X1_12/B NOR3X1_12/C gnd NOR3X1_12/Y vdd NOR3X1
XNOR2X1_360 INVX2_8/Y BUFX4_189/Y gnd AND2X2_20/A vdd NOR2X1
XNOR2X1_393 BUFX4_410/Y OAI22X1_13/Y gnd NOR2X1_393/Y vdd NOR2X1
XNOR2X1_382 NOR2X1_246/A BUFX4_336/Y gnd OAI22X1_9/A vdd NOR2X1
XNOR2X1_371 NOR2X1_371/A NOR2X1_371/B gnd NOR2X1_371/Y vdd NOR2X1
XOAI21X1_800 INVX1_24/A AND2X2_51/B BUFX4_86/Y gnd AOI21X1_352/C vdd OAI21X1
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XOAI21X1_822 INVX1_43/Y BUFX4_249/Y NAND2X1_247/Y gnd AOI21X1_359/B vdd OAI21X1
XOAI21X1_811 OAI22X1_23/Y BUFX4_31/Y BUFX4_202/Y gnd OAI22X1_24/B vdd OAI21X1
XOAI21X1_833 INVX1_62/Y BUFX4_256/Y NAND2X1_249/Y gnd MUX2X1_219/B vdd OAI21X1
XOAI21X1_866 NOR2X1_449/Y OAI21X1_864/Y OAI21X1_866/C gnd NOR2X1_450/B vdd OAI21X1
XOAI21X1_855 INVX1_94/Y BUFX4_34/Y BUFX4_327/Y gnd OAI21X1_856/A vdd OAI21X1
XOAI21X1_844 OAI21X1_194/C AND2X2_25/B BUFX4_103/Y gnd OAI21X1_844/Y vdd OAI21X1
XOAI21X1_899 BUFX4_370/Y NOR2X1_198/A BUFX4_156/Y gnd OAI22X1_33/C vdd OAI21X1
XOAI21X1_877 BUFX4_350/Y NOR2X1_272/A BUFX4_146/Y gnd OAI21X1_877/Y vdd OAI21X1
XOAI21X1_888 NOR2X1_457/Y AND2X2_37/Y BUFX4_153/Y gnd OAI21X1_888/Y vdd OAI21X1
XMUX2X1_300 INVX1_416/Y MUX2X1_29/B MUX2X1_59/S gnd MUX2X1_300/Y vdd MUX2X1
XMUX2X1_322 INVX1_313/Y BUFX4_424/Y MUX2X1_81/S gnd MUX2X1_322/Y vdd MUX2X1
XMUX2X1_311 INVX1_345/Y BUFX4_71/Y MUX2X1_71/S gnd MUX2X1_311/Y vdd MUX2X1
XMUX2X1_366 INVX1_316/Y BUFX4_420/Y MUX2X1_366/S gnd MUX2X1_366/Y vdd MUX2X1
XMUX2X1_333 BUFX4_65/Y INVX1_354/Y MUX2X1_89/S gnd MUX2X1_333/Y vdd MUX2X1
XMUX2X1_355 BUFX4_66/Y INVX1_358/Y MUX2X1_108/S gnd MUX2X1_355/Y vdd MUX2X1
XOAI21X1_1190 NOR2X1_105/A BUFX4_358/Y AOI21X1_497/Y gnd OAI21X1_1191/C vdd OAI21X1
XMUX2X1_344 INVX1_357/Y BUFX4_68/Y MUX2X1_97/S gnd MUX2X1_344/Y vdd MUX2X1
XMUX2X1_377 BUFX4_317/Y INVX1_434/Y MUX2X1_376/S gnd MUX2X1_377/Y vdd MUX2X1
XMUX2X1_388 BUFX4_322/Y INVX1_437/Y NOR2X1_233/Y gnd MUX2X1_388/Y vdd MUX2X1
XMUX2X1_399 BUFX4_428/Y INVX1_326/Y MUX2X1_400/S gnd MUX2X1_399/Y vdd MUX2X1
XDFFPOSX1_780 INVX1_78/A CLKBUF1_77/Y MUX2X1_68/Y gnd vdd DFFPOSX1
XDFFPOSX1_791 NOR2X1_410/A CLKBUF1_77/Y AOI21X1_56/Y gnd vdd DFFPOSX1
XFILL_44_6_0 gnd vdd FILL
XFILL_35_6_0 gnd vdd FILL
XOAI21X1_107 BUFX4_193/Y BUFX4_478/Y NOR2X1_569/A gnd OAI21X1_108/C vdd OAI21X1
XOAI21X1_129 BUFX4_58/Y BUFX4_395/Y NAND2X1_311/A gnd OAI21X1_129/Y vdd OAI21X1
XOAI21X1_118 NAND2X1_40/Y MUX2X1_59/B OAI21X1_117/Y gnd OAI21X1_118/Y vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd traffic_Street[0] vdd BUFX2
XNAND2X1_102 AND2X2_3/B AND2X2_3/A gnd NAND3X1_6/C vdd NAND2X1
XNAND2X1_135 INVX1_188/A NOR2X1_321/Y gnd XNOR2X1_1/A vdd NAND2X1
XNAND2X1_124 AND2X2_7/B AND2X2_7/A gnd NOR2X1_311/B vdd NAND2X1
XNAND2X1_113 NAND3X1_17/Y NAND3X1_31/C gnd NOR3X1_6/B vdd NAND2X1
XNAND2X1_146 AND2X2_10/Y NOR3X1_9/Y gnd NAND2X1_146/Y vdd NAND2X1
XNAND2X1_157 NOR2X1_342/Y OAI21X1_483/Y gnd AOI21X1_242/B vdd NAND2X1
XNAND2X1_168 NAND2X1_168/A NOR3X1_7/Y gnd OR2X2_7/B vdd NAND2X1
XNAND2X1_179 BUFX4_258/Y NOR2X1_666/A gnd OAI21X1_591/C vdd NAND2X1
XFILL_26_6_0 gnd vdd FILL
XFILL_1_6_0 gnd vdd FILL
XNOR2X1_190 NOR2X1_190/A NOR2X1_188/B gnd NOR2X1_190/Y vdd NOR2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XOAI21X1_641 INVX1_276/Y BUFX4_235/Y NAND2X1_198/Y gnd MUX2X1_192/A vdd OAI21X1
XOAI21X1_630 INVX1_38/Y AND2X2_37/B OAI21X1_630/C gnd MUX2X1_189/A vdd OAI21X1
XAOI21X1_5 MUX2X1_1/B AOI21X1_7/B AOI21X1_5/C gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_663 NOR2X1_235/A BUFX4_329/Y AOI21X1_301/Y gnd NAND3X1_73/C vdd OAI21X1
XOAI21X1_652 BUFX4_338/Y OAI21X1_413/C BUFX4_158/Y gnd OAI22X1_7/C vdd OAI21X1
XOAI21X1_674 INVX1_133/Y BUFX4_273/Y BUFX4_81/Y gnd AOI21X1_306/C vdd OAI21X1
XOAI21X1_685 BUFX4_361/Y NOR2X1_132/A BUFX4_154/Y gnd OAI22X1_14/C vdd OAI21X1
XOAI21X1_696 OAI21X1_696/A BUFX4_225/Y BUFX4_91/Y gnd OAI22X1_15/B vdd OAI21X1
XMUX2X1_141 INVX1_154/Y BUFX4_473/Y MUX2X1_406/S gnd MUX2X1_141/Y vdd MUX2X1
XMUX2X1_130 MUX2X1_86/B INVX1_143/Y NOR2X1_233/Y gnd MUX2X1_130/Y vdd MUX2X1
XMUX2X1_163 INVX1_176/Y BUFX4_173/Y MUX2X1_21/S gnd MUX2X1_163/Y vdd MUX2X1
XMUX2X1_152 INVX1_165/Y BUFX4_375/Y MUX2X1_9/S gnd MUX2X1_152/Y vdd MUX2X1
XMUX2X1_174 INVX1_189/Y MUX2X1_174/B NOR3X1_1/B gnd NOR3X1_2/C vdd MUX2X1
XFILL_9_7_0 gnd vdd FILL
XMUX2X1_185 MUX2X1_185/A MUX2X1_185/B AND2X2_32/B gnd MUX2X1_185/Y vdd MUX2X1
XMUX2X1_196 MUX2X1_195/Y MUX2X1_194/Y BUFX4_31/Y gnd MUX2X1_196/Y vdd MUX2X1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XFILL_17_6_0 gnd vdd FILL
XNOR2X1_3 INVX1_27/A INVX4_1/Y gnd INVX2_1/A vdd NOR2X1
XFILL_50_4_0 gnd vdd FILL
XAOI21X1_13 BUFX4_64/Y NOR2X1_33/Y NOR2X1_35/Y gnd AOI21X1_13/Y vdd AOI21X1
XAOI21X1_24 BUFX4_214/Y NOR2X1_54/Y NOR2X1_55/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_35 BUFX4_468/Y NOR2X1_65/Y NOR2X1_69/Y gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_46 BUFX4_217/Y MUX2X1_50/S NOR2X1_87/Y gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_68 BUFX4_218/Y MUX2X1_320/S AOI21X1_68/C gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_57 BUFX4_371/Y MUX2X1_75/S AOI21X1_57/C gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_79 BUFX4_214/Y NOR2X1_137/B NOR2X1_136/Y gnd AOI21X1_79/Y vdd AOI21X1
XOAI21X1_8 BUFX4_71/Y OAI21X1_7/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XOAI22X1_32 OAI22X1_32/A OAI22X1_32/B OAI22X1_32/C NOR2X1_461/Y gnd NOR2X1_463/B vdd
+ OAI22X1
XOAI22X1_21 NOR2X1_425/Y OAI22X1_21/B OAI22X1_21/C NOR2X1_424/Y gnd OAI22X1_21/Y vdd
+ OAI22X1
XOAI22X1_10 OAI22X1_10/A OAI22X1_10/B OAI22X1_10/C NOR2X1_383/Y gnd OAI22X1_10/Y vdd
+ OAI22X1
XOAI22X1_43 OAI22X1_43/A OAI22X1_43/B OAI22X1_43/C OAI22X1_43/D gnd MUX2X1_242/B vdd
+ OAI22X1
XFILL_41_4_0 gnd vdd FILL
XFILL_42_9_1 gnd vdd FILL
XOAI22X1_76 NOR2X1_592/Y OAI22X1_76/B OAI22X1_76/C OAI22X1_76/D gnd MUX2X1_262/B vdd
+ OAI22X1
XOAI22X1_65 NOR2X1_559/Y OAI22X1_65/B OAI22X1_65/C AND2X2_50/Y gnd OAI22X1_65/Y vdd
+ OAI22X1
XOAI22X1_54 NOR2X1_537/Y OAI22X1_54/B OAI22X1_54/C NOR2X1_536/Y gnd OAI22X1_54/Y vdd
+ OAI22X1
XOAI22X1_87 NOR2X1_613/Y OAI22X1_87/B OAI22X1_87/C OAI22X1_87/D gnd NOR2X1_614/B vdd
+ OAI22X1
XOAI21X1_482 BUFX4_305/Y INVX4_11/Y INVX2_22/A gnd INVX1_198/A vdd OAI21X1
XOAI21X1_493 NOR2X1_336/B INVX4_10/A AOI22X1_5/D gnd NAND3X1_44/C vdd OAI21X1
XOAI21X1_460 AND2X2_6/B NOR2X1_308/B NAND2X1_116/Y gnd NAND3X1_23/B vdd OAI21X1
XOAI21X1_471 AOI22X1_3/Y INVX1_190/A INVX4_6/Y gnd OAI21X1_471/Y vdd OAI21X1
XFILL_49_5_0 gnd vdd FILL
XFILL_32_4_0 gnd vdd FILL
XFILL_33_9_1 gnd vdd FILL
XAOI21X1_506 NAND2X1_89/A BUFX4_346/Y BUFX4_101/Y gnd AOI21X1_506/Y vdd AOI21X1
XAOI21X1_528 BUFX4_437/Y NOR2X1_83/B NOR2X1_640/Y gnd AOI21X1_528/Y vdd AOI21X1
XAOI21X1_517 BUFX4_442/Y NOR2X1_60/Y NOR2X1_629/Y gnd AOI21X1_517/Y vdd AOI21X1
XAOI21X1_539 BUFX4_430/Y NOR2X1_97/B NOR2X1_651/Y gnd AOI21X1_539/Y vdd AOI21X1
XFILL_23_4_0 gnd vdd FILL
XFILL_24_9_1 gnd vdd FILL
XFILL_6_5_0 gnd vdd FILL
XBUFX4_107 BUFX4_14/Y gnd AND2X2_33/B vdd BUFX4
XBUFX4_118 BUFX4_75/A gnd BUFX4_118/Y vdd BUFX4
XBUFX4_129 INVX8_20/Y gnd BUFX4_129/Y vdd BUFX4
XFILL_14_4_0 gnd vdd FILL
XFILL_15_9_1 gnd vdd FILL
XOAI21X1_1019 BUFX4_351/Y INVX1_42/A BUFX4_154/Y gnd AOI21X1_437/C vdd OAI21X1
XOAI21X1_1008 INVX1_396/Y BUFX4_261/Y NAND2X1_305/Y gnd MUX2X1_244/B vdd OAI21X1
XDFFPOSX1_609 INVX1_16/A CLKBUF1_78/Y MUX2X1_11/Y gnd vdd DFFPOSX1
XOAI21X1_290 BUFX4_458/Y BUFX4_298/Y NOR2X1_459/A gnd OAI21X1_291/C vdd OAI21X1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XINVX1_321 INVX1_321/A gnd INVX1_321/Y vdd INVX1
XINVX1_332 INVX1_332/A gnd INVX1_332/Y vdd INVX1
XINVX1_343 INVX1_343/A gnd INVX1_343/Y vdd INVX1
XINVX1_376 INVX1_376/A gnd INVX1_376/Y vdd INVX1
XINVX1_387 INVX1_387/A gnd INVX1_387/Y vdd INVX1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XINVX1_365 INVX1_365/A gnd INVX1_365/Y vdd INVX1
XINVX1_398 INVX1_398/A gnd INVX1_398/Y vdd INVX1
XNOR2X1_701 NOR2X1_701/A INVX1_219/A gnd NOR2X1_701/Y vdd NOR2X1
XNOR2X1_734 NOR2X1_734/A MUX2X1_400/S gnd NOR2X1_734/Y vdd NOR2X1
XNOR2X1_723 NOR2X1_723/A NOR2X1_234/Y gnd NOR2X1_723/Y vdd NOR2X1
XNOR2X1_712 NOR2X1_712/A MUX2X1_120/S gnd NOR2X1_712/Y vdd NOR2X1
XAOI21X1_314 INVX1_86/Y BUFX4_339/Y OAI21X1_716/Y gnd OAI21X1_718/A vdd AOI21X1
XAOI21X1_303 BUFX4_77/Y AOI21X1_303/B NOR2X1_387/Y gnd OAI21X1_669/A vdd AOI21X1
XAOI21X1_325 BUFX4_410/Y OAI21X1_736/Y AOI21X1_325/C gnd OAI21X1_746/A vdd AOI21X1
XAOI21X1_358 INVX1_332/Y BUFX4_351/Y OAI21X1_821/Y gnd AOI21X1_358/Y vdd AOI21X1
XAOI21X1_336 BUFX4_412/Y MUX2X1_210/Y BUFX4_206/Y gnd AOI21X1_336/Y vdd AOI21X1
XAOI21X1_347 BUFX4_146/Y INVX1_326/Y OAI21X1_793/Y gnd OAI21X1_795/A vdd AOI21X1
XAOI21X1_369 INVX1_85/Y BUFX4_266/Y AOI21X1_369/C gnd AOI21X1_369/Y vdd AOI21X1
XDFFPOSX1_24 NOR2X1_268/A CLKBUF1_5/Y AOI21X1_172/Y gnd vdd DFFPOSX1
XOAI21X1_1531 BUFX4_451/Y BUFX4_312/Y INVX1_322/A gnd OAI21X1_1532/C vdd OAI21X1
XDFFPOSX1_35 OAI21X1_878/A CLKBUF1_25/Y OAI21X1_355/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 NOR2X1_601/A CLKBUF1_72/Y AOI21X1_165/Y gnd vdd DFFPOSX1
XOAI21X1_1520 NAND2X1_78/Y AND2X2_6/B OAI21X1_1520/C gnd DFFPOSX1_530/D vdd OAI21X1
XDFFPOSX1_46 INVX1_155/A CLKBUF1_98/Y MUX2X1_142/Y gnd vdd DFFPOSX1
XOAI21X1_1564 BUFX4_426/Y NAND2X1_85/Y OAI21X1_1563/Y gnd OAI21X1_1564/Y vdd OAI21X1
XOAI21X1_1542 BUFX4_67/Y NAND2X1_81/Y OAI21X1_1542/C gnd DFFPOSX1_557/D vdd OAI21X1
XDFFPOSX1_57 INVX1_162/A CLKBUF1_84/Y MUX2X1_149/Y gnd vdd DFFPOSX1
XOAI21X1_1553 BUFX4_124/Y BUFX4_196/Y OAI21X1_616/B gnd OAI21X1_1554/C vdd OAI21X1
XDFFPOSX1_68 INVX1_173/A CLKBUF1_66/Y MUX2X1_160/Y gnd vdd DFFPOSX1
XDFFPOSX1_79 NOR2X1_276/A CLKBUF1_80/Y AOI21X1_179/Y gnd vdd DFFPOSX1
XFILL_47_8_1 gnd vdd FILL
XFILL_46_3_0 gnd vdd FILL
XFILL_30_7_1 gnd vdd FILL
XDFFPOSX1_406 INVX1_236/A CLKBUF1_86/Y MUX2X1_342/Y gnd vdd DFFPOSX1
XDFFPOSX1_417 OAI21X1_1116/B CLKBUF1_8/Y OAI21X1_1421/Y gnd vdd DFFPOSX1
XDFFPOSX1_428 BUFX2_5/A CLKBUF1_96/Y OAI21X1_723/Y gnd vdd DFFPOSX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XDFFPOSX1_439 NOR2X1_629/A CLKBUF1_43/Y AOI21X1_517/Y gnd vdd DFFPOSX1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XINVX1_195 NOR3X1_4/Y gnd INVX1_195/Y vdd INVX1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XFILL_37_3_0 gnd vdd FILL
XFILL_38_8_1 gnd vdd FILL
XBUFX4_460 INVX8_10/Y gnd BUFX4_460/Y vdd BUFX4
XBUFX4_471 INVX8_15/Y gnd MUX2X1_58/A vdd BUFX4
XNOR2X1_531 BUFX4_337/Y INVX1_419/Y gnd NOR2X1_531/Y vdd NOR2X1
XNOR2X1_553 INVX1_11/A BUFX4_333/Y gnd OAI22X1_61/A vdd NOR2X1
XNOR2X1_542 BUFX4_290/Y NOR2X1_542/B gnd NOR2X1_542/Y vdd NOR2X1
XNOR2X1_520 NOR2X1_520/A NOR2X1_520/B gnd NOR2X1_520/Y vdd NOR2X1
XNOR2X1_575 NOR2X1_72/A BUFX4_352/Y gnd NOR2X1_575/Y vdd NOR2X1
XNOR2X1_564 NOR2X1_564/A BUFX4_153/Y gnd NOR2X1_564/Y vdd NOR2X1
XNOR2X1_586 NOR2X1_586/A BUFX4_335/Y gnd OAI22X1_73/A vdd NOR2X1
XNOR2X1_597 BUFX4_419/Y NOR2X1_597/B gnd OAI22X1_80/B vdd NOR2X1
XAOI21X1_100 BUFX4_174/Y NOR2X1_167/B NOR2X1_165/Y gnd AOI21X1_100/Y vdd AOI21X1
XAOI21X1_122 MUX2X1_97/B NOR2X1_703/B NOR2X1_197/Y gnd AOI21X1_122/Y vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XFILL_21_7_1 gnd vdd FILL
XAOI21X1_111 BUFX4_216/Y INVX1_219/A NOR2X1_181/Y gnd AOI21X1_111/Y vdd AOI21X1
XAOI21X1_133 MUX2X1_66/B MUX2X1_120/S NOR2X1_212/Y gnd AOI21X1_133/Y vdd AOI21X1
XAOI21X1_166 MUX2X1_39/B NOR2X1_261/B NOR2X1_261/Y gnd AOI21X1_166/Y vdd AOI21X1
XAOI21X1_155 BUFX4_469/Y NOR2X1_727/B NOR2X1_244/Y gnd AOI21X1_155/Y vdd AOI21X1
XAOI21X1_144 BUFX4_218/Y NOR2X1_231/B NOR2X1_228/Y gnd AOI21X1_144/Y vdd AOI21X1
XAOI21X1_177 BUFX4_473/Y MUX2X1_410/S NOR2X1_274/Y gnd DFFPOSX1_33/D vdd AOI21X1
XAOI21X1_188 BUFX4_468/Y NOR2X1_30/B NOR2X1_285/Y gnd DFFPOSX1_97/D vdd AOI21X1
XAOI21X1_199 MUX2X1_61/B NOR2X1_47/B NOR2X1_296/Y gnd AOI21X1_199/Y vdd AOI21X1
XOAI21X1_1350 BUFX4_386/Y BUFX4_187/Y OAI21X1_590/B gnd OAI21X1_1351/C vdd OAI21X1
XDFFPOSX1_940 INVX1_124/A CLKBUF1_9/Y MUX2X1_111/Y gnd vdd DFFPOSX1
XDFFPOSX1_951 NOR2X1_187/A CLKBUF1_61/Y AOI21X1_114/Y gnd vdd DFFPOSX1
XOAI21X1_1361 NAND2X1_53/Y BUFX4_424/Y OAI21X1_1361/C gnd DFFPOSX1_307/D vdd OAI21X1
XOAI21X1_1372 BUFX4_129/Y BUFX4_297/Y AOI21X1_476/B gnd OAI21X1_1372/Y vdd OAI21X1
XOAI21X1_1383 BUFX4_441/Y NAND2X1_58/Y OAI21X1_1383/C gnd DFFPOSX1_246/D vdd OAI21X1
XDFFPOSX1_962 NOR2X1_200/A CLKBUF1_37/Y AOI21X1_125/Y gnd vdd DFFPOSX1
XDFFPOSX1_984 NOR2X1_467/A CLKBUF1_95/Y AOI21X1_135/Y gnd vdd DFFPOSX1
XDFFPOSX1_973 INVX1_132/A CLKBUF1_46/Y MUX2X1_119/Y gnd vdd DFFPOSX1
XOAI21X1_1394 BUFX4_387/Y BUFX4_406/Y MUX2X1_230/B gnd OAI21X1_1395/C vdd OAI21X1
XDFFPOSX1_995 INVX1_135/A CLKBUF1_89/Y MUX2X1_122/Y gnd vdd DFFPOSX1
XFILL_4_8_1 gnd vdd FILL
XFILL_28_3_0 gnd vdd FILL
XFILL_29_8_1 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_203 NOR2X1_421/B CLKBUF1_8/Y AOI21X1_570/Y gnd vdd DFFPOSX1
XDFFPOSX1_214 NOR2X1_637/A CLKBUF1_86/Y AOI21X1_525/Y gnd vdd DFFPOSX1
XDFFPOSX1_236 INVX1_367/A CLKBUF1_50/Y MUX2X1_296/Y gnd vdd DFFPOSX1
XBUFX4_9 clock gnd BUFX4_9/Y vdd BUFX4
XDFFPOSX1_225 NOR2X1_528/A CLKBUF1_15/Y AOI21X1_537/Y gnd vdd DFFPOSX1
XDFFPOSX1_247 OAI21X1_766/B CLKBUF1_26/Y OAI21X1_1385/Y gnd vdd DFFPOSX1
XDFFPOSX1_258 INVX1_246/A CLKBUF1_69/Y MUX2X1_332/Y gnd vdd DFFPOSX1
XDFFPOSX1_269 NOR2X1_701/A CLKBUF1_8/Y AOI21X1_589/Y gnd vdd DFFPOSX1
XNAND2X1_306 INVX1_99/A BUFX4_262/Y gnd NAND2X1_306/Y vdd NAND2X1
XNAND2X1_317 INVX4_14/Y AOI22X1_31/Y gnd AOI22X1_33/A vdd NAND2X1
XNAND2X1_339 BUFX4_250/Y NOR2X1_726/A gnd NAND2X1_339/Y vdd NAND2X1
XNAND2X1_328 BUFX4_410/Y NAND2X1_328/B gnd AOI22X1_32/D vdd NAND2X1
XNOR3X1_13 INVX4_10/A NOR3X1_13/B NOR3X1_13/C gnd NOR3X1_13/Y vdd NOR3X1
XBUFX4_290 BUFX4_23/Y gnd BUFX4_290/Y vdd BUFX4
XNOR2X1_361 INVX1_3/A AND2X2_20/A gnd NOR2X1_361/Y vdd NOR2X1
XNOR2X1_350 INVX1_193/Y BUFX4_307/Y gnd INVX1_218/A vdd NOR2X1
XNOR2X1_372 BUFX4_356/Y INVX1_244/Y gnd NOR2X1_372/Y vdd NOR2X1
XNOR2X1_394 NOR2X1_394/A BUFX4_85/Y gnd NOR2X1_394/Y vdd NOR2X1
XNOR2X1_383 NOR2X1_383/A BUFX4_260/Y gnd NOR2X1_383/Y vdd NOR2X1
XINVX4_9 INVX4_9/A gnd INVX4_9/Y vdd INVX4
XOAI21X1_812 BUFX4_326/Y NOR2X1_18/A BUFX4_159/Y gnd OAI21X1_814/B vdd OAI21X1
XOAI21X1_823 BUFX4_352/Y NOR2X1_67/A BUFX4_157/Y gnd NOR2X1_445/B vdd OAI21X1
XOAI21X1_801 BUFX4_241/Y NAND2X1_362/A OAI21X1_801/C gnd OAI21X1_803/C vdd OAI21X1
XOAI21X1_867 BUFX4_347/Y NOR2X1_283/A BUFX4_146/Y gnd OAI22X1_27/C vdd OAI21X1
XOAI21X1_856 OAI21X1_856/A AND2X2_34/Y BUFX4_109/Y gnd OAI21X1_859/B vdd OAI21X1
XOAI21X1_834 INVX1_66/Y BUFX4_258/Y OAI21X1_834/C gnd MUX2X1_219/A vdd OAI21X1
XOAI21X1_845 BUFX4_335/Y NOR2X1_160/A BUFX4_152/Y gnd OAI22X1_26/C vdd OAI21X1
XOAI21X1_878 OAI21X1_878/A BUFX4_289/Y BUFX4_74/Y gnd OAI21X1_878/Y vdd OAI21X1
XOAI21X1_889 OAI21X1_889/A BUFX4_230/Y BUFX4_78/Y gnd OAI21X1_890/B vdd OAI21X1
XMUX2X1_301 INVX1_229/Y BUFX4_437/Y MUX2X1_66/S gnd MUX2X1_301/Y vdd MUX2X1
XMUX2X1_323 INVX1_373/Y BUFX4_67/Y MUX2X1_81/S gnd MUX2X1_323/Y vdd MUX2X1
XMUX2X1_312 INVX1_418/Y BUFX4_316/Y MUX2X1_71/S gnd MUX2X1_312/Y vdd MUX2X1
XMUX2X1_345 INVX1_420/Y BUFX4_317/Y MUX2X1_97/S gnd MUX2X1_345/Y vdd MUX2X1
XMUX2X1_334 BUFX4_441/Y INVX1_247/Y MUX2X1_92/S gnd MUX2X1_334/Y vdd MUX2X1
XOAI21X1_1180 NOR2X1_569/Y OAI21X1_1180/B OAI21X1_1178/Y gnd NOR2X1_570/B vdd OAI21X1
XOAI21X1_1191 NOR2X1_577/Y OAI21X1_1189/Y OAI21X1_1191/C gnd NOR2X1_578/B vdd OAI21X1
XMUX2X1_356 BUFX4_317/Y INVX1_421/Y MUX2X1_108/S gnd MUX2X1_356/Y vdd MUX2X1
XDFFPOSX1_770 NOR2X1_100/A CLKBUF1_4/Y AOI21X1_55/Y gnd vdd DFFPOSX1
XMUX2X1_389 BUFX4_440/Y INVX1_261/Y NOR2X1_727/B gnd MUX2X1_389/Y vdd MUX2X1
XDFFPOSX1_792 INVX1_85/A CLKBUF1_20/Y MUX2X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_781 INVX1_79/A CLKBUF1_99/Y MUX2X1_69/Y gnd vdd DFFPOSX1
XMUX2X1_378 BUFX4_445/Y INVX1_253/Y NOR2X1_220/B gnd MUX2X1_378/Y vdd MUX2X1
XMUX2X1_367 INVX1_382/Y BUFX4_68/Y MUX2X1_366/S gnd MUX2X1_367/Y vdd MUX2X1
XFILL_44_6_1 gnd vdd FILL
XFILL_43_1_0 gnd vdd FILL
XFILL_34_1_0 gnd vdd FILL
XFILL_35_6_1 gnd vdd FILL
XNOR2X1_90 BUFX4_55/Y BUFX4_383/Y gnd MUX2X1_55/S vdd NOR2X1
XOAI21X1_108 BUFX4_469/Y NAND2X1_37/Y OAI21X1_108/C gnd OAI21X1_108/Y vdd OAI21X1
XOAI21X1_119 BUFX4_449/Y BUFX4_53/Y INVX1_333/A gnd OAI21X1_119/Y vdd OAI21X1
XBUFX2_6 BUFX2_6/A gnd traffic_Street[1] vdd BUFX2
XNAND2X1_103 traffic_Street_1[0] BUFX4_174/Y gnd AOI22X1_2/C vdd NAND2X1
XNAND2X1_125 NAND3X1_27/Y OAI21X1_468/Y gnd NAND3X1_35/A vdd NAND2X1
XNAND2X1_114 INVX1_214/A NAND3X1_20/C gnd NAND3X1_19/B vdd NAND2X1
XNAND2X1_147 NAND2X1_147/A NOR3X1_7/Y gnd NAND2X1_148/B vdd NAND2X1
XNAND2X1_158 NAND2X1_158/A NOR3X1_7/Y gnd INVX1_211/A vdd NAND2X1
XNAND2X1_136 INVX1_200/A NOR3X1_7/Y gnd OAI21X1_497/A vdd NAND2X1
XNAND2X1_169 police_Interrupt INVX2_13/Y gnd NOR2X1_355/A vdd NAND2X1
XNAND2X1_1 NOR2X1_4/Y INVX2_6/A gnd NOR2X1_6/B vdd NAND2X1
XFILL_0_1_0 gnd vdd FILL
XFILL_1_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XNOR2X1_180 BUFX4_140/Y BUFX4_188/Y gnd INVX1_219/A vdd NOR2X1
XNOR2X1_191 BUFX4_434/Y BUFX4_449/Y gnd MUX2X1_364/S vdd NOR2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XOAI21X1_620 INVX1_18/Y BUFX4_333/Y BUFX4_146/Y gnd OAI21X1_620/Y vdd OAI21X1
XOAI21X1_642 INVX1_149/Y BUFX4_237/Y OAI21X1_642/C gnd MUX2X1_193/B vdd OAI21X1
XOAI21X1_631 BUFX4_339/Y OAI21X1_43/C BUFX4_158/Y gnd OAI22X1_6/C vdd OAI21X1
XAOI21X1_6 BUFX4_421/Y AOI21X1_7/B NOR2X1_24/Y gnd AOI21X1_6/Y vdd AOI21X1
XOAI21X1_664 OAI22X1_10/Y BUFX4_419/Y NAND3X1_73/Y gnd NOR2X1_385/B vdd OAI21X1
XOAI21X1_653 INVX1_180/A BUFX4_253/Y BUFX4_117/Y gnd OAI22X1_7/B vdd OAI21X1
XOAI21X1_675 OAI21X1_675/A OAI21X1_675/B BUFX4_37/Y gnd AND2X2_26/A vdd OAI21X1
XOAI21X1_686 OAI21X1_686/A BUFX4_284/Y BUFX4_87/Y gnd OAI22X1_14/B vdd OAI21X1
XOAI21X1_697 OAI22X1_15/Y BUFX4_413/Y AND2X2_48/B gnd OAI21X1_697/Y vdd OAI21X1
XMUX2X1_131 BUFX4_467/Y INVX1_144/Y NOR2X1_233/Y gnd MUX2X1_131/Y vdd MUX2X1
XMUX2X1_120 MUX2X1_59/B INVX1_133/Y MUX2X1_120/S gnd MUX2X1_120/Y vdd MUX2X1
XMUX2X1_164 INVX1_177/Y BUFX4_375/Y MUX2X1_21/S gnd MUX2X1_164/Y vdd MUX2X1
XMUX2X1_153 INVX1_166/Y BUFX4_470/Y MUX2X1_9/S gnd MUX2X1_153/Y vdd MUX2X1
XMUX2X1_142 INVX1_155/Y BUFX4_209/Y MUX2X1_2/S gnd MUX2X1_142/Y vdd MUX2X1
XFILL_9_7_1 gnd vdd FILL
XFILL_8_2_0 gnd vdd FILL
XMUX2X1_197 MUX2X1_197/A MUX2X1_197/B BUFX4_116/Y gnd MUX2X1_197/Y vdd MUX2X1
XMUX2X1_186 MUX2X1_185/Y MUX2X1_186/B INVX8_30/A gnd AOI22X1_15/D vdd MUX2X1
XMUX2X1_175 OR2X2_3/Y AND2X2_6/A traffic_Street_0[3] gnd AND2X2_5/A vdd MUX2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XDFFPOSX1_1 DFFPOSX1_1/Q CLKBUF1_57/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_16_1_0 gnd vdd FILL
XFILL_17_6_1 gnd vdd FILL
XNOR2X1_4 INVX1_2/Y INVX2_2/Y gnd NOR2X1_4/Y vdd NOR2X1
XFILL_50_4_1 gnd vdd FILL
XAOI21X1_14 MUX2X1_8/B NOR2X1_33/Y NOR2X1_36/Y gnd AOI21X1_14/Y vdd AOI21X1
XAOI21X1_25 BUFX4_473/Y NOR2X1_54/Y NOR2X1_56/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_47 MUX2X1_82/B MUX2X1_50/S NOR2X1_88/Y gnd AOI21X1_47/Y vdd AOI21X1
XAOI21X1_36 BUFX4_213/Y NOR2X1_70/Y NOR2X1_71/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_58 MUX2X1_58/A MUX2X1_75/S AOI21X1_58/C gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_69 BUFX4_176/Y MUX2X1_320/S NOR2X1_122/Y gnd AOI21X1_69/Y vdd AOI21X1
XOAI21X1_9 MUX2X1_4/B OAI21X1_7/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_33 OAI22X1_33/A OAI22X1_33/B OAI22X1_33/C OAI22X1_33/D gnd OAI22X1_33/Y vdd
+ OAI22X1
XOAI22X1_11 NOR2X1_389/Y OAI22X1_11/B OAI22X1_11/C NOR2X1_388/Y gnd OAI22X1_11/Y vdd
+ OAI22X1
XFILL_41_4_1 gnd vdd FILL
XOAI22X1_22 NOR2X1_429/Y OAI22X1_22/B OAI22X1_22/C OAI22X1_22/D gnd NOR2X1_430/B vdd
+ OAI22X1
XOAI22X1_44 OAI22X1_44/A OAI22X1_44/B MUX2X1_241/Y BUFX4_39/Y gnd OAI22X1_44/Y vdd
+ OAI22X1
XOAI22X1_66 OAI22X1_66/A OAI22X1_66/B NOR2X1_568/Y OAI22X1_66/D gnd OAI22X1_66/Y vdd
+ OAI22X1
XOAI22X1_55 NOR2X1_535/Y OAI22X1_55/B OAI22X1_55/C BUFX4_168/Y gnd NOR2X1_538/B vdd
+ OAI22X1
XOAI22X1_77 OAI22X1_77/A OAI22X1_77/B OAI22X1_77/C NOR2X1_593/Y gnd OAI22X1_77/Y vdd
+ OAI22X1
XOAI22X1_88 NOR2X1_616/Y OAI22X1_88/B OAI22X1_88/C NOR2X1_615/Y gnd OAI22X1_88/Y vdd
+ OAI22X1
XOAI21X1_450 NOR2X1_304/Y AND2X2_4/Y INVX2_15/Y gnd AOI22X1_3/C vdd OAI21X1
XOAI21X1_461 AOI21X1_212/B INVX2_17/Y MUX2X1_176/B gnd OAI21X1_461/Y vdd OAI21X1
XOAI21X1_483 AOI21X1_224/Y NAND3X1_39/Y AOI21X1_225/Y gnd OAI21X1_483/Y vdd OAI21X1
XOAI21X1_472 AND2X2_6/B NOR2X1_308/B MUX2X1_174/B gnd OAI21X1_472/Y vdd OAI21X1
XOAI21X1_494 AND2X2_3/B NOR2X1_300/B NAND3X1_7/C gnd INVX1_209/A vdd OAI21X1
XFILL_49_5_1 gnd vdd FILL
XFILL_48_0_0 gnd vdd FILL
XFILL_32_4_1 gnd vdd FILL
XAOI21X1_507 BUFX4_204/Y AOI21X1_507/B AOI21X1_503/Y gnd AND2X2_54/A vdd AOI21X1
XAOI21X1_518 BUFX4_421/Y NOR2X1_60/Y NOR2X1_630/Y gnd AOI21X1_518/Y vdd AOI21X1
XAOI21X1_529 BUFX4_430/Y NOR2X1_83/B NOR2X1_641/Y gnd AOI21X1_529/Y vdd AOI21X1
XFILL_39_0_0 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XBUFX4_108 BUFX4_82/A gnd BUFX4_108/Y vdd BUFX4
XBUFX4_119 BUFX4_124/A gnd BUFX4_119/Y vdd BUFX4
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_1009 INVX1_95/Y BUFX4_263/Y NAND2X1_306/Y gnd MUX2X1_244/A vdd OAI21X1
XINVX1_300 INVX1_300/A gnd INVX1_300/Y vdd INVX1
XOAI21X1_291 NAND2X1_75/Y BUFX4_176/Y OAI21X1_291/C gnd OAI21X1_291/Y vdd OAI21X1
XOAI21X1_280 BUFX4_192/Y BUFX4_163/Y AND2X2_25/A gnd OAI21X1_281/C vdd OAI21X1
XINVX1_322 INVX1_322/A gnd INVX1_322/Y vdd INVX1
XINVX1_344 INVX1_344/A gnd INVX1_344/Y vdd INVX1
XINVX1_333 INVX1_333/A gnd INVX1_333/Y vdd INVX1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XINVX1_377 INVX1_377/A gnd INVX1_377/Y vdd INVX1
XINVX1_366 INVX1_366/A gnd INVX1_366/Y vdd INVX1
XINVX1_355 INVX1_355/A gnd INVX1_355/Y vdd INVX1
XINVX1_388 INVX1_388/A gnd INVX1_388/Y vdd INVX1
XINVX1_399 INVX1_399/A gnd INVX1_399/Y vdd INVX1
XNOR2X1_702 NOR2X1_702/A NOR2X1_188/B gnd NOR2X1_702/Y vdd NOR2X1
XNOR2X1_713 NOR2X1_713/A MUX2X1_376/S gnd NOR2X1_713/Y vdd NOR2X1
XNOR2X1_724 NOR2X1_724/A NOR2X1_234/Y gnd NOR2X1_724/Y vdd NOR2X1
XNOR2X1_735 NOR2X1_735/A NOR2X1_261/B gnd NOR2X1_735/Y vdd NOR2X1
XFILL_29_1 gnd vdd FILL
XAOI21X1_304 AOI21X1_304/A AND2X2_29/A BUFX4_79/Y gnd OAI21X1_670/C vdd AOI21X1
XAOI21X1_315 INVX1_290/Y BUFX4_242/Y OAI21X1_717/Y gnd OAI21X1_718/B vdd AOI21X1
XAOI21X1_326 BUFX4_109/Y INVX1_303/Y BUFX4_334/Y gnd AOI21X1_326/Y vdd AOI21X1
XAOI21X1_337 BUFX4_329/Y INVX1_314/Y BUFX4_150/Y gnd AOI21X1_337/Y vdd AOI21X1
XAOI21X1_348 BUFX4_146/Y INVX1_327/Y AOI21X1_348/C gnd OAI21X1_795/B vdd AOI21X1
XAOI21X1_359 BUFX4_90/Y AOI21X1_359/B AOI21X1_358/Y gnd AOI21X1_359/Y vdd AOI21X1
XDFFPOSX1_36 INVX1_404/A CLKBUF1_25/Y OAI21X1_357/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 NOR2X1_269/A CLKBUF1_72/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XOAI21X1_1532 NAND2X1_80/Y BUFX4_428/Y OAI21X1_1532/C gnd DFFPOSX1_544/D vdd OAI21X1
XDFFPOSX1_14 NOR2X1_261/A CLKBUF1_78/Y AOI21X1_166/Y gnd vdd DFFPOSX1
XOAI21X1_1510 BUFX4_63/Y NAND2X1_77/Y OAI21X1_1510/C gnd OAI21X1_1510/Y vdd OAI21X1
XOAI21X1_1521 BUFX4_386/Y BUFX4_311/Y MUX2X1_182/A gnd OAI21X1_1522/C vdd OAI21X1
XOAI21X1_1554 NAND2X1_84/Y BUFX4_442/Y OAI21X1_1554/C gnd DFFPOSX1_583/D vdd OAI21X1
XDFFPOSX1_69 INVX1_174/A CLKBUF1_72/Y MUX2X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 INVX1_156/A CLKBUF1_81/Y MUX2X1_143/Y gnd vdd DFFPOSX1
XOAI21X1_1543 BUFX4_189/Y BUFX4_312/Y AND2X2_53/B gnd OAI21X1_1544/C vdd OAI21X1
XOAI21X1_1565 BUFX4_188/Y BUFX4_197/Y NOR2X1_486/A gnd OAI21X1_1566/C vdd OAI21X1
XDFFPOSX1_58 INVX1_163/A CLKBUF1_47/Y MUX2X1_150/Y gnd vdd DFFPOSX1
XFILL_46_3_1 gnd vdd FILL
XDFFPOSX1_429 BUFX2_6/A CLKBUF1_96/Y OAI21X1_910/Y gnd vdd DFFPOSX1
XDFFPOSX1_407 INVX1_307/A CLKBUF1_22/Y MUX2X1_343/Y gnd vdd DFFPOSX1
XDFFPOSX1_418 INVX1_193/A CLKBUF1_71/Y NAND2X1_167/Y gnd vdd DFFPOSX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_141 INVX1_141/A gnd INVX1_141/Y vdd INVX1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XCLKBUF1_100 BUFX4_3/Y gnd CLKBUF1_100/Y vdd CLKBUF1
XFILL_37_3_1 gnd vdd FILL
XBUFX4_450 BUFX4_449/A gnd BUFX4_450/Y vdd BUFX4
XBUFX4_472 INVX8_15/Y gnd MUX2X1_83/B vdd BUFX4
XNOR2X1_510 NOR2X1_509/Y NOR2X1_510/B gnd NOR2X1_510/Y vdd NOR2X1
XBUFX4_461 INVX8_10/Y gnd BUFX4_461/Y vdd BUFX4
XNOR2X1_521 NOR2X1_521/A BUFX4_351/Y gnd NOR2X1_521/Y vdd NOR2X1
XNOR2X1_543 INVX1_458/A BUFX4_325/Y gnd OAI22X1_57/A vdd NOR2X1
XNOR2X1_532 NOR2X1_701/A BUFX4_335/Y gnd NOR2X1_532/Y vdd NOR2X1
XNOR2X1_554 BUFX4_419/Y NOR2X1_554/B gnd OAI22X1_63/A vdd NOR2X1
XNOR2X1_576 BUFX4_50/Y OAI22X1_69/Y gnd NOR2X1_576/Y vdd NOR2X1
XNOR2X1_565 BUFX4_76/Y NOR2X1_565/B gnd NOR2X1_565/Y vdd NOR2X1
XNOR2X1_598 NOR2X1_598/A BUFX4_223/Y gnd NOR2X1_598/Y vdd NOR2X1
XNOR2X1_587 BUFX4_417/Y OAI22X1_73/Y gnd NOR2X1_587/Y vdd NOR2X1
XAOI21X1_123 BUFX4_177/Y NOR2X1_703/B NOR2X1_198/Y gnd AOI21X1_123/Y vdd AOI21X1
XAOI21X1_101 MUX2X1_57/A NOR2X1_167/B NOR2X1_166/Y gnd AOI21X1_101/Y vdd AOI21X1
XAOI21X1_112 MUX2X1_44/A INVX1_219/A NOR2X1_182/Y gnd AOI21X1_112/Y vdd AOI21X1
XAOI21X1_167 MUX2X1_40/B NOR2X1_261/B NOR2X1_262/Y gnd DFFPOSX1_15/D vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_156 BUFX4_218/Y NOR2X1_729/B NOR2X1_246/Y gnd AOI21X1_156/Y vdd AOI21X1
XAOI21X1_145 BUFX4_176/Y NOR2X1_231/B NOR2X1_229/Y gnd AOI21X1_145/Y vdd AOI21X1
XAOI21X1_134 MUX2X1_97/B MUX2X1_376/S NOR2X1_214/Y gnd AOI21X1_134/Y vdd AOI21X1
XAOI21X1_178 BUFX4_213/Y NOR2X1_16/Y NOR2X1_275/Y gnd AOI21X1_178/Y vdd AOI21X1
XAOI21X1_189 BUFX4_213/Y NOR2X1_33/Y NOR2X1_286/Y gnd AOI21X1_189/Y vdd AOI21X1
XOAI21X1_1340 INVX1_248/Y NAND2X1_50/B NAND2X1_356/Y gnd OAI21X1_1340/Y vdd OAI21X1
XDFFPOSX1_930 INVX1_121/A CLKBUF1_27/Y MUX2X1_108/Y gnd vdd DFFPOSX1
XDFFPOSX1_941 INVX1_125/A CLKBUF1_49/Y MUX2X1_112/Y gnd vdd DFFPOSX1
XOAI21X1_1362 BUFX4_454/Y BUFX4_185/Y INVX1_372/A gnd OAI21X1_1363/C vdd OAI21X1
XOAI21X1_1373 NAND2X1_56/Y BUFX4_321/Y OAI21X1_1372/Y gnd OAI21X1_1373/Y vdd OAI21X1
XOAI21X1_1351 NAND2X1_52/Y BUFX4_440/Y OAI21X1_1351/C gnd DFFPOSX1_318/D vdd OAI21X1
XDFFPOSX1_963 NAND2X1_210/A CLKBUF1_9/Y OAI21X1_257/Y gnd vdd DFFPOSX1
XDFFPOSX1_952 NOR2X1_188/A CLKBUF1_61/Y AOI21X1_115/Y gnd vdd DFFPOSX1
XOAI21X1_1384 BUFX4_136/Y BUFX4_127/Y OAI21X1_766/B gnd OAI21X1_1384/Y vdd OAI21X1
XDFFPOSX1_985 NOR2X1_216/A CLKBUF1_15/Y AOI21X1_136/Y gnd vdd DFFPOSX1
XOAI21X1_1395 NAND2X1_59/Y BUFX4_73/Y OAI21X1_1395/C gnd DFFPOSX1_196/D vdd OAI21X1
XDFFPOSX1_974 NOR2X1_204/A CLKBUF1_1/Y AOI21X1_127/Y gnd vdd DFFPOSX1
XDFFPOSX1_996 NOR2X1_219/A CLKBUF1_68/Y AOI21X1_138/Y gnd vdd DFFPOSX1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFPOSX1_204 INVX1_369/A CLKBUF1_86/Y MUX2X1_338/Y gnd vdd DFFPOSX1
XDFFPOSX1_226 INVX1_247/A CLKBUF1_69/Y MUX2X1_334/Y gnd vdd DFFPOSX1
XDFFPOSX1_215 INVX1_301/A CLKBUF1_44/Y DFFPOSX1_215/D gnd vdd DFFPOSX1
XDFFPOSX1_237 NOR2X1_645/A CLKBUF1_15/Y AOI21X1_533/Y gnd vdd DFFPOSX1
XDFFPOSX1_259 NOR2X1_427/B CLKBUF1_26/Y AOI21X1_563/Y gnd vdd DFFPOSX1
XDFFPOSX1_248 OAI21X1_924/B CLKBUF1_26/Y OAI21X1_1387/Y gnd vdd DFFPOSX1
XNAND2X1_318 NOR2X1_280/A AND2X2_36/B gnd NAND2X1_318/Y vdd NAND2X1
XNAND2X1_307 OAI21X1_220/C BUFX4_418/Y gnd NAND2X1_307/Y vdd NAND2X1
XNAND2X1_329 NAND2X1_329/A BUFX4_249/Y gnd NAND2X1_329/Y vdd NAND2X1
XNOR3X1_14 BUFX4_36/Y NOR3X1_14/B NOR3X1_14/C gnd NOR3X1_14/Y vdd NOR3X1
XBUFX4_291 BUFX4_18/Y gnd BUFX4_291/Y vdd BUFX4
XBUFX4_280 BUFX4_19/Y gnd BUFX4_280/Y vdd BUFX4
XNOR2X1_340 INVX2_21/A XNOR2X1_4/A gnd NOR2X1_341/A vdd NOR2X1
XNOR2X1_351 traffic_Street_0[3] NOR2X1_351/B gnd OAI22X1_3/A vdd NOR2X1
XNOR2X1_373 BUFX4_362/Y INVX1_255/Y gnd NOR2X1_373/Y vdd NOR2X1
XNOR2X1_395 NOR2X1_393/Y NOR2X1_395/B gnd NOR2X1_395/Y vdd NOR2X1
XNOR2X1_362 NOR2X1_361/Y AND2X2_20/Y gnd NOR2X1_362/Y vdd NOR2X1
XNOR2X1_384 NOR2X1_384/A BUFX4_331/Y gnd OAI22X1_10/A vdd NOR2X1
XOAI21X1_824 OAI21X1_85/C BUFX4_251/Y BUFX4_91/Y gnd OAI21X1_824/Y vdd OAI21X1
XOAI21X1_813 NOR2X1_24/A BUFX4_326/Y AOI21X1_355/Y gnd OAI21X1_813/Y vdd OAI21X1
XOAI21X1_802 NAND2X1_6/A BUFX4_242/Y BUFX4_88/Y gnd OAI21X1_803/B vdd OAI21X1
XOAI21X1_857 INVX1_336/Y INVX8_30/A AOI21X1_377/Y gnd NAND3X1_74/C vdd OAI21X1
XOAI21X1_835 INVX1_333/Y BUFX4_260/Y OAI21X1_835/C gnd OAI21X1_835/Y vdd OAI21X1
XOAI21X1_846 OAI21X1_846/A BUFX4_272/Y BUFX4_104/Y gnd OAI22X1_26/B vdd OAI21X1
XOAI21X1_879 OAI21X1_879/A AOI21X1_385/Y BUFX4_416/Y gnd OAI21X1_879/Y vdd OAI21X1
XOAI21X1_868 OAI21X1_868/A BUFX4_281/Y BUFX4_115/Y gnd OAI22X1_27/B vdd OAI21X1
XMUX2X1_313 MUX2X1_9/B INVX1_231/Y MUX2X1_75/S gnd MUX2X1_313/Y vdd MUX2X1
XMUX2X1_302 INVX1_293/Y BUFX4_430/Y MUX2X1_66/S gnd MUX2X1_302/Y vdd MUX2X1
XMUX2X1_346 BUFX4_437/Y INVX1_235/Y NOR2X1_172/B gnd MUX2X1_346/Y vdd MUX2X1
XMUX2X1_357 INVX1_257/Y BUFX4_444/Y MUX2X1_360/S gnd MUX2X1_357/Y vdd MUX2X1
XOAI21X1_1181 BUFX4_361/Y NOR2X1_56/A BUFX4_154/Y gnd OAI22X1_67/C vdd OAI21X1
XMUX2X1_335 BUFX4_426/Y INVX1_314/Y MUX2X1_92/S gnd MUX2X1_335/Y vdd MUX2X1
XMUX2X1_324 INVX1_454/Y BUFX4_322/Y MUX2X1_81/S gnd MUX2X1_324/Y vdd MUX2X1
XOAI21X1_1170 AND2X2_27/A INVX1_438/Y AOI21X1_491/Y gnd OAI21X1_1170/Y vdd OAI21X1
XOAI21X1_1192 INVX1_64/Y BUFX4_272/Y NAND2X1_343/Y gnd MUX2X1_261/B vdd OAI21X1
XDFFPOSX1_771 INVX1_69/A CLKBUF1_95/Y MUX2X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_760 NOR2X1_93/A CLKBUF1_68/Y AOI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_793 NOR2X1_104/A CLKBUF1_55/Y AOI21X1_57/Y gnd vdd DFFPOSX1
XMUX2X1_379 BUFX4_66/Y INVX1_375/Y NOR2X1_220/B gnd MUX2X1_379/Y vdd MUX2X1
XDFFPOSX1_782 INVX1_80/A CLKBUF1_63/Y MUX2X1_70/Y gnd vdd DFFPOSX1
XMUX2X1_368 INVX1_430/Y MUX2X1_29/B MUX2X1_366/S gnd MUX2X1_368/Y vdd MUX2X1
XFILL_43_1_1 gnd vdd FILL
XNAND3X1_80 BUFX4_32/Y NAND3X1_80/B NAND3X1_80/C gnd NAND3X1_80/Y vdd NAND3X1
XNOR2X1_80 NOR2X1_80/A NOR2X1_83/B gnd NOR2X1_80/Y vdd NOR2X1
XFILL_34_1_1 gnd vdd FILL
XNOR2X1_91 BUFX4_55/Y NOR2X1_39/B gnd NOR2X1_92/B vdd NOR2X1
XFILL_11_1 gnd vdd FILL
XOAI21X1_109 BUFX4_61/Y BUFX4_54/Y NAND2X1_224/A gnd OAI21X1_110/C vdd OAI21X1
XBUFX2_7 BUFX2_7/A gnd traffic_Street[2] vdd BUFX2
XNAND2X1_104 traffic_Street_1[1] AND2X2_2/B gnd AOI22X1_2/D vdd NAND2X1
XNAND2X1_115 BUFX4_73/Y NAND3X1_14/B gnd NAND3X1_22/C vdd NAND2X1
XNAND2X1_126 OAI21X1_471/Y NAND3X1_30/Y gnd NAND3X1_37/A vdd NAND2X1
XNAND2X1_148 ped_Vert_Interrupt NAND2X1_148/B gnd INVX1_208/A vdd NAND2X1
XNAND2X1_159 NAND2X1_148/B AND2X2_14/B gnd NAND2X1_159/Y vdd NAND2X1
XNAND2X1_137 NAND2X1_137/A XNOR2X1_1/A gnd INVX1_203/A vdd NAND2X1
XNAND2X1_2 NOR2X1_2/Y NOR2X1_6/Y gnd NAND2X1_2/Y vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_170 NOR2X1_170/A NOR2X1_172/B gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_192 NOR2X1_192/A MUX2X1_364/S gnd NOR2X1_192/Y vdd NOR2X1
XNOR2X1_181 NOR2X1_181/A INVX1_219/A gnd NOR2X1_181/Y vdd NOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XOAI21X1_621 OAI21X1_620/Y NOR2X1_374/Y BUFX4_411/Y gnd OAI21X1_624/B vdd OAI21X1
XOAI21X1_610 INVX1_265/Y BUFX4_280/Y OAI21X1_610/C gnd MUX2X1_184/A vdd OAI21X1
XOAI21X1_632 INVX1_34/A BUFX4_230/Y BUFX4_111/Y gnd OAI22X1_6/B vdd OAI21X1
XOAI21X1_665 BUFX4_337/Y NOR2X1_197/A BUFX4_151/Y gnd NOR2X1_387/B vdd OAI21X1
XAOI21X1_7 BUFX4_64/Y AOI21X1_7/B NOR2X1_25/Y gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_643 INVX1_277/Y AND2X2_22/A OAI21X1_643/C gnd MUX2X1_193/A vdd OAI21X1
XOAI21X1_654 OAI22X1_7/Y BUFX4_416/Y BUFX4_206/Y gnd AOI21X1_298/C vdd OAI21X1
XOAI21X1_687 OAI22X1_14/Y BUFX4_411/Y BUFX4_202/Y gnd OAI21X1_687/Y vdd OAI21X1
XOAI21X1_698 BUFX4_394/Y OAI21X1_698/B OAI21X1_688/Y gnd MUX2X1_207/B vdd OAI21X1
XOAI21X1_676 AND2X2_26/Y BUFX4_170/Y BUFX4_391/Y gnd OAI22X1_12/B vdd OAI21X1
XMUX2X1_110 INVX1_123/Y MUX2X1_97/B MUX2X1_360/S gnd MUX2X1_110/Y vdd MUX2X1
XMUX2X1_132 BUFX4_217/Y INVX1_145/Y MUX2X1_397/S gnd DFFPOSX1_2/D vdd MUX2X1
XMUX2X1_121 BUFX4_371/Y INVX1_134/Y MUX2X1_120/S gnd MUX2X1_121/Y vdd MUX2X1
XMUX2X1_165 INVX1_178/Y BUFX4_470/Y MUX2X1_21/S gnd MUX2X1_165/Y vdd MUX2X1
XMUX2X1_143 INVX1_156/Y BUFX4_178/Y MUX2X1_2/S gnd MUX2X1_143/Y vdd MUX2X1
XMUX2X1_154 INVX1_167/Y BUFX4_209/Y MUX2X1_14/S gnd MUX2X1_154/Y vdd MUX2X1
XMUX2X1_176 MUX2X1_176/A MUX2X1_176/B AND2X2_15/B gnd MUX2X1_176/Y vdd MUX2X1
XDFFPOSX1_590 NOR2X1_551/A CLKBUF1_72/Y DFFPOSX1_590/D gnd vdd DFFPOSX1
XMUX2X1_198 MUX2X1_198/A MUX2X1_198/B BUFX4_118/Y gnd MUX2X1_198/Y vdd MUX2X1
XMUX2X1_187 MUX2X1_187/A MUX2X1_187/B BUFX4_108/Y gnd MUX2X1_187/Y vdd MUX2X1
XFILL_8_2_1 gnd vdd FILL
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XFILL_45_9_0 gnd vdd FILL
XDFFPOSX1_2 INVX1_145/A CLKBUF1_52/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 INVX1_3/Y INVX2_3/Y gnd INVX2_6/A vdd NOR2X1
XFILL_36_9_0 gnd vdd FILL
XAOI21X1_15 BUFX4_443/Y NOR2X1_43/B NOR2X1_40/Y gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 BUFX4_214/Y NOR2X1_57/Y NOR2X1_58/Y gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_37 BUFX4_468/Y NOR2X1_70/Y NOR2X1_72/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_59 MUX2X1_71/B NOR2X1_107/B AOI21X1_59/C gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_48 MUX2X1_59/B NOR2X1_92/B NOR2X1_92/Y gnd AOI21X1_48/Y vdd AOI21X1
XFILL_2_9_0 gnd vdd FILL
XFILL_27_9_0 gnd vdd FILL
XOAI22X1_23 OAI22X1_23/A OAI22X1_23/B OAI22X1_23/C OAI22X1_23/D gnd OAI22X1_23/Y vdd
+ OAI22X1
XOAI22X1_12 OAI22X1_12/A OAI22X1_12/B OAI22X1_12/C BUFX4_391/Y gnd MUX2X1_199/A vdd
+ OAI22X1
XOAI22X1_34 OAI22X1_34/A OAI22X1_34/B OAI22X1_34/C OAI22X1_34/D gnd NOR2X1_468/B vdd
+ OAI22X1
XOAI22X1_45 NOR2X1_506/Y OAI22X1_45/B OAI22X1_45/C NOR2X1_505/Y gnd OAI22X1_45/Y vdd
+ OAI22X1
XOAI22X1_67 OAI22X1_67/A OAI22X1_67/B OAI22X1_67/C NOR2X1_571/Y gnd OAI22X1_67/Y vdd
+ OAI22X1
XOAI22X1_56 NOR2X1_540/Y OAI22X1_56/B OAI22X1_56/C NOR2X1_539/Y gnd NOR2X1_541/B vdd
+ OAI22X1
XOAI22X1_78 NOR2X1_596/Y OAI22X1_78/B OAI22X1_78/C NOR2X1_595/Y gnd NOR2X1_597/B vdd
+ OAI22X1
XOAI22X1_89 OAI22X1_89/A OAI22X1_89/B OAI22X1_89/C OAI22X1_89/D gnd MUX2X1_264/B vdd
+ OAI22X1
XOAI21X1_440 AOI22X1_1/Y INVX1_187/A INVX4_6/A gnd NAND2X1_105/B vdd OAI21X1
XFILL_10_8_0 gnd vdd FILL
XOAI21X1_462 INVX2_16/Y AND2X2_2/A OAI21X1_462/C gnd AOI21X1_213/C vdd OAI21X1
XOAI21X1_484 NOR2X1_321/B INVX4_8/Y INVX1_188/Y gnd NAND2X1_137/A vdd OAI21X1
XOAI21X1_473 INVX1_189/A OAI21X1_473/B OAI21X1_472/Y gnd NAND3X1_32/B vdd OAI21X1
XOAI21X1_451 AOI22X1_3/Y INVX1_190/A INVX4_6/A gnd OAI21X1_451/Y vdd OAI21X1
XOAI21X1_495 NAND3X1_28/C OAI22X1_2/A AOI22X1_6/A gnd NAND2X1_141/A vdd OAI21X1
XFILL_48_0_1 gnd vdd FILL
XFILL_18_9_0 gnd vdd FILL
XAOI21X1_508 INVX1_183/Y BUFX4_368/Y BUFX4_156/Y gnd AOI21X1_508/Y vdd AOI21X1
XAOI21X1_519 BUFX4_321/Y NOR2X1_60/Y NOR2X1_631/Y gnd AOI21X1_519/Y vdd AOI21X1
XFILL_39_0_1 gnd vdd FILL
XBUFX4_109 BUFX4_85/A gnd BUFX4_109/Y vdd BUFX4
XFILL_5_0_1 gnd vdd FILL
XFILL_42_7_0 gnd vdd FILL
XOAI21X1_292 BUFX4_456/Y BUFX4_298/Y NOR2X1_518/A gnd OAI21X1_293/C vdd OAI21X1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XOAI21X1_281 BUFX4_216/Y NAND2X1_74/Y OAI21X1_281/C gnd OAI21X1_281/Y vdd OAI21X1
XOAI21X1_270 BUFX4_452/Y BUFX4_164/Y NOR2X1_615/A gnd OAI21X1_270/Y vdd OAI21X1
XINVX1_312 INVX1_312/A gnd INVX1_312/Y vdd INVX1
XINVX1_323 INVX1_323/A gnd INVX1_323/Y vdd INVX1
XINVX1_334 INVX1_334/A gnd INVX1_334/Y vdd INVX1
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XINVX1_367 INVX1_367/A gnd INVX1_367/Y vdd INVX1
XINVX1_345 INVX1_345/A gnd INVX1_345/Y vdd INVX1
XINVX1_356 INVX1_356/A gnd INVX1_356/Y vdd INVX1
XINVX1_389 INVX1_389/A gnd INVX1_389/Y vdd INVX1
XNOR2X1_703 NOR2X1_703/A NOR2X1_703/B gnd NOR2X1_703/Y vdd NOR2X1
XNOR2X1_725 NOR2X1_725/A NOR2X1_234/Y gnd NOR2X1_725/Y vdd NOR2X1
XNOR2X1_714 NOR2X1_714/A NOR2X1_220/B gnd NOR2X1_714/Y vdd NOR2X1
XNOR2X1_736 NOR2X1_736/A NOR2X1_737/B gnd NOR2X1_736/Y vdd NOR2X1
XFILL_33_7_0 gnd vdd FILL
XAOI21X1_316 AOI21X1_316/A AOI21X1_316/B BUFX4_166/Y gnd NOR2X1_411/A vdd AOI21X1
XAOI21X1_305 NOR2X1_206/A BUFX4_272/Y AOI21X1_305/C gnd OAI21X1_675/A vdd AOI21X1
XAOI21X1_349 BUFX4_154/Y INVX1_328/Y AOI21X1_349/C gnd AOI21X1_349/Y vdd AOI21X1
XAOI21X1_327 BUFX4_157/Y INVX1_304/Y OAI21X1_742/Y gnd AOI21X1_327/Y vdd AOI21X1
XAOI21X1_338 BUFX4_51/Y AOI22X1_20/Y OAI21X1_771/Y gnd AOI21X1_339/C vdd AOI21X1
XOAI21X1_1511 BUFX4_137/Y BUFX4_455/Y NAND2X1_338/B gnd OAI21X1_1511/Y vdd OAI21X1
XDFFPOSX1_15 NOR2X1_262/A CLKBUF1_25/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX1_151/A CLKBUF1_11/Y MUX2X1_138/Y gnd vdd DFFPOSX1
XOAI21X1_1522 NAND2X1_79/Y BUFX4_440/Y OAI21X1_1522/C gnd DFFPOSX1_535/D vdd OAI21X1
XOAI21X1_1500 NAND2X1_76/Y BUFX4_429/Y OAI21X1_1500/C gnd DFFPOSX1_504/D vdd OAI21X1
XOAI21X1_1533 NOR2X1_84/B BUFX4_309/Y INVX1_387/A gnd OAI21X1_1534/C vdd OAI21X1
XOAI21X1_1555 BUFX4_124/Y BUFX4_196/Y OAI21X1_796/B gnd OAI21X1_1556/C vdd OAI21X1
XOAI21X1_1544 BUFX4_322/Y NAND2X1_81/Y OAI21X1_1544/C gnd DFFPOSX1_558/D vdd OAI21X1
XDFFPOSX1_37 DFFPOSX1_37/Q CLKBUF1_11/Y OAI21X1_359/Y gnd vdd DFFPOSX1
XOAI21X1_1566 BUFX4_63/Y NAND2X1_85/Y OAI21X1_1566/C gnd DFFPOSX1_589/D vdd OAI21X1
XDFFPOSX1_59 INVX1_164/A CLKBUF1_81/Y MUX2X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 INVX1_157/A CLKBUF1_98/Y MUX2X1_144/Y gnd vdd DFFPOSX1
XFILL_24_7_0 gnd vdd FILL
XFILL_7_8_0 gnd vdd FILL
XCLKBUF1_90 BUFX4_5/Y gnd CLKBUF1_90/Y vdd CLKBUF1
XFILL_15_7_0 gnd vdd FILL
XDFFPOSX1_408 INVX1_357/A CLKBUF1_83/Y MUX2X1_344/Y gnd vdd DFFPOSX1
XDFFPOSX1_419 NAND2X1_168/A CLKBUF1_71/Y XOR2X1_4/Y gnd vdd DFFPOSX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XCLKBUF1_101 BUFX4_8/Y gnd CLKBUF1_101/Y vdd CLKBUF1
XBUFX4_440 INVX8_2/Y gnd BUFX4_440/Y vdd BUFX4
XNOR2X1_500 NOR2X1_500/A NOR2X1_500/B gnd NOR2X1_500/Y vdd NOR2X1
XBUFX4_473 INVX8_15/Y gnd BUFX4_473/Y vdd BUFX4
XBUFX4_462 INVX8_10/Y gnd BUFX4_462/Y vdd BUFX4
XBUFX4_451 BUFX4_449/A gnd BUFX4_451/Y vdd BUFX4
XFILL_41_1 gnd vdd FILL
XNOR2X1_511 NOR2X1_511/A AND2X2_51/B gnd NOR2X1_512/A vdd NOR2X1
XNOR2X1_544 AND2X2_46/B NOR2X1_676/A gnd OAI22X1_58/D vdd NOR2X1
XNOR2X1_522 BUFX4_266/Y NOR2X1_522/B gnd OAI22X1_49/D vdd NOR2X1
XNOR2X1_533 BUFX4_284/Y NOR2X1_683/A gnd NOR2X1_533/Y vdd NOR2X1
XNOR2X1_555 INVX1_17/A BUFX4_229/Y gnd OAI22X1_62/D vdd NOR2X1
XNOR2X1_566 NOR2X1_566/A BUFX4_153/Y gnd NOR2X1_566/Y vdd NOR2X1
XNOR2X1_577 INVX1_80/A BUFX4_270/Y gnd NOR2X1_577/Y vdd NOR2X1
XNOR2X1_599 NOR2X1_599/A BUFX4_329/Y gnd NOR2X1_599/Y vdd NOR2X1
XNOR2X1_588 NOR2X1_588/A BUFX4_284/Y gnd OAI22X1_74/D vdd NOR2X1
XAOI21X1_124 BUFX4_377/Y NOR2X1_703/B NOR2X1_199/Y gnd AOI21X1_124/Y vdd AOI21X1
XAOI21X1_113 BUFX4_466/Y INVX1_219/A NOR2X1_183/Y gnd AOI21X1_113/Y vdd AOI21X1
XAOI21X1_102 AND2X2_3/B NOR2X1_167/B NOR2X1_167/Y gnd AOI21X1_102/Y vdd AOI21X1
XAOI21X1_135 BUFX4_177/Y MUX2X1_376/S NOR2X1_215/Y gnd AOI21X1_135/Y vdd AOI21X1
XAOI21X1_157 BUFX4_176/Y NOR2X1_729/B NOR2X1_247/Y gnd AOI21X1_157/Y vdd AOI21X1
XAOI21X1_146 BUFX4_380/Y NOR2X1_231/B NOR2X1_230/Y gnd AOI21X1_146/Y vdd AOI21X1
XAOI21X1_168 BUFX4_372/Y NOR2X1_261/B NOR2X1_263/Y gnd DFFPOSX1_16/D vdd AOI21X1
XAOI21X1_179 BUFX4_173/Y NOR2X1_16/Y NOR2X1_276/Y gnd AOI21X1_179/Y vdd AOI21X1
XOAI21X1_1341 INVX1_370/Y NAND2X1_50/B NAND2X1_357/Y gnd DFFPOSX1_328/D vdd OAI21X1
XOAI21X1_1330 BUFX4_316/Y NAND2X1_44/Y OAI21X1_1329/Y gnd OAI21X1_1330/Y vdd OAI21X1
XDFFPOSX1_920 INVX1_115/A CLKBUF1_37/Y MUX2X1_102/Y gnd vdd DFFPOSX1
XOAI21X1_1363 NAND2X1_53/Y BUFX4_67/Y OAI21X1_1363/C gnd DFFPOSX1_308/D vdd OAI21X1
XOAI21X1_1374 BUFX4_385/Y BUFX4_131/Y INVX1_243/A gnd OAI21X1_1374/Y vdd OAI21X1
XOAI21X1_1352 NOR2X1_77/B BUFX4_184/Y OAI21X1_760/B gnd OAI21X1_1352/Y vdd OAI21X1
XDFFPOSX1_931 INVX1_288/A CLKBUF1_39/Y OAI21X1_233/Y gnd vdd DFFPOSX1
XDFFPOSX1_942 INVX1_126/A CLKBUF1_50/Y MUX2X1_113/Y gnd vdd DFFPOSX1
XDFFPOSX1_964 OAI21X1_900/A CLKBUF1_49/Y OAI21X1_259/Y gnd vdd DFFPOSX1
XDFFPOSX1_953 NOR2X1_514/A CLKBUF1_50/Y AOI21X1_116/Y gnd vdd DFFPOSX1
XOAI21X1_1385 BUFX4_426/Y NAND2X1_58/Y OAI21X1_1384/Y gnd OAI21X1_1385/Y vdd OAI21X1
XDFFPOSX1_975 NOR2X1_206/A CLKBUF1_15/Y AOI21X1_128/Y gnd vdd DFFPOSX1
XOAI21X1_1396 BUFX4_387/Y BUFX4_407/Y OAI21X1_1396/C gnd OAI21X1_1397/C vdd OAI21X1
XDFFPOSX1_986 NOR2X1_613/A CLKBUF1_102/Y AOI21X1_137/Y gnd vdd DFFPOSX1
XDFFPOSX1_997 INVX1_136/A CLKBUF1_44/Y MUX2X1_123/Y gnd vdd DFFPOSX1
XFILL_47_6_0 gnd vdd FILL
XFILL_30_5_0 gnd vdd FILL
XDFFPOSX1_227 INVX1_314/A CLKBUF1_93/Y MUX2X1_335/Y gnd vdd DFFPOSX1
XDFFPOSX1_216 NOR2X1_638/A CLKBUF1_65/Y AOI21X1_526/Y gnd vdd DFFPOSX1
XDFFPOSX1_205 NOR2X1_683/A CLKBUF1_45/Y AOI21X1_571/Y gnd vdd DFFPOSX1
XDFFPOSX1_249 DFFPOSX1_249/Q CLKBUF1_31/Y DFFPOSX1_249/D gnd vdd DFFPOSX1
XDFFPOSX1_238 NOR2X1_363/A CLKBUF1_43/Y OAI21X1_1266/Y gnd vdd DFFPOSX1
XNAND2X1_308 BUFX4_167/Y NAND2X1_308/B gnd NAND2X1_308/Y vdd NAND2X1
XNAND2X1_319 BUFX4_418/Y OAI22X1_45/Y gnd NAND2X1_319/Y vdd NAND2X1
XFILL_38_6_0 gnd vdd FILL
XBUFX4_281 BUFX4_17/Y gnd BUFX4_281/Y vdd BUFX4
XBUFX4_270 BUFX4_19/Y gnd BUFX4_270/Y vdd BUFX4
XNOR2X1_330 OR2X2_6/B INVX1_205/A gnd OAI22X1_2/A vdd NOR2X1
XNOR2X1_341 NOR2X1_341/A NOR2X1_341/B gnd NAND3X1_64/B vdd NOR2X1
XNOR2X1_352 NOR2X1_352/A XOR2X1_3/A gnd OAI22X1_3/D vdd NOR2X1
XBUFX4_292 INVX8_5/Y gnd BUFX4_292/Y vdd BUFX4
XNOR2X1_363 NOR2X1_363/A BUFX4_222/Y gnd NOR2X1_363/Y vdd NOR2X1
XNOR2X1_374 BUFX4_289/Y INVX1_12/Y gnd NOR2X1_374/Y vdd NOR2X1
XNOR2X1_385 BUFX4_207/Y NOR2X1_385/B gnd NOR2X1_385/Y vdd NOR2X1
XNOR2X1_396 NOR2X1_396/A BUFX4_283/Y gnd NOR2X1_396/Y vdd NOR2X1
XOAI21X1_814 NOR2X1_442/Y OAI21X1_814/B OAI21X1_813/Y gnd MUX2X1_217/B vdd OAI21X1
XOAI21X1_803 NOR2X1_436/Y OAI21X1_803/B OAI21X1_803/C gnd OAI21X1_804/A vdd OAI21X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_825 NOR2X1_445/Y AOI21X1_360/Y BUFX4_412/Y gnd OAI21X1_826/C vdd OAI21X1
XOAI21X1_858 INVX1_91/Y BUFX4_411/Y OAI21X1_858/C gnd NAND3X1_74/B vdd OAI21X1
XOAI21X1_836 INVX1_70/A BUFX4_261/Y BUFX4_100/Y gnd OAI21X1_836/Y vdd OAI21X1
XOAI21X1_847 BUFX4_417/Y OAI21X1_847/B NAND2X1_255/Y gnd AOI22X1_22/A vdd OAI21X1
XOAI21X1_869 OAI22X1_27/Y BUFX4_36/Y BUFX4_169/Y gnd OAI22X1_28/B vdd OAI21X1
XMUX2X1_303 INVX1_366/Y BUFX4_68/Y MUX2X1_66/S gnd MUX2X1_303/Y vdd MUX2X1
XMUX2X1_314 MUX2X1_6/B INVX1_295/Y MUX2X1_75/S gnd MUX2X1_314/Y vdd MUX2X1
XOAI21X1_1182 NOR2X1_59/A BUFX4_263/Y BUFX4_83/Y gnd OAI22X1_67/B vdd OAI21X1
XMUX2X1_325 INVX1_455/Y BUFX4_439/Y MUX2X1_84/S gnd MUX2X1_325/Y vdd MUX2X1
XMUX2X1_336 BUFX4_65/Y INVX1_355/Y MUX2X1_92/S gnd MUX2X1_336/Y vdd MUX2X1
XOAI21X1_1171 INVX1_439/Y BUFX4_256/Y BUFX4_79/Y gnd OAI21X1_1171/Y vdd OAI21X1
XOAI21X1_1160 INVX1_432/Y BUFX4_246/Y BUFX4_117/Y gnd OAI21X1_1160/Y vdd OAI21X1
XMUX2X1_347 BUFX4_66/Y INVX1_356/Y NOR2X1_172/B gnd MUX2X1_347/Y vdd MUX2X1
XDFFPOSX1_750 INVX1_64/A CLKBUF1_46/Y MUX2X1_54/Y gnd vdd DFFPOSX1
XMUX2X1_369 BUFX4_444/Y INVX1_254/Y MUX2X1_369/S gnd MUX2X1_369/Y vdd MUX2X1
XMUX2X1_358 INVX1_317/Y BUFX4_420/Y MUX2X1_360/S gnd MUX2X1_358/Y vdd MUX2X1
XDFFPOSX1_772 INVX1_70/A CLKBUF1_68/Y MUX2X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_783 OAI21X1_125/C CLKBUF1_55/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_761 NOR2X1_94/A CLKBUF1_54/Y AOI21X1_50/Y gnd vdd DFFPOSX1
XOAI21X1_1193 INVX1_68/Y BUFX4_274/Y NAND2X1_344/Y gnd MUX2X1_261/A vdd OAI21X1
XDFFPOSX1_794 NOR2X1_105/A CLKBUF1_58/Y AOI21X1_58/Y gnd vdd DFFPOSX1
XFILL_4_6_0 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XNAND3X1_81 BUFX4_36/Y NAND3X1_81/B NAND3X1_81/C gnd NAND3X1_81/Y vdd NAND3X1
XNAND3X1_70 INVX1_215/Y NAND3X1_70/B AND2X2_16/A gnd OR2X2_7/A vdd NAND3X1
XNOR2X1_70 BUFX4_46/Y BUFX4_191/Y gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_81 NOR2X1_81/A NOR2X1_83/B gnd NOR2X1_81/Y vdd NOR2X1
XNOR2X1_92 NOR2X1_92/A NOR2X1_92/B gnd NOR2X1_92/Y vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd traffic_Street[3] vdd BUFX2
XNAND2X1_105 NAND3X1_7/Y NAND2X1_105/B gnd NOR3X1_3/A vdd NAND2X1
XNAND2X1_116 INVX1_188/A INVX1_191/Y gnd NAND2X1_116/Y vdd NAND2X1
XNAND2X1_149 NAND3X1_46/Y OAI21X1_500/Y gnd NAND3X1_56/A vdd NAND2X1
XNAND2X1_138 AND2X2_9/A AND2X2_9/B gnd AOI21X1_241/C vdd NAND2X1
XNAND2X1_127 INVX2_18/A NOR2X1_319/Y gnd AOI21X1_224/A vdd NAND2X1
XNAND2X1_3 NAND2X1_3/A NAND2X1_2/Y gnd NAND2X1_3/Y vdd NAND2X1
XNOR2X1_160 NOR2X1_160/A MUX2X1_340/S gnd NOR2X1_160/Y vdd NOR2X1
XNOR2X1_171 NOR2X1_171/A NOR2X1_172/B gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_193 NOR2X1_464/A MUX2X1_364/S gnd NOR2X1_193/Y vdd NOR2X1
XNOR2X1_182 NOR2X1_182/A INVX1_219/A gnd NOR2X1_182/Y vdd NOR2X1
XOAI21X1_611 INVX1_266/Y BUFX4_282/Y OAI21X1_611/C gnd MUX2X1_185/B vdd OAI21X1
XOAI21X1_622 INVX1_8/Y BUFX4_332/Y OAI21X1_622/C gnd NAND3X1_72/B vdd OAI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XOAI21X1_633 BUFX4_31/Y MUX2X1_189/Y OAI21X1_633/C gnd AOI22X1_16/C vdd OAI21X1
XOAI21X1_600 AND2X2_29/A OAI21X1_600/B BUFX4_98/Y gnd AOI21X1_276/C vdd OAI21X1
XOAI21X1_666 INVX1_127/Y BUFX4_369/Y OAI21X1_666/C gnd AOI21X1_303/B vdd OAI21X1
XAOI21X1_8 BUFX4_442/Y NOR2X1_30/B AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XOAI21X1_655 INVX1_282/Y BUFX4_255/Y OAI21X1_655/C gnd MUX2X1_198/B vdd OAI21X1
XOAI21X1_644 MUX2X1_193/Y BUFX4_415/Y BUFX4_170/Y gnd OAI21X1_645/A vdd OAI21X1
XOAI21X1_699 BUFX4_352/Y NOR2X1_55/A BUFX4_157/Y gnd OAI22X1_16/C vdd OAI21X1
XOAI21X1_677 BUFX4_327/Y OAI21X1_677/B BUFX4_153/Y gnd OAI22X1_13/C vdd OAI21X1
XOAI21X1_688 NOR2X1_395/Y AOI21X1_308/Y BUFX4_394/Y gnd OAI21X1_688/Y vdd OAI21X1
XMUX2X1_111 INVX1_124/Y MUX2X1_96/A MUX2X1_360/S gnd MUX2X1_111/Y vdd MUX2X1
XMUX2X1_100 INVX1_113/Y BUFX4_466/Y MUX2X1_97/S gnd MUX2X1_100/Y vdd MUX2X1
XMUX2X1_122 BUFX4_216/Y INVX1_135/Y NOR2X1_220/B gnd MUX2X1_122/Y vdd MUX2X1
XMUX2X1_133 BUFX4_180/Y INVX1_146/Y MUX2X1_397/S gnd DFFPOSX1_3/D vdd MUX2X1
XMUX2X1_155 INVX1_168/Y BUFX4_178/Y MUX2X1_14/S gnd MUX2X1_155/Y vdd MUX2X1
XMUX2X1_144 INVX1_157/Y MUX2X1_61/B MUX2X1_2/S gnd MUX2X1_144/Y vdd MUX2X1
XDFFPOSX1_591 NAND2X1_361/A CLKBUF1_40/Y DFFPOSX1_591/D gnd vdd DFFPOSX1
XDFFPOSX1_580 INVX1_329/A CLKBUF1_35/Y MUX2X1_409/Y gnd vdd DFFPOSX1
XMUX2X1_188 MUX2X1_188/A MUX2X1_188/B BUFX4_109/Y gnd MUX2X1_188/Y vdd MUX2X1
XMUX2X1_199 MUX2X1_199/A OAI22X1_8/Y INVX8_33/Y gnd MUX2X1_199/Y vdd MUX2X1
XMUX2X1_177 MUX2X1_177/A MUX2X1_177/B BUFX4_80/Y gnd MUX2X1_177/Y vdd MUX2X1
XMUX2X1_166 INVX1_180/Y MUX2X1_71/B MUX2X1_29/S gnd MUX2X1_166/Y vdd MUX2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XFILL_45_9_1 gnd vdd FILL
XFILL_44_4_0 gnd vdd FILL
XDFFPOSX1_3 INVX1_146/A CLKBUF1_90/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XNOR2X1_6 INVX2_1/Y NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_35_4_0 gnd vdd FILL
XFILL_36_9_1 gnd vdd FILL
XAOI21X1_16 MUX2X1_27/B NOR2X1_43/B NOR2X1_41/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_27 BUFX4_473/Y NOR2X1_57/Y NOR2X1_59/Y gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_38 MUX2X1_39/B NOR2X1_76/B NOR2X1_75/Y gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_49 MUX2X1_64/B NOR2X1_92/B NOR2X1_93/Y gnd AOI21X1_49/Y vdd AOI21X1
XFILL_2_9_1 gnd vdd FILL
XFILL_27_9_1 gnd vdd FILL
XFILL_1_4_0 gnd vdd FILL
XFILL_26_4_0 gnd vdd FILL
XOAI22X1_13 OAI22X1_13/A OAI22X1_13/B OAI22X1_13/C OAI22X1_13/D gnd OAI22X1_13/Y vdd
+ OAI22X1
XOAI22X1_24 OAI22X1_24/A OAI22X1_24/B MUX2X1_217/Y AND2X2_48/B gnd OAI22X1_24/Y vdd
+ OAI22X1
XOAI22X1_57 OAI22X1_57/A OAI22X1_57/B OAI22X1_57/C NOR2X1_542/Y gnd OAI22X1_57/Y vdd
+ OAI22X1
XOAI22X1_46 BUFX4_48/Y MUX2X1_253/Y OAI22X1_46/C NOR2X1_507/Y gnd OAI22X1_46/Y vdd
+ OAI22X1
XOAI22X1_35 OAI22X1_35/A OAI22X1_35/B OAI22X1_35/C OAI22X1_35/D gnd OAI22X1_35/Y vdd
+ OAI22X1
XOAI22X1_68 NOR2X1_575/Y OAI22X1_68/B OAI22X1_68/C OAI22X1_68/D gnd OAI22X1_68/Y vdd
+ OAI22X1
XOAI22X1_79 NOR2X1_599/Y OAI22X1_79/B OAI22X1_79/C NOR2X1_598/Y gnd OAI22X1_79/Y vdd
+ OAI22X1
XOAI21X1_441 OAI21X1_441/A AOI22X1_2/Y NAND3X1_8/B gnd NAND3X1_7/C vdd OAI21X1
XFILL_10_8_1 gnd vdd FILL
XOAI21X1_430 BUFX4_209/Y OAI21X1_64/B OAI21X1_429/Y gnd OAI21X1_430/Y vdd OAI21X1
XOAI21X1_452 NOR2X1_304/Y BUFX4_73/Y AND2X2_6/B gnd NAND3X1_15/C vdd OAI21X1
XOAI21X1_463 NAND2X1_168/A INVX2_15/A OAI21X1_463/C gnd AOI21X1_215/C vdd OAI21X1
XOAI21X1_474 BUFX4_320/Y NOR2X1_351/B NAND3X1_16/C gnd INVX2_19/A vdd OAI21X1
XOAI21X1_496 INVX1_205/A OR2X2_6/B NOR3X1_1/B gnd AOI22X1_6/B vdd OAI21X1
XOAI21X1_485 INVX1_201/A INVX1_196/A NOR3X1_4/B gnd INVX2_23/A vdd OAI21X1
XFILL_9_5_0 gnd vdd FILL
XFILL_18_9_1 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XAOI21X1_509 BUFX4_415/Y MUX2X1_265/Y BUFX4_201/Y gnd AOI21X1_509/Y vdd AOI21X1
XFILL_50_2_0 gnd vdd FILL
XOAI21X1_90 NAND2X1_32/Y BUFX4_468/Y OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XFILL_41_2_0 gnd vdd FILL
XFILL_42_7_1 gnd vdd FILL
XOAI21X1_260 BUFX4_126/Y BUFX4_432/Y OAI21X1_260/C gnd OAI21X1_260/Y vdd OAI21X1
XOAI21X1_282 BUFX4_192/Y BUFX4_162/Y NOR2X1_470/A gnd OAI21X1_282/Y vdd OAI21X1
XOAI21X1_271 NAND2X1_72/Y BUFX4_465/Y OAI21X1_270/Y gnd OAI21X1_271/Y vdd OAI21X1
XINVX1_313 INVX1_313/A gnd INVX1_313/Y vdd INVX1
XOAI21X1_293 NAND2X1_75/Y BUFX4_380/Y OAI21X1_293/C gnd OAI21X1_293/Y vdd OAI21X1
XINVX1_324 INVX1_324/A gnd INVX1_324/Y vdd INVX1
XINVX1_302 INVX1_302/A gnd INVX1_302/Y vdd INVX1
XINVX1_335 INVX1_335/A gnd INVX1_335/Y vdd INVX1
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XINVX1_346 INVX1_346/A gnd INVX1_346/Y vdd INVX1
XINVX1_357 INVX1_357/A gnd INVX1_357/Y vdd INVX1
XINVX1_379 INVX1_379/A gnd INVX1_379/Y vdd INVX1
XFILL_49_3_0 gnd vdd FILL
XNOR2X1_726 NOR2X1_726/A NOR2X1_234/Y gnd NOR2X1_726/Y vdd NOR2X1
XNOR2X1_715 NOR2X1_715/A NOR2X1_716/B gnd NOR2X1_715/Y vdd NOR2X1
XNOR2X1_704 NOR2X1_704/A NOR2X1_703/B gnd NOR2X1_704/Y vdd NOR2X1
XNOR2X1_737 NOR2X1_737/A NOR2X1_737/B gnd NOR2X1_737/Y vdd NOR2X1
XFILL_32_2_0 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XAOI21X1_306 NOR2X1_214/A BUFX4_274/Y AOI21X1_306/C gnd OAI21X1_675/B vdd AOI21X1
XAOI21X1_328 AOI21X1_328/A NOR2X1_419/Y OAI21X1_745/Y gnd AOI21X1_328/Y vdd AOI21X1
XAOI21X1_339 INVX8_33/Y AOI21X1_339/B AOI21X1_339/C gnd AOI21X1_339/Y vdd AOI21X1
XAOI21X1_317 INVX4_14/Y MUX2X1_207/Y INVX4_13/Y gnd AOI22X1_18/C vdd AOI21X1
XOAI21X1_1512 BUFX4_322/Y NAND2X1_77/Y OAI21X1_1511/Y gnd OAI21X1_1512/Y vdd OAI21X1
XDFFPOSX1_16 NOR2X1_263/A CLKBUF1_35/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XDFFPOSX1_27 INVX1_152/A CLKBUF1_11/Y MUX2X1_139/Y gnd vdd DFFPOSX1
XOAI21X1_1523 BUFX4_389/Y BUFX4_313/Y OAI21X1_791/B gnd OAI21X1_1524/C vdd OAI21X1
XOAI21X1_1501 NOR2X1_77/B BUFX4_457/Y NOR2X1_484/A gnd OAI21X1_1502/C vdd OAI21X1
XOAI21X1_1545 BUFX4_385/Y BUFX4_195/Y OAI21X1_613/B gnd OAI21X1_1546/C vdd OAI21X1
XOAI21X1_1534 NAND2X1_80/Y BUFX4_67/Y OAI21X1_1534/C gnd DFFPOSX1_545/D vdd OAI21X1
XOAI21X1_1556 NAND2X1_84/Y BUFX4_426/Y OAI21X1_1556/C gnd OAI21X1_1556/Y vdd OAI21X1
XDFFPOSX1_49 INVX1_158/A CLKBUF1_66/Y MUX2X1_145/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 NAND2X1_198/A CLKBUF1_11/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XOAI21X1_1567 BUFX4_191/Y BUFX4_196/Y NOR2X1_551/A gnd OAI21X1_1568/C vdd OAI21X1
XFILL_23_2_0 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_7_8_1 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XCLKBUF1_91 BUFX4_7/Y gnd CLKBUF1_91/Y vdd CLKBUF1
XCLKBUF1_80 BUFX4_7/Y gnd CLKBUF1_80/Y vdd CLKBUF1
XFILL_15_7_1 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XDFFPOSX1_409 INVX1_420/A CLKBUF1_27/Y MUX2X1_345/Y gnd vdd DFFPOSX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XCLKBUF1_102 BUFX4_10/Y gnd CLKBUF1_102/Y vdd CLKBUF1
XBUFX4_430 INVX8_3/Y gnd BUFX4_430/Y vdd BUFX4
XBUFX4_474 INVX8_15/Y gnd AND2X2_3/B vdd BUFX4
XBUFX4_441 INVX8_2/Y gnd BUFX4_441/Y vdd BUFX4
XNOR2X1_501 NOR2X1_501/A BUFX4_278/Y gnd NOR2X1_502/A vdd NOR2X1
XBUFX4_452 BUFX4_449/A gnd BUFX4_452/Y vdd BUFX4
XBUFX4_463 INVX8_10/Y gnd NOR2X1_39/A vdd BUFX4
XNOR2X1_512 NOR2X1_512/A NOR2X1_512/B gnd NOR2X1_512/Y vdd NOR2X1
XNOR2X1_523 NOR2X1_523/A BUFX4_334/Y gnd OAI22X1_49/A vdd NOR2X1
XNOR2X1_534 NOR2X1_534/A BUFX4_335/Y gnd NOR2X1_534/Y vdd NOR2X1
XFILL_41_2 gnd vdd FILL
XNOR2X1_556 NAND2X1_14/A BUFX4_363/Y gnd OAI22X1_62/A vdd NOR2X1
XNOR2X1_545 NOR2X1_545/A BUFX4_354/Y gnd NOR2X1_545/Y vdd NOR2X1
XNOR2X1_567 BUFX4_77/Y NOR2X1_567/B gnd NOR2X1_567/Y vdd NOR2X1
XNOR2X1_578 BUFX4_416/Y NOR2X1_578/B gnd NOR2X1_578/Y vdd NOR2X1
XNOR2X1_589 NOR2X1_589/A BUFX4_342/Y gnd OAI22X1_74/A vdd NOR2X1
XAOI21X1_114 MUX2X1_97/B NOR2X1_188/B NOR2X1_187/Y gnd AOI21X1_114/Y vdd AOI21X1
XAOI21X1_103 BUFX4_216/Y NOR2X1_172/B NOR2X1_170/Y gnd AOI21X1_103/Y vdd AOI21X1
XAOI21X1_125 BUFX4_466/Y NOR2X1_703/B NOR2X1_200/Y gnd AOI21X1_125/Y vdd AOI21X1
XAOI21X1_158 BUFX4_380/Y NOR2X1_729/B NOR2X1_248/Y gnd AOI21X1_158/Y vdd AOI21X1
XAOI21X1_147 BUFX4_465/Y NOR2X1_231/B NOR2X1_231/Y gnd AOI21X1_147/Y vdd AOI21X1
XAOI21X1_136 BUFX4_377/Y MUX2X1_376/S NOR2X1_216/Y gnd AOI21X1_136/Y vdd AOI21X1
XAOI21X1_169 BUFX4_473/Y NOR2X1_261/B NOR2X1_264/Y gnd DFFPOSX1_17/D vdd AOI21X1
XOAI21X1_1331 INVX1_415/Y NOR2X1_107/B NAND2X1_355/Y gnd OAI21X1_1331/Y vdd OAI21X1
XOAI21X1_1320 BUFX4_449/Y BUFX4_55/Y NOR2X1_530/B gnd OAI21X1_1321/C vdd OAI21X1
XDFFPOSX1_910 INVX1_113/A CLKBUF1_27/Y MUX2X1_100/Y gnd vdd DFFPOSX1
XOAI21X1_1364 BUFX4_454/Y BUFX4_186/Y NOR2X1_542/B gnd OAI21X1_1365/C vdd OAI21X1
XOAI21X1_1342 BUFX4_59/Y BUFX4_187/Y NAND2X1_177/B gnd OAI21X1_1343/C vdd OAI21X1
XOAI21X1_1353 NAND2X1_52/Y BUFX4_428/Y OAI21X1_1352/Y gnd OAI21X1_1353/Y vdd OAI21X1
XDFFPOSX1_921 NOR2X1_175/A CLKBUF1_12/Y AOI21X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_932 AND2X2_33/A CLKBUF1_29/Y OAI21X1_235/Y gnd vdd DFFPOSX1
XDFFPOSX1_943 OAI21X1_667/B CLKBUF1_9/Y OAI21X1_241/Y gnd vdd DFFPOSX1
XDFFPOSX1_965 OAI21X1_260/C CLKBUF1_49/Y OAI21X1_261/Y gnd vdd DFFPOSX1
XDFFPOSX1_976 NOR2X1_207/A CLKBUF1_102/Y AOI21X1_129/Y gnd vdd DFFPOSX1
XDFFPOSX1_954 NOR2X1_190/A CLKBUF1_9/Y AOI21X1_117/Y gnd vdd DFFPOSX1
XOAI21X1_1375 NAND2X1_57/Y BUFX4_441/Y OAI21X1_1374/Y gnd DFFPOSX1_270/D vdd OAI21X1
XOAI21X1_1386 BUFX4_136/Y BUFX4_127/Y OAI21X1_924/B gnd OAI21X1_1386/Y vdd OAI21X1
XOAI21X1_1397 NAND2X1_59/Y BUFX4_320/Y OAI21X1_1397/C gnd DFFPOSX1_197/D vdd OAI21X1
XDFFPOSX1_987 INVX1_284/A CLKBUF1_67/Y OAI21X1_265/Y gnd vdd DFFPOSX1
XDFFPOSX1_998 NOR2X1_220/A CLKBUF1_7/Y AOI21X1_139/Y gnd vdd DFFPOSX1
XFILL_47_6_1 gnd vdd FILL
XFILL_46_1_0 gnd vdd FILL
XFILL_30_5_1 gnd vdd FILL
XDFFPOSX1_228 INVX1_355/A CLKBUF1_93/Y MUX2X1_336/Y gnd vdd DFFPOSX1
XDFFPOSX1_206 AND2X2_21/B CLKBUF1_23/Y DFFPOSX1_206/D gnd vdd DFFPOSX1
XDFFPOSX1_217 NOR2X1_639/A CLKBUF1_38/Y AOI21X1_527/Y gnd vdd DFFPOSX1
XDFFPOSX1_239 NOR2X1_420/B CLKBUF1_94/Y DFFPOSX1_239/D gnd vdd DFFPOSX1
XNAND2X1_309 NOR2X1_63/A AND2X2_29/A gnd NAND2X1_309/Y vdd NAND2X1
XFILL_37_1_0 gnd vdd FILL
XFILL_38_6_1 gnd vdd FILL
XBUFX4_260 BUFX4_21/Y gnd BUFX4_260/Y vdd BUFX4
XBUFX4_271 BUFX4_23/Y gnd BUFX4_271/Y vdd BUFX4
XBUFX4_282 BUFX4_19/Y gnd BUFX4_282/Y vdd BUFX4
XNOR2X1_331 NOR3X1_1/B AND2X2_3/Y gnd NOR2X1_331/Y vdd NOR2X1
XNOR2X1_320 INVX2_20/Y BUFX4_305/Y gnd AOI22X1_9/C vdd NOR2X1
XNOR2X1_342 INVX2_23/A INVX4_12/A gnd NOR2X1_342/Y vdd NOR2X1
XBUFX4_293 INVX8_5/Y gnd BUFX4_293/Y vdd BUFX4
XNOR2X1_386 NOR2X1_192/A AND2X2_23/A gnd NOR2X1_386/Y vdd NOR2X1
XNOR2X1_353 AND2X2_5/B AOI22X1_5/D gnd NOR2X1_353/Y vdd NOR2X1
XNOR2X1_364 NOR2X1_363/Y NOR2X1_364/B gnd NOR2X1_364/Y vdd NOR2X1
XNOR2X1_375 OAI21X1_35/C BUFX4_229/Y gnd OAI22X1_6/D vdd NOR2X1
XNOR2X1_397 NOR2X1_397/A BUFX4_356/Y gnd NOR2X1_397/Y vdd NOR2X1
XOAI21X1_815 BUFX4_360/Y NOR2X1_29/A BUFX4_149/Y gnd OAI21X1_815/Y vdd OAI21X1
XFILL_20_0_0 gnd vdd FILL
XOAI21X1_804 OAI21X1_804/A INVX8_30/A BUFX4_201/Y gnd OAI21X1_805/B vdd OAI21X1
XFILL_21_5_1 gnd vdd FILL
XOAI21X1_826 AOI21X1_359/Y BUFX4_413/Y OAI21X1_826/C gnd MUX2X1_218/A vdd OAI21X1
XOAI21X1_837 BUFX4_353/Y INVX1_90/A BUFX4_158/Y gnd AOI21X1_366/C vdd OAI21X1
XOAI21X1_848 INVX1_111/Y BUFX4_106/Y BUFX4_344/Y gnd OAI21X1_850/B vdd OAI21X1
XOAI21X1_859 AOI21X1_376/Y OAI21X1_859/B NAND3X1_74/Y gnd MUX2X1_222/A vdd OAI21X1
XMUX2X1_304 INVX1_451/Y MUX2X1_29/B MUX2X1_66/S gnd MUX2X1_304/Y vdd MUX2X1
XMUX2X1_348 BUFX4_317/Y INVX1_419/Y NOR2X1_172/B gnd MUX2X1_348/Y vdd MUX2X1
XMUX2X1_337 AND2X2_5/B INVX1_241/Y MUX2X1_96/S gnd MUX2X1_337/Y vdd MUX2X1
XMUX2X1_326 INVX1_456/Y BUFX4_424/Y MUX2X1_84/S gnd MUX2X1_326/Y vdd MUX2X1
XOAI21X1_1183 BUFX4_352/Y NOR2X1_69/A BUFX4_157/Y gnd OAI22X1_68/C vdd OAI21X1
XDFFPOSX1_740 AND2X2_31/A CLKBUF1_85/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XOAI21X1_1172 OAI21X1_1171/Y AND2X2_53/Y OAI21X1_1170/Y gnd MUX2X1_260/B vdd OAI21X1
XOAI21X1_1161 OAI21X1_1160/Y AND2X2_52/Y OAI21X1_1159/Y gnd MUX2X1_258/B vdd OAI21X1
XMUX2X1_315 INVX1_232/Y BUFX4_443/Y MUX2X1_76/S gnd MUX2X1_315/Y vdd MUX2X1
XOAI21X1_1150 BUFX4_113/Y AOI21X1_481/Y OAI21X1_1150/C gnd OAI21X1_1151/A vdd OAI21X1
XMUX2X1_359 INVX1_379/Y BUFX4_70/Y MUX2X1_360/S gnd MUX2X1_359/Y vdd MUX2X1
XOAI21X1_1194 BUFX4_355/Y NOR2X1_100/A BUFX4_156/Y gnd OAI22X1_70/C vdd OAI21X1
XDFFPOSX1_773 INVX1_71/A CLKBUF1_55/Y MUX2X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_784 OAI21X1_839/B CLKBUF1_51/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XDFFPOSX1_751 NAND2X1_224/A CLKBUF1_15/Y OAI21X1_110/Y gnd vdd DFFPOSX1
XDFFPOSX1_762 NOR2X1_95/A CLKBUF1_46/Y AOI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_795 INVX1_86/A CLKBUF1_77/Y MUX2X1_76/Y gnd vdd DFFPOSX1
XFILL_4_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNAND3X1_60 INVX4_10/Y XOR2X1_2/Y NAND3X1_54/C gnd NAND3X1_60/Y vdd NAND3X1
XNAND3X1_82 INVX8_28/A NAND3X1_82/B NAND3X1_82/C gnd NAND3X1_82/Y vdd NAND3X1
XNAND3X1_71 BUFX4_40/Y NAND3X1_71/B NAND3X1_71/C gnd AOI22X1_11/A vdd NAND3X1
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_60 BUFX4_42/Y BUFX4_144/Y gnd NOR2X1_60/Y vdd NOR2X1
XNOR2X1_71 NOR2X1_71/A NOR2X1_70/Y gnd NOR2X1_71/Y vdd NOR2X1
XNOR2X1_82 NOR2X1_82/A NOR2X1_83/B gnd NOR2X1_82/Y vdd NOR2X1
XNOR2X1_93 NOR2X1_93/A NOR2X1_92/B gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd west_East[0] vdd BUFX2
XNAND2X1_106 OR2X2_2/A NAND2X1_106/B gnd NAND3X1_11/C vdd NAND2X1
XNAND2X1_117 INVX1_193/A AND2X2_5/A gnd NAND2X1_117/Y vdd NAND2X1
XNAND2X1_139 NAND3X1_8/B NAND3X1_8/C gnd INVX2_24/A vdd NAND2X1
XNAND2X1_128 INVX2_14/A NOR2X1_312/Y gnd NOR2X1_321/B vdd NAND2X1
XNAND2X1_4 NOR2X1_8/Y NOR2X1_6/Y gnd NAND2X1_6/B vdd NAND2X1
XNOR2X1_161 MUX2X1_247/A MUX2X1_340/S gnd AOI21X1_97/C vdd NOR2X1
XNOR2X1_150 INVX4_2/A BUFX4_406/Y gnd MUX2X1_96/S vdd NOR2X1
XNOR2X1_172 NOR2X1_172/A NOR2X1_172/B gnd NOR2X1_172/Y vdd NOR2X1
XNOR2X1_194 NOR2X1_511/A MUX2X1_364/S gnd NOR2X1_194/Y vdd NOR2X1
XNOR2X1_183 NOR2X1_183/A INVX1_219/A gnd NOR2X1_183/Y vdd NOR2X1
XOAI21X1_612 INVX1_267/Y BUFX4_284/Y NAND2X1_188/Y gnd MUX2X1_185/A vdd OAI21X1
XOAI21X1_623 INVX1_4/Y BUFX4_346/Y AOI21X1_291/Y gnd NAND3X1_72/C vdd OAI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XOAI21X1_601 OAI21X1_601/A OAI21X1_601/B BUFX4_35/Y gnd AOI21X1_279/A vdd OAI21X1
XOAI21X1_656 INVX1_145/Y BUFX4_257/Y OAI21X1_656/C gnd MUX2X1_198/A vdd OAI21X1
XOAI21X1_634 INVX1_159/Y BUFX4_414/Y AOI21X1_294/Y gnd OAI21X1_634/Y vdd OAI21X1
XOAI21X1_645 OAI21X1_645/A NOR2X1_378/Y BUFX4_390/Y gnd OAI22X1_8/B vdd OAI21X1
XOAI21X1_667 BUFX4_359/Y OAI21X1_667/B BUFX4_147/Y gnd OAI22X1_11/C vdd OAI21X1
XAOI21X1_9 MUX2X1_6/B NOR2X1_30/B NOR2X1_29/Y gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_678 OAI21X1_678/A BUFX4_276/Y BUFX4_82/Y gnd OAI22X1_13/B vdd OAI21X1
XOAI21X1_689 INVX1_285/Y AND2X2_36/B NAND2X1_216/Y gnd MUX2X1_201/B vdd OAI21X1
XMUX2X1_112 INVX1_125/Y BUFX4_377/Y MUX2X1_360/S gnd MUX2X1_112/Y vdd MUX2X1
XMUX2X1_101 MUX2X1_57/A INVX1_114/Y NOR2X1_172/B gnd MUX2X1_101/Y vdd MUX2X1
XMUX2X1_123 BUFX4_380/Y INVX1_136/Y NOR2X1_220/B gnd MUX2X1_123/Y vdd MUX2X1
XMUX2X1_134 MUX2X1_86/B INVX1_147/Y MUX2X1_397/S gnd DFFPOSX1_4/D vdd MUX2X1
XMUX2X1_156 INVX1_169/Y BUFX4_375/Y MUX2X1_14/S gnd MUX2X1_156/Y vdd MUX2X1
XMUX2X1_145 INVX1_158/Y BUFX4_470/Y MUX2X1_2/S gnd MUX2X1_145/Y vdd MUX2X1
XMUX2X1_167 INVX1_181/Y BUFX4_177/Y MUX2X1_29/S gnd MUX2X1_167/Y vdd MUX2X1
XDFFPOSX1_570 DFFPOSX1_570/Q CLKBUF1_5/Y DFFPOSX1_570/D gnd vdd DFFPOSX1
XDFFPOSX1_592 NAND2X1_362/A CLKBUF1_81/Y DFFPOSX1_592/D gnd vdd DFFPOSX1
XDFFPOSX1_581 INVX1_391/A CLKBUF1_78/Y MUX2X1_410/Y gnd vdd DFFPOSX1
XMUX2X1_189 MUX2X1_189/A MUX2X1_189/B BUFX4_110/Y gnd MUX2X1_189/Y vdd MUX2X1
XMUX2X1_178 MUX2X1_178/A MUX2X1_178/B BUFX4_31/Y gnd AOI22X1_12/B vdd MUX2X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XFILL_44_4_1 gnd vdd FILL
XDFFPOSX1_4 INVX1_147/A CLKBUF1_52/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XNOR2X1_7 NOR2X1_1/B INVX2_4/Y gnd INVX2_5/A vdd NOR2X1
XFILL_35_4_1 gnd vdd FILL
XAOI21X1_17 BUFX4_70/Y NOR2X1_43/B NOR2X1_42/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 BUFX4_213/Y NOR2X1_60/Y NOR2X1_61/Y gnd AOI21X1_28/Y vdd AOI21X1
XAOI21X1_39 MUX2X1_44/A NOR2X1_76/B NOR2X1_76/Y gnd AOI21X1_39/Y vdd AOI21X1
XFILL_1_4_1 gnd vdd FILL
XFILL_26_4_1 gnd vdd FILL
XOAI22X1_14 NOR2X1_397/Y OAI22X1_14/B OAI22X1_14/C NOR2X1_396/Y gnd OAI22X1_14/Y vdd
+ OAI22X1
XOAI22X1_25 OAI22X1_25/A OAI22X1_25/B OAI22X1_25/C OAI22X1_25/D gnd OAI22X1_25/Y vdd
+ OAI22X1
XOAI22X1_47 NOR2X1_514/Y OAI22X1_47/B OAI22X1_47/C OAI22X1_47/D gnd OAI22X1_47/Y vdd
+ OAI22X1
XOAI22X1_58 NOR2X1_545/Y OAI22X1_58/B OAI22X1_58/C OAI22X1_58/D gnd OAI22X1_58/Y vdd
+ OAI22X1
XOAI22X1_36 OAI22X1_36/A OAI22X1_36/B OAI22X1_36/C OAI22X1_36/D gnd OAI22X1_36/Y vdd
+ OAI22X1
XOAI22X1_69 NOR2X1_573/Y OAI22X1_69/B OAI22X1_69/C NOR2X1_570/Y gnd OAI22X1_69/Y vdd
+ OAI22X1
XOAI21X1_431 BUFX4_190/Y BUFX4_461/Y NAND2X1_261/A gnd OAI21X1_431/Y vdd OAI21X1
XOAI21X1_420 MUX2X1_66/B OAI21X1_48/B OAI21X1_419/Y gnd OAI21X1_420/Y vdd OAI21X1
XOAI21X1_475 AND2X2_2/Y NOR2X1_301/Y INVX4_7/Y gnd OAI21X1_475/Y vdd OAI21X1
XOAI21X1_442 AND2X2_2/Y NOR2X1_301/Y INVX4_7/A gnd NAND3X1_9/C vdd OAI21X1
XOAI21X1_453 AOI21X1_208/Y AOI21X1_207/Y NAND3X1_17/B gnd NAND3X1_16/C vdd OAI21X1
XOAI21X1_464 NOR3X1_4/C INVX2_15/Y INVX1_193/Y gnd AOI21X1_215/B vdd OAI21X1
XOAI21X1_497 OAI21X1_497/A INVX4_12/A AOI22X1_6/D gnd OAI21X1_497/Y vdd OAI21X1
XOAI21X1_486 INVX4_12/Y INVX2_23/Y OAI21X1_497/A gnd INVX1_199/A vdd OAI21X1
XFILL_9_5_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XFILL_17_4_1 gnd vdd FILL
XFILL_50_2_1 gnd vdd FILL
XOAI21X1_80 NAND2X1_31/Y BUFX4_372/Y OAI21X1_79/Y gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 INVX1_47/Y NOR2X1_76/B NAND2X1_33/Y gnd OAI21X1_91/Y vdd OAI21X1
XFILL_41_2_1 gnd vdd FILL
XOAI21X1_250 BUFX4_384/Y BUFX4_434/Y OAI21X1_898/A gnd OAI21X1_250/Y vdd OAI21X1
XOAI21X1_261 NAND2X1_70/Y BUFX4_377/Y OAI21X1_260/Y gnd OAI21X1_261/Y vdd OAI21X1
XOAI21X1_272 BUFX4_132/Y BUFX4_162/Y AOI21X1_304/A gnd OAI21X1_272/Y vdd OAI21X1
XOAI21X1_283 BUFX4_174/Y NAND2X1_74/Y OAI21X1_282/Y gnd OAI21X1_283/Y vdd OAI21X1
XINVX1_314 INVX1_314/A gnd INVX1_314/Y vdd INVX1
XINVX1_303 INVX1_303/A gnd INVX1_303/Y vdd INVX1
XOAI21X1_294 BUFX4_457/Y BUFX4_298/Y NOR2X1_621/A gnd OAI21X1_294/Y vdd OAI21X1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XINVX1_336 INVX1_336/A gnd INVX1_336/Y vdd INVX1
XAND2X2_50 AND2X2_50/A BUFX4_410/Y gnd AND2X2_50/Y vdd AND2X2
XINVX1_347 INVX1_347/A gnd INVX1_347/Y vdd INVX1
XINVX1_358 INVX1_358/A gnd INVX1_358/Y vdd INVX1
XINVX1_369 INVX1_369/A gnd INVX1_369/Y vdd INVX1
XFILL_49_3_1 gnd vdd FILL
XNOR2X1_705 NOR2X1_705/A NOR2X1_703/B gnd NOR2X1_705/Y vdd NOR2X1
XNOR2X1_716 NOR2X1_716/A NOR2X1_716/B gnd NOR2X1_716/Y vdd NOR2X1
XNOR2X1_738 NOR2X1_738/A NOR2X1_737/B gnd NOR2X1_738/Y vdd NOR2X1
XNOR2X1_727 NOR2X1_727/A NOR2X1_727/B gnd NOR2X1_727/Y vdd NOR2X1
XAOI21X1_307 BUFX4_83/Y INVX1_93/Y BUFX4_277/Y gnd AOI21X1_307/Y vdd AOI21X1
XFILL_32_2_1 gnd vdd FILL
XAOI21X1_318 BUFX4_101/Y INVX1_293/Y NOR2X1_412/Y gnd AOI21X1_318/Y vdd AOI21X1
XAOI21X1_329 BUFX4_265/Y NOR2X1_697/A BUFX4_113/Y gnd AOI21X1_329/Y vdd AOI21X1
XDFFPOSX1_17 NOR2X1_264/A CLKBUF1_72/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XOAI21X1_1513 BUFX4_311/Y BUFX4_298/Y MUX2X1_182/B gnd OAI21X1_1513/Y vdd OAI21X1
XOAI21X1_1502 NAND2X1_76/Y BUFX4_72/Y OAI21X1_1502/C gnd DFFPOSX1_505/D vdd OAI21X1
XOAI21X1_1546 NAND2X1_82/Y BUFX4_441/Y OAI21X1_1546/C gnd DFFPOSX1_567/D vdd OAI21X1
XDFFPOSX1_28 INVX1_153/A CLKBUF1_35/Y MUX2X1_140/Y gnd vdd DFFPOSX1
XOAI21X1_1535 BUFX4_451/Y BUFX4_312/Y INVX1_438/A gnd OAI21X1_1536/C vdd OAI21X1
XDFFPOSX1_39 INVX1_339/A CLKBUF1_25/Y OAI21X1_363/Y gnd vdd DFFPOSX1
XOAI21X1_1557 INVX4_5/A BUFX4_197/Y OAI21X1_974/B gnd OAI21X1_1558/C vdd OAI21X1
XOAI21X1_1524 NAND2X1_79/Y BUFX4_429/Y OAI21X1_1524/C gnd OAI21X1_1524/Y vdd OAI21X1
XOAI21X1_1568 MUX2X1_4/B NAND2X1_85/Y OAI21X1_1568/C gnd DFFPOSX1_590/D vdd OAI21X1
XFILL_23_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XCLKBUF1_70 BUFX4_1/Y gnd CLKBUF1_70/Y vdd CLKBUF1
XCLKBUF1_92 BUFX4_5/Y gnd CLKBUF1_92/Y vdd CLKBUF1
XCLKBUF1_81 BUFX4_3/Y gnd CLKBUF1_81/Y vdd CLKBUF1
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_166 INVX1_166/A gnd INVX1_166/Y vdd INVX1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XINVX1_177 INVX1_177/A gnd INVX1_177/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd NOR3X1_13/B vdd INVX1
XCLKBUF1_103 BUFX4_7/Y gnd CLKBUF1_103/Y vdd CLKBUF1
XBUFX4_420 INVX8_3/Y gnd BUFX4_420/Y vdd BUFX4
XBUFX4_431 INVX8_23/Y gnd BUFX4_431/Y vdd BUFX4
XBUFX4_453 BUFX4_449/A gnd NOR2X1_84/B vdd BUFX4
XBUFX4_442 INVX8_2/Y gnd BUFX4_442/Y vdd BUFX4
XBUFX4_464 INVX8_10/Y gnd BUFX4_464/Y vdd BUFX4
XBUFX4_475 INVX8_15/Y gnd MUX2X1_66/B vdd BUFX4
XNOR2X1_513 INVX1_125/A AND2X2_22/A gnd OAI22X1_47/D vdd NOR2X1
XNOR2X1_524 BUFX4_51/Y OAI22X1_50/Y gnd NOR2X1_524/Y vdd NOR2X1
XNOR2X1_502 NOR2X1_502/A NOR2X1_502/B gnd NOR2X1_502/Y vdd NOR2X1
XNOR2X1_535 BUFX4_415/Y OAI22X1_53/Y gnd NOR2X1_535/Y vdd NOR2X1
XFILL_41_3 gnd vdd FILL
XNOR2X1_546 BUFX4_39/Y OAI22X1_58/Y gnd NOR2X1_546/Y vdd NOR2X1
XNOR2X1_557 BUFX4_48/Y OAI22X1_63/Y gnd NOR2X1_557/Y vdd NOR2X1
XNOR2X1_568 BUFX4_204/Y NOR2X1_568/B gnd NOR2X1_568/Y vdd NOR2X1
XFILL_27_1 gnd vdd FILL
XNOR2X1_579 NOR2X1_579/A BUFX4_275/Y gnd NOR2X1_579/Y vdd NOR2X1
XAOI21X1_104 MUX2X1_96/A NOR2X1_172/B NOR2X1_171/Y gnd AOI21X1_104/Y vdd AOI21X1
XAOI21X1_115 MUX2X1_96/A NOR2X1_188/B NOR2X1_188/Y gnd AOI21X1_115/Y vdd AOI21X1
XAOI21X1_137 MUX2X1_66/B MUX2X1_376/S NOR2X1_217/Y gnd AOI21X1_137/Y vdd AOI21X1
XAOI21X1_148 BUFX4_217/Y NOR2X1_234/Y NOR2X1_235/Y gnd AOI21X1_148/Y vdd AOI21X1
XAOI21X1_126 BUFX4_177/Y NOR2X1_707/B NOR2X1_203/Y gnd AOI21X1_126/Y vdd AOI21X1
XAOI21X1_159 BUFX4_469/Y NOR2X1_729/B NOR2X1_249/Y gnd AOI21X1_159/Y vdd AOI21X1
XOAI21X1_1332 BUFX4_121/Y BUFX4_396/Y INVX1_233/A gnd OAI21X1_1332/Y vdd OAI21X1
XOAI21X1_1310 BUFX4_61/Y BUFX4_55/Y AOI21X1_407/B gnd OAI21X1_1311/C vdd OAI21X1
XOAI21X1_1321 NAND2X1_40/Y BUFX4_317/Y OAI21X1_1321/C gnd OAI21X1_1321/Y vdd OAI21X1
XDFFPOSX1_922 NOR2X1_176/A CLKBUF1_83/Y AOI21X1_108/Y gnd vdd DFFPOSX1
XOAI21X1_1365 NAND2X1_53/Y BUFX4_322/Y OAI21X1_1365/C gnd DFFPOSX1_309/D vdd OAI21X1
XOAI21X1_1343 BUFX4_440/Y NAND2X1_51/Y OAI21X1_1343/C gnd OAI21X1_1343/Y vdd OAI21X1
XOAI21X1_1354 NOR2X1_77/B BUFX4_184/Y OAI21X1_947/B gnd OAI21X1_1355/C vdd OAI21X1
XDFFPOSX1_900 OAI21X1_846/A CLKBUF1_33/Y OAI21X1_219/Y gnd vdd DFFPOSX1
XDFFPOSX1_911 NOR2X1_170/A CLKBUF1_12/Y AOI21X1_103/Y gnd vdd DFFPOSX1
XDFFPOSX1_933 AND2X2_43/A CLKBUF1_39/Y OAI21X1_237/Y gnd vdd DFFPOSX1
XDFFPOSX1_955 NOR2X1_192/A CLKBUF1_37/Y AOI21X1_118/Y gnd vdd DFFPOSX1
XDFFPOSX1_966 OAI21X1_262/C CLKBUF1_49/Y OAI21X1_263/Y gnd vdd DFFPOSX1
XDFFPOSX1_944 OAI21X1_242/C CLKBUF1_9/Y OAI21X1_243/Y gnd vdd DFFPOSX1
XOAI21X1_1387 BUFX4_65/Y NAND2X1_58/Y OAI21X1_1386/Y gnd OAI21X1_1387/Y vdd OAI21X1
XOAI21X1_1376 BUFX4_385/Y BUFX4_128/Y OAI21X1_765/B gnd OAI21X1_1377/C vdd OAI21X1
XOAI21X1_1398 BUFX4_143/Y BUFX4_407/Y OAI21X1_582/B gnd OAI21X1_1398/Y vdd OAI21X1
XDFFPOSX1_988 NOR2X1_469/A CLKBUF1_74/Y OAI21X1_267/Y gnd vdd DFFPOSX1
XDFFPOSX1_999 AND2X2_25/A CLKBUF1_74/Y OAI21X1_281/Y gnd vdd DFFPOSX1
XDFFPOSX1_977 NOR2X1_208/A CLKBUF1_46/Y AOI21X1_130/Y gnd vdd DFFPOSX1
XFILL_46_1_1 gnd vdd FILL
XDFFPOSX1_218 INVX1_224/A CLKBUF1_24/Y MUX2X1_272/Y gnd vdd DFFPOSX1
XDFFPOSX1_207 AND2X2_28/B CLKBUF1_90/Y DFFPOSX1_207/D gnd vdd DFFPOSX1
XDFFPOSX1_229 NOR2X1_677/A CLKBUF1_62/Y AOI21X1_565/Y gnd vdd DFFPOSX1
XBUFX4_250 BUFX4_24/Y gnd BUFX4_250/Y vdd BUFX4
XBUFX4_261 BUFX4_22/Y gnd BUFX4_261/Y vdd BUFX4
XBUFX4_272 BUFX4_19/Y gnd BUFX4_272/Y vdd BUFX4
XFILL_37_1_1 gnd vdd FILL
XNOR2X1_310 NOR2X1_306/Y AND2X2_5/Y gnd INVX2_18/A vdd NOR2X1
XNOR2X1_343 INVX2_16/Y BUFX4_306/Y gnd XNOR2X1_7/B vdd NOR2X1
XNOR2X1_332 INVX1_204/Y INVX1_205/Y gnd OAI22X1_2/B vdd NOR2X1
XNOR2X1_321 INVX4_8/Y NOR2X1_321/B gnd NOR2X1_321/Y vdd NOR2X1
XBUFX4_294 INVX8_5/Y gnd BUFX4_294/Y vdd BUFX4
XBUFX4_283 BUFX4_20/Y gnd BUFX4_283/Y vdd BUFX4
XNOR2X1_365 BUFX4_81/Y NOR2X1_650/A gnd NOR2X1_365/Y vdd NOR2X1
XNOR2X1_354 AND2X2_18/B INVX4_9/A gnd INVX1_217/A vdd NOR2X1
XNOR2X1_376 NOR2X1_40/A BUFX4_339/Y gnd OAI22X1_6/A vdd NOR2X1
XNOR2X1_387 NOR2X1_386/Y NOR2X1_387/B gnd NOR2X1_387/Y vdd NOR2X1
XNOR2X1_398 INVX1_110/A BUFX4_224/Y gnd OAI22X1_15/D vdd NOR2X1
XOAI21X1_805 NOR3X1_14/Y OAI21X1_805/B NAND2X1_246/Y gnd NOR2X1_437/B vdd OAI21X1
XOAI21X1_849 INVX1_115/Y BUFX4_151/Y AOI21X1_373/Y gnd OAI21X1_850/C vdd OAI21X1
XOAI21X1_816 INVX1_33/A BUFX4_343/Y OAI21X1_816/C gnd OAI21X1_816/Y vdd OAI21X1
XFILL_20_0_1 gnd vdd FILL
XOAI21X1_827 INVX1_50/Y BUFX4_92/Y BUFX4_253/Y gnd OAI21X1_827/Y vdd OAI21X1
XOAI21X1_838 INVX1_334/Y AND2X2_23/A NAND2X1_253/Y gnd OAI21X1_838/Y vdd OAI21X1
XOAI21X1_1140 OAI22X1_62/Y BUFX4_41/Y BUFX4_201/Y gnd OAI22X1_63/B vdd OAI21X1
XMUX2X1_305 INVX1_230/Y MUX2X1_9/B MUX2X1_70/S gnd MUX2X1_305/Y vdd MUX2X1
XDFFPOSX1_730 NOR2X1_83/A CLKBUF1_27/Y AOI21X1_44/Y gnd vdd DFFPOSX1
XMUX2X1_327 INVX1_457/Y BUFX4_67/Y MUX2X1_84/S gnd MUX2X1_327/Y vdd MUX2X1
XDFFPOSX1_741 AND2X2_45/A CLKBUF1_92/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XOAI21X1_1173 BUFX4_336/Y INVX1_440/Y NAND2X1_340/Y gnd AOI21X1_493/B vdd OAI21X1
XMUX2X1_316 INVX1_297/Y MUX2X1_18/B MUX2X1_76/S gnd MUX2X1_316/Y vdd MUX2X1
XOAI21X1_1151 OAI21X1_1151/A BUFX4_411/Y BUFX4_202/Y gnd OAI22X1_65/C vdd OAI21X1
XOAI21X1_1162 BUFX4_328/Y INVX1_433/Y AOI21X1_488/Y gnd OAI21X1_1164/C vdd OAI21X1
XMUX2X1_338 BUFX4_68/Y INVX1_369/Y MUX2X1_96/S gnd MUX2X1_338/Y vdd MUX2X1
XOAI21X1_1184 OAI21X1_89/C BUFX4_265/Y BUFX4_84/Y gnd OAI22X1_68/B vdd OAI21X1
XDFFPOSX1_752 OAI21X1_111/C CLKBUF1_54/Y OAI21X1_112/Y gnd vdd DFFPOSX1
XMUX2X1_349 BUFX4_430/Y INVX1_308/Y MUX2X1_102/S gnd MUX2X1_349/Y vdd MUX2X1
XOAI21X1_1195 INVX1_72/A BUFX4_276/Y BUFX4_87/Y gnd OAI22X1_70/B vdd OAI21X1
XDFFPOSX1_763 NOR2X1_408/A CLKBUF1_46/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XDFFPOSX1_774 INVX1_72/A CLKBUF1_1/Y MUX2X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_785 NAND2X1_311/A CLKBUF1_99/Y OAI21X1_130/Y gnd vdd DFFPOSX1
XDFFPOSX1_796 INVX1_87/A CLKBUF1_55/Y MUX2X1_77/Y gnd vdd DFFPOSX1
XFILL_3_1_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_40_8_0 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XAOI21X1_490 BUFX4_414/Y MUX2X1_259/Y AOI21X1_489/Y gnd NOR2X1_568/B vdd AOI21X1
XNAND3X1_50 AOI22X1_5/Y AND2X2_11/A AOI22X1_6/Y gnd NAND3X1_50/Y vdd NAND3X1
XFILL_48_9_0 gnd vdd FILL
XNAND3X1_61 INVX4_9/A NAND3X1_60/Y NAND3X1_61/C gnd NAND3X1_61/Y vdd NAND3X1
XNAND3X1_72 BUFX4_36/Y NAND3X1_72/B NAND3X1_72/C gnd NAND3X1_72/Y vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_72 NOR2X1_72/A NOR2X1_70/Y gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_61 NOR2X1_61/A NOR2X1_60/Y gnd NOR2X1_61/Y vdd NOR2X1
XNOR2X1_50 NOR2X1_50/A MUX2X1_31/S gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_83 NOR2X1_83/A NOR2X1_83/B gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_94 NOR2X1_94/A NOR2X1_92/B gnd NOR2X1_94/Y vdd NOR2X1
XFILL_31_8_0 gnd vdd FILL
XNAND2X1_107 XNOR2X1_1/B INVX1_188/Y gnd INVX1_189/A vdd NAND2X1
XNAND2X1_118 BUFX2_3/A NOR3X1_7/Y gnd NOR2X1_349/B vdd NAND2X1
XNAND2X1_129 NAND2X1_129/A NOR2X1_321/B gnd OAI22X1_2/D vdd NAND2X1
XNAND2X1_5 NAND2X1_5/A NAND2X1_6/B gnd OAI21X1_2/C vdd NAND2X1
XFILL_39_9_0 gnd vdd FILL
XNOR2X1_140 BUFX4_127/Y BUFX4_454/Y gnd MUX2X1_89/S vdd NOR2X1
XMUX2X1_90 BUFX4_180/Y INVX1_103/Y MUX2X1_89/S gnd MUX2X1_90/Y vdd MUX2X1
XNOR2X1_151 MUX2X1_246/B MUX2X1_96/S gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_162 NOR2X1_162/A MUX2X1_340/S gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_184 INVX1_3/A INVX2_3/Y gnd INVX2_12/A vdd NOR2X1
XNOR2X1_173 BUFX4_138/Y NOR2X1_39/B gnd MUX2X1_102/S vdd NOR2X1
XNOR2X1_195 NOR2X1_619/A MUX2X1_364/S gnd NOR2X1_195/Y vdd NOR2X1
XFILL_22_8_0 gnd vdd FILL
XOAI21X1_602 BUFX4_369/Y NOR2X1_703/A BUFX4_151/Y gnd OAI21X1_602/Y vdd OAI21X1
XOAI21X1_613 BUFX4_154/Y OAI21X1_613/B BUFX4_361/Y gnd OAI21X1_613/Y vdd OAI21X1
XOAI21X1_624 AOI21X1_289/Y OAI21X1_624/B NAND3X1_72/Y gnd AOI21X1_292/B vdd OAI21X1
XOAI21X1_646 INVX1_278/Y BUFX4_241/Y NAND2X1_201/Y gnd MUX2X1_194/B vdd OAI21X1
XOAI21X1_635 INVX1_171/Y BUFX4_31/Y BUFX4_364/Y gnd AOI21X1_295/C vdd OAI21X1
XOAI21X1_657 BUFX4_336/Y NOR2X1_241/A BUFX4_155/Y gnd OAI22X1_9/C vdd OAI21X1
XOAI21X1_668 OAI21X1_248/C BUFX4_266/Y BUFX4_78/Y gnd OAI22X1_11/B vdd OAI21X1
XOAI21X1_679 OAI21X1_160/C BUFX4_84/Y AOI21X1_307/Y gnd OAI21X1_679/Y vdd OAI21X1
XMUX2X1_102 MUX2X1_96/A INVX1_115/Y MUX2X1_102/S gnd MUX2X1_102/Y vdd MUX2X1
XMUX2X1_113 INVX1_126/Y MUX2X1_66/B MUX2X1_360/S gnd MUX2X1_113/Y vdd MUX2X1
XMUX2X1_135 BUFX4_467/Y INVX1_148/Y MUX2X1_397/S gnd DFFPOSX1_5/D vdd MUX2X1
XMUX2X1_146 INVX1_159/Y BUFX4_213/Y MUX2X1_6/S gnd MUX2X1_146/Y vdd MUX2X1
XMUX2X1_124 MUX2X1_39/B INVX1_137/Y NOR2X1_232/Y gnd MUX2X1_124/Y vdd MUX2X1
XDFFPOSX1_582 INVX1_425/A CLKBUF1_72/Y MUX2X1_411/Y gnd vdd DFFPOSX1
XMUX2X1_179 MUX2X1_179/A MUX2X1_179/B BUFX4_93/Y gnd MUX2X1_179/Y vdd MUX2X1
XDFFPOSX1_571 NOR2X1_736/A CLKBUF1_53/Y AOI21X1_624/Y gnd vdd DFFPOSX1
XMUX2X1_157 INVX1_170/Y BUFX4_468/Y MUX2X1_14/S gnd MUX2X1_157/Y vdd MUX2X1
XDFFPOSX1_560 INVX1_326/A CLKBUF1_14/Y MUX2X1_399/Y gnd vdd DFFPOSX1
XMUX2X1_168 INVX1_182/Y BUFX4_371/Y MUX2X1_29/S gnd MUX2X1_168/Y vdd MUX2X1
XDFFPOSX1_593 NAND2X1_363/A CLKBUF1_47/Y DFFPOSX1_593/D gnd vdd DFFPOSX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XFILL_5_9_0 gnd vdd FILL
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XDFFPOSX1_5 INVX1_148/A CLKBUF1_97/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XFILL_13_8_0 gnd vdd FILL
XNOR2X1_8 NOR2X1_2/A INVX2_5/Y gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 MUX2X1_29/B NOR2X1_43/B NOR2X1_43/Y gnd AOI21X1_18/Y vdd AOI21X1
XAOI21X1_29 BUFX4_173/Y NOR2X1_60/Y NOR2X1_62/Y gnd AOI21X1_29/Y vdd AOI21X1
XOAI22X1_15 OAI22X1_15/A OAI22X1_15/B OAI22X1_15/C OAI22X1_15/D gnd OAI22X1_15/Y vdd
+ OAI22X1
XOAI22X1_37 OAI22X1_37/A OAI22X1_37/B OAI22X1_37/C BUFX4_39/Y gnd OAI22X1_37/Y vdd
+ OAI22X1
XOAI22X1_48 BUFX4_50/Y OAI22X1_48/B OAI22X1_48/C OAI22X1_48/D gnd MUX2X1_255/A vdd
+ OAI22X1
XOAI22X1_26 NOR2X1_448/Y OAI22X1_26/B OAI22X1_26/C NOR2X1_447/Y gnd OAI22X1_26/Y vdd
+ OAI22X1
XOAI22X1_59 NOR2X1_541/Y OAI22X1_59/B OAI22X1_59/C NOR2X1_546/Y gnd OAI22X1_59/Y vdd
+ OAI22X1
XOAI21X1_421 BUFX4_450/Y BUFX4_461/Y INVX1_281/A gnd OAI21X1_421/Y vdd OAI21X1
XOAI21X1_432 MUX2X1_77/B OAI21X1_64/B OAI21X1_431/Y gnd OAI21X1_432/Y vdd OAI21X1
XOAI21X1_410 OAI21X1_40/A MUX2X1_61/B OAI21X1_410/C gnd OAI21X1_410/Y vdd OAI21X1
XOAI21X1_443 AND2X2_3/Y AOI21X1_212/B traffic_Street_1[0] gnd NAND3X1_8/C vdd OAI21X1
XOAI21X1_465 AND2X2_5/Y NOR2X1_306/Y INVX4_7/Y gnd OAI21X1_465/Y vdd OAI21X1
XOAI21X1_454 AND2X2_5/Y NOR2X1_306/Y INVX4_7/A gnd NAND3X1_31/C vdd OAI21X1
XOAI21X1_498 AND2X2_3/Y NOR3X1_1/B OAI22X1_2/A gnd AND2X2_10/A vdd OAI21X1
XOAI21X1_476 NOR3X1_4/B MUX2X1_174/B BUFX2_3/A gnd OAI21X1_476/Y vdd OAI21X1
XOAI21X1_487 BUFX4_307/Y INVX4_7/A INVX2_18/A gnd OAI21X1_487/Y vdd OAI21X1
XDFFPOSX1_390 BUFX2_1/A CLKBUF1_59/Y AND2X2_19/Y gnd vdd DFFPOSX1
XFILL_8_0_1 gnd vdd FILL
XFILL_45_7_0 gnd vdd FILL
XFILL_36_7_0 gnd vdd FILL
XOAI21X1_70 NAND2X1_30/Y BUFX4_173/Y OAI21X1_69/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_81 BUFX4_448/Y BUFX4_43/Y NOR2X1_574/A gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_92 INVX1_48/Y NOR2X1_76/B NAND2X1_34/Y gnd OAI21X1_92/Y vdd OAI21X1
XFILL_2_7_0 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XOAI21X1_240 BUFX4_60/Y BUFX4_432/Y OAI21X1_667/B gnd OAI21X1_241/C vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_262 BUFX4_126/Y BUFX4_435/Y OAI21X1_262/C gnd OAI21X1_263/C vdd OAI21X1
XOAI21X1_251 NAND2X1_69/Y MUX2X1_96/A OAI21X1_250/Y gnd OAI21X1_251/Y vdd OAI21X1
XOAI21X1_273 BUFX4_216/Y NAND2X1_73/Y OAI21X1_272/Y gnd OAI21X1_273/Y vdd OAI21X1
XINVX1_315 INVX1_315/A gnd INVX1_315/Y vdd INVX1
XINVX1_304 INVX1_304/A gnd INVX1_304/Y vdd INVX1
XINVX1_326 INVX1_326/A gnd INVX1_326/Y vdd INVX1
XOAI21X1_295 NAND2X1_75/Y BUFX4_469/Y OAI21X1_294/Y gnd OAI21X1_295/Y vdd OAI21X1
XOAI21X1_284 BUFX4_192/Y BUFX4_163/Y AND2X2_47/A gnd OAI21X1_285/C vdd OAI21X1
XINVX1_337 INVX1_337/A gnd INVX1_337/Y vdd INVX1
XINVX1_348 INVX1_348/A gnd INVX1_348/Y vdd INVX1
XAND2X2_40 BUFX4_99/Y AND2X2_40/B gnd AND2X2_40/Y vdd AND2X2
XINVX1_359 INVX1_359/A gnd INVX1_359/Y vdd INVX1
XAND2X2_51 AND2X2_51/A AND2X2_51/B gnd AND2X2_51/Y vdd AND2X2
XNAND2X1_290 BUFX4_38/Y MUX2X1_237/Y gnd AOI22X1_26/A vdd NAND2X1
XNOR2X1_706 NOR2X1_706/A NOR2X1_703/B gnd NOR2X1_706/Y vdd NOR2X1
XFILL_18_7_0 gnd vdd FILL
XNOR2X1_717 NOR2X1_483/B NOR2X1_716/B gnd NOR2X1_717/Y vdd NOR2X1
XNOR2X1_739 NOR2X1_739/A NOR2X1_737/B gnd NOR2X1_739/Y vdd NOR2X1
XNOR2X1_728 NOR2X1_728/A NOR2X1_729/B gnd NOR2X1_728/Y vdd NOR2X1
XAOI21X1_308 BUFX4_412/Y MUX2X1_200/Y OAI21X1_687/Y gnd AOI21X1_308/Y vdd AOI21X1
XAOI21X1_319 BUFX4_250/Y AOI21X1_319/B OAI21X1_728/Y gnd OAI21X1_730/A vdd AOI21X1
XDFFPOSX1_18 INVX1_277/A CLKBUF1_14/Y OAI21X1_345/Y gnd vdd DFFPOSX1
XOAI21X1_1503 BUFX4_386/Y BUFX4_456/Y NOR2X1_566/A gnd OAI21X1_1504/C vdd OAI21X1
XOAI21X1_1514 NAND2X1_78/Y BUFX4_445/Y OAI21X1_1513/Y gnd DFFPOSX1_527/D vdd OAI21X1
XDFFPOSX1_29 INVX1_154/A CLKBUF1_19/Y MUX2X1_141/Y gnd vdd DFFPOSX1
XOAI21X1_1547 INVX4_3/A BUFX4_199/Y OAI21X1_793/B gnd OAI21X1_1548/C vdd OAI21X1
XOAI21X1_1536 NAND2X1_80/Y BUFX4_322/Y OAI21X1_1536/C gnd DFFPOSX1_546/D vdd OAI21X1
XOAI21X1_1525 BUFX4_389/Y BUFX4_311/Y INVX1_386/A gnd OAI21X1_1525/Y vdd OAI21X1
XOAI21X1_1569 MUX2X1_1/B NAND2X1_2/Y NAND2X1_361/Y gnd DFFPOSX1_591/D vdd OAI21X1
XOAI21X1_1558 NAND2X1_84/Y BUFX4_63/Y OAI21X1_1558/C gnd OAI21X1_1558/Y vdd OAI21X1
XCLKBUF1_60 BUFX4_4/Y gnd CLKBUF1_60/Y vdd CLKBUF1
XCLKBUF1_82 BUFX4_10/Y gnd CLKBUF1_82/Y vdd CLKBUF1
XCLKBUF1_93 BUFX4_6/Y gnd CLKBUF1_93/Y vdd CLKBUF1
XCLKBUF1_71 BUFX4_4/Y gnd CLKBUF1_71/Y vdd CLKBUF1
XFILL_42_5_0 gnd vdd FILL
XINVX1_101 INVX1_101/A gnd MUX2X1_88/B vdd INVX1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd MUX2X1_99/A vdd INVX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XBUFX4_421 INVX8_3/Y gnd BUFX4_421/Y vdd BUFX4
XBUFX4_410 address[2] gnd BUFX4_410/Y vdd BUFX4
XBUFX4_432 INVX8_23/Y gnd BUFX4_432/Y vdd BUFX4
XBUFX4_454 BUFX4_449/A gnd BUFX4_454/Y vdd BUFX4
XBUFX4_443 INVX8_2/Y gnd BUFX4_443/Y vdd BUFX4
XBUFX4_465 INVX8_15/Y gnd BUFX4_465/Y vdd BUFX4
XNOR2X1_514 NOR2X1_514/A BUFX4_340/Y gnd NOR2X1_514/Y vdd NOR2X1
XNOR2X1_503 NOR2X1_503/A BUFX4_285/Y gnd NOR2X1_503/Y vdd NOR2X1
XBUFX4_476 INVX8_16/Y gnd BUFX4_476/Y vdd BUFX4
XNOR2X1_525 NOR2X1_525/A BUFX4_338/Y gnd NOR2X1_525/Y vdd NOR2X1
XNOR2X1_558 OAI21X1_16/C BUFX4_231/Y gnd NOR2X1_558/Y vdd NOR2X1
XNOR2X1_547 BUFX4_356/Y INVX1_422/Y gnd NOR2X1_547/Y vdd NOR2X1
XNOR2X1_536 AND2X2_36/B NOR2X1_536/B gnd NOR2X1_536/Y vdd NOR2X1
XNOR2X1_569 NOR2X1_569/A BUFX4_330/Y gnd NOR2X1_569/Y vdd NOR2X1
XFILL_27_2 gnd vdd FILL
XFILL_33_5_0 gnd vdd FILL
XAOI21X1_105 BUFX4_466/Y NOR2X1_172/B NOR2X1_172/Y gnd AOI21X1_105/Y vdd AOI21X1
XAOI21X1_116 BUFX4_377/Y NOR2X1_188/B NOR2X1_189/Y gnd AOI21X1_116/Y vdd AOI21X1
XAOI21X1_149 BUFX4_180/Y NOR2X1_234/Y NOR2X1_236/Y gnd AOI21X1_149/Y vdd AOI21X1
XAOI21X1_138 MUX2X1_64/B NOR2X1_220/B NOR2X1_219/Y gnd AOI21X1_138/Y vdd AOI21X1
XAOI21X1_127 MUX2X1_66/B NOR2X1_707/B NOR2X1_204/Y gnd AOI21X1_127/Y vdd AOI21X1
XOAI21X1_1300 BUFX4_194/Y BUFX4_476/Y AND2X2_28/B gnd OAI21X1_1300/Y vdd OAI21X1
XOAI21X1_1322 INVX1_363/Y NOR2X1_97/B NAND2X1_354/Y gnd DFFPOSX1_372/D vdd OAI21X1
XOAI21X1_1311 BUFX4_68/Y NAND2X1_39/Y OAI21X1_1311/C gnd DFFPOSX1_184/D vdd OAI21X1
XDFFPOSX1_912 NOR2X1_171/A CLKBUF1_41/Y AOI21X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_923 INVX1_116/A CLKBUF1_29/Y MUX2X1_103/Y gnd vdd DFFPOSX1
XOAI21X1_1344 BUFX4_59/Y BUFX4_183/Y OAI21X1_759/B gnd OAI21X1_1345/C vdd OAI21X1
XOAI21X1_1355 NAND2X1_52/Y BUFX4_72/Y OAI21X1_1355/C gnd DFFPOSX1_320/D vdd OAI21X1
XOAI21X1_1333 NAND2X1_48/Y BUFX4_443/Y OAI21X1_1332/Y gnd OAI21X1_1333/Y vdd OAI21X1
XDFFPOSX1_901 OAI21X1_220/C CLKBUF1_12/Y OAI21X1_221/Y gnd vdd DFFPOSX1
XDFFPOSX1_956 NOR2X1_464/A CLKBUF1_82/Y AOI21X1_119/Y gnd vdd DFFPOSX1
XDFFPOSX1_945 OAI21X1_244/C CLKBUF1_82/Y OAI21X1_245/Y gnd vdd DFFPOSX1
XOAI21X1_1366 BUFX4_130/Y BUFX4_297/Y INVX1_245/A gnd OAI21X1_1367/C vdd OAI21X1
XOAI21X1_1388 BUFX4_133/Y BUFX4_129/Y DFFPOSX1_249/Q gnd OAI21X1_1389/C vdd OAI21X1
XOAI21X1_1377 NAND2X1_57/Y BUFX4_428/Y OAI21X1_1377/C gnd OAI21X1_1377/Y vdd OAI21X1
XOAI21X1_1399 BUFX4_445/Y NAND2X1_60/Y OAI21X1_1398/Y gnd OAI21X1_1399/Y vdd OAI21X1
XDFFPOSX1_934 OAI21X1_238/C CLKBUF1_12/Y OAI21X1_239/Y gnd vdd DFFPOSX1
XDFFPOSX1_967 INVX1_127/A CLKBUF1_37/Y MUX2X1_114/Y gnd vdd DFFPOSX1
XDFFPOSX1_978 NOR2X1_209/A CLKBUF1_102/Y AOI21X1_131/Y gnd vdd DFFPOSX1
XDFFPOSX1_989 INVX1_405/A CLKBUF1_44/Y OAI21X1_269/Y gnd vdd DFFPOSX1
XFILL_24_5_0 gnd vdd FILL
XFILL_7_6_0 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XDFFPOSX1_219 INVX1_303/A CLKBUF1_80/Y MUX2X1_273/Y gnd vdd DFFPOSX1
XDFFPOSX1_208 AND2X2_38/B CLKBUF1_48/Y OAI21X1_1303/Y gnd vdd DFFPOSX1
XBUFX4_240 BUFX4_17/Y gnd BUFX4_240/Y vdd BUFX4
XNOR2X1_300 AND2X2_3/B NOR2X1_300/B gnd INVX1_187/A vdd NOR2X1
XBUFX4_273 BUFX4_21/Y gnd BUFX4_273/Y vdd BUFX4
XBUFX4_262 BUFX4_21/Y gnd BUFX4_262/Y vdd BUFX4
XBUFX4_251 BUFX4_21/Y gnd BUFX4_251/Y vdd BUFX4
XNOR2X1_333 OAI22X1_2/A OAI22X1_2/B gnd XNOR2X1_4/B vdd NOR2X1
XNOR2X1_322 NOR2X1_321/Y INVX1_197/Y gnd INVX4_11/A vdd NOR2X1
XBUFX4_295 INVX8_5/Y gnd BUFX4_295/Y vdd BUFX4
XBUFX4_284 BUFX4_18/Y gnd BUFX4_284/Y vdd BUFX4
XNOR2X1_311 NAND3X1_32/Y NOR2X1_311/B gnd NOR2X1_311/Y vdd NOR2X1
XNOR2X1_366 INVX1_449/A BUFX4_151/Y gnd NOR2X1_366/Y vdd NOR2X1
XNOR2X1_344 OR2X2_2/A XNOR2X1_4/A gnd NOR2X1_344/Y vdd NOR2X1
XNOR2X1_377 BUFX4_149/Y NOR2X1_377/B gnd NOR2X1_377/Y vdd NOR2X1
XNOR2X1_355 NOR2X1_355/A INVX1_218/Y gnd NAND3X1_70/B vdd NOR2X1
XNOR2X1_388 INVX1_123/A BUFX4_265/Y gnd NOR2X1_388/Y vdd NOR2X1
XNOR2X1_399 NOR2X1_399/A BUFX4_344/Y gnd OAI22X1_15/A vdd NOR2X1
XOAI21X1_806 BUFX4_338/Y OAI21X1_45/C BUFX4_156/Y gnd OAI21X1_808/B vdd OAI21X1
XOAI21X1_817 NOR2X1_443/Y OAI21X1_815/Y OAI21X1_816/Y gnd MUX2X1_217/A vdd OAI21X1
XOAI21X1_828 INVX1_47/Y BUFX4_94/Y BUFX4_365/Y gnd OAI21X1_829/A vdd OAI21X1
XOAI21X1_839 BUFX4_358/Y OAI21X1_839/B BUFX4_158/Y gnd AOI21X1_368/C vdd OAI21X1
XOAI21X1_1130 BUFX4_223/Y DFFPOSX1_570/Q BUFX4_106/Y gnd OAI21X1_1130/Y vdd OAI21X1
XMUX2X1_339 AND2X2_5/B INVX1_242/Y NOR2X1_155/B gnd MUX2X1_339/Y vdd MUX2X1
XDFFPOSX1_731 INVX1_56/A CLKBUF1_97/Y MUX2X1_46/Y gnd vdd DFFPOSX1
XMUX2X1_328 INVX1_458/Y BUFX4_322/Y MUX2X1_84/S gnd MUX2X1_328/Y vdd MUX2X1
XOAI21X1_1141 BUFX4_326/Y NOR2X1_20/A BUFX4_159/Y gnd OAI21X1_1141/Y vdd OAI21X1
XMUX2X1_306 INVX1_294/Y MUX2X1_18/B MUX2X1_70/S gnd MUX2X1_306/Y vdd MUX2X1
XOAI21X1_1174 BUFX4_257/Y OAI21X1_1527/C BUFX4_80/Y gnd AOI21X1_492/C vdd OAI21X1
XOAI21X1_1152 OAI22X1_65/Y BUFX4_392/Y BUFX4_401/Y gnd OAI21X1_1176/B vdd OAI21X1
XDFFPOSX1_720 INVX1_50/A CLKBUF1_38/Y MUX2X1_40/Y gnd vdd DFFPOSX1
XMUX2X1_317 INVX1_342/Y BUFX4_69/Y MUX2X1_76/S gnd MUX2X1_317/Y vdd MUX2X1
XOAI21X1_1163 INVX1_435/Y BUFX4_247/Y BUFX4_74/Y gnd OAI21X1_1163/Y vdd OAI21X1
XDFFPOSX1_775 INVX1_73/A CLKBUF1_102/Y MUX2X1_63/Y gnd vdd DFFPOSX1
XOAI21X1_1185 OAI22X1_68/Y BUFX4_41/Y BUFX4_169/Y gnd OAI22X1_69/B vdd OAI21X1
XDFFPOSX1_742 OAI21X1_99/C CLKBUF1_48/Y OAI21X1_100/Y gnd vdd DFFPOSX1
XDFFPOSX1_764 INVX1_333/A CLKBUF1_13/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XDFFPOSX1_753 OAI21X1_113/C CLKBUF1_13/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XOAI21X1_1196 BUFX4_33/Y OAI22X1_70/Y NAND2X1_345/Y gnd OAI22X1_72/C vdd OAI21X1
XDFFPOSX1_797 INVX1_88/A CLKBUF1_6/Y MUX2X1_78/Y gnd vdd DFFPOSX1
XDFFPOSX1_786 OAI21X1_131/C CLKBUF1_58/Y OAI21X1_132/Y gnd vdd DFFPOSX1
XFILL_40_8_1 gnd vdd FILL
XAOI21X1_480 INVX1_31/Y BUFX4_326/Y BUFX4_159/Y gnd AOI21X1_480/Y vdd AOI21X1
XAOI21X1_491 BUFX4_253/Y NOR2X1_733/A BUFX4_78/Y gnd AOI21X1_491/Y vdd AOI21X1
XNAND3X1_40 INVX2_18/Y INVX4_10/Y NAND3X1_54/C gnd NAND3X1_40/Y vdd NAND3X1
XFILL_48_9_1 gnd vdd FILL
XNAND3X1_51 INVX4_9/Y NAND3X1_48/Y NAND3X1_51/C gnd NAND3X1_51/Y vdd NAND3X1
XNAND3X1_62 INVX4_10/Y NOR2X1_339/Y NAND3X1_54/C gnd NAND3X1_62/Y vdd NAND3X1
XNAND3X1_73 BUFX4_418/Y NAND3X1_73/B NAND3X1_73/C gnd NAND3X1_73/Y vdd NAND3X1
XFILL_47_4_0 gnd vdd FILL
XNOR2X1_62 NOR2X1_62/A NOR2X1_60/Y gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_51 INVX1_3/A INVX2_3/A gnd INVX2_9/A vdd NOR2X1
XNOR2X1_73 INVX2_9/Y INVX2_1/Y gnd INVX8_16/A vdd NOR2X1
XNOR2X1_40 NOR2X1_40/A NOR2X1_43/B gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_84 BUFX4_476/Y NOR2X1_84/B gnd NOR2X1_85/B vdd NOR2X1
XNOR2X1_95 NOR2X1_95/A NOR2X1_92/B gnd NOR2X1_95/Y vdd NOR2X1
XFILL_31_8_1 gnd vdd FILL
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_108 BUFX4_73/Y NOR2X1_304/Y gnd NOR2X1_351/B vdd NAND2X1
XNAND2X1_119 NAND3X1_25/Y OAI21X1_465/Y gnd NAND3X1_26/B vdd NAND2X1
XNAND2X1_6 NAND2X1_6/A NAND2X1_6/B gnd OAI21X1_3/C vdd NAND2X1
XFILL_39_9_1 gnd vdd FILL
XFILL_38_4_0 gnd vdd FILL
XNOR2X1_141 NOR2X1_598/A MUX2X1_89/S gnd NOR2X1_141/Y vdd NOR2X1
XMUX2X1_80 INVX1_93/Y BUFX4_214/Y MUX2X1_81/S gnd MUX2X1_80/Y vdd MUX2X1
XNOR2X1_130 INVX2_1/Y INVX2_11/Y gnd INVX8_20/A vdd NOR2X1
XNOR2X1_152 NOR2X1_585/A MUX2X1_96/S gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_174 NOR2X1_399/A MUX2X1_102/S gnd NOR2X1_174/Y vdd NOR2X1
XMUX2X1_91 MUX2X1_82/B MUX2X1_91/B MUX2X1_89/S gnd MUX2X1_91/Y vdd MUX2X1
XNOR2X1_185 INVX2_10/Y INVX2_12/Y gnd INVX8_23/A vdd NOR2X1
XNOR2X1_163 BUFX4_405/Y BUFX4_192/Y gnd NOR2X1_167/B vdd NOR2X1
XFILL_22_8_1 gnd vdd FILL
XNOR2X1_196 BUFX4_431/Y NOR2X1_96/B gnd NOR2X1_703/B vdd NOR2X1
XOAI21X1_614 BUFX4_154/Y NOR2X1_736/A BUFX4_285/Y gnd OAI21X1_614/Y vdd OAI21X1
XFILL_21_3_0 gnd vdd FILL
XOAI21X1_603 AND2X2_25/B OAI21X1_603/B BUFX4_99/Y gnd AOI21X1_278/C vdd OAI21X1
XOAI21X1_625 INVX1_272/Y BUFX4_291/Y NAND2X1_189/Y gnd MUX2X1_187/B vdd OAI21X1
XOAI21X1_636 INVX1_167/Y BUFX4_31/Y BUFX4_231/Y gnd AOI21X1_296/C vdd OAI21X1
XOAI21X1_647 INVX1_279/Y AND2X2_47/B NAND2X1_202/Y gnd MUX2X1_194/A vdd OAI21X1
XOAI21X1_669 OAI21X1_669/A BUFX4_35/Y OAI21X1_669/C gnd NOR2X1_390/B vdd OAI21X1
XOAI21X1_658 OAI21X1_320/C BUFX4_259/Y BUFX4_74/Y gnd OAI22X1_9/B vdd OAI21X1
XMUX2X1_114 INVX1_127/Y MUX2X1_97/B MUX2X1_366/S gnd MUX2X1_114/Y vdd MUX2X1
XMUX2X1_103 INVX1_116/Y MUX2X1_97/B MUX2X1_353/S gnd MUX2X1_103/Y vdd MUX2X1
XMUX2X1_125 BUFX4_180/Y INVX1_138/Y NOR2X1_232/Y gnd MUX2X1_125/Y vdd MUX2X1
XDFFPOSX1_550 NOR2X1_733/A CLKBUF1_97/Y AOI21X1_621/Y gnd vdd DFFPOSX1
XMUX2X1_147 INVX1_160/Y BUFX4_178/Y MUX2X1_6/S gnd MUX2X1_147/Y vdd MUX2X1
XMUX2X1_136 MUX2X1_39/B INVX1_149/Y MUX2X1_400/S gnd MUX2X1_136/Y vdd MUX2X1
XMUX2X1_169 INVX1_183/Y MUX2X1_66/B MUX2X1_29/S gnd MUX2X1_169/Y vdd MUX2X1
XDFFPOSX1_583 OAI21X1_616/B CLKBUF1_94/Y DFFPOSX1_583/D gnd vdd DFFPOSX1
XDFFPOSX1_561 INVX1_389/A CLKBUF1_25/Y MUX2X1_400/Y gnd vdd DFFPOSX1
XDFFPOSX1_572 NOR2X1_737/A CLKBUF1_73/Y AOI21X1_625/Y gnd vdd DFFPOSX1
XMUX2X1_158 INVX1_171/Y BUFX4_209/Y MUX2X1_18/S gnd MUX2X1_158/Y vdd MUX2X1
XDFFPOSX1_594 NAND2X1_3/A CLKBUF1_76/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XFILL_5_9_1 gnd vdd FILL
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XFILL_4_4_0 gnd vdd FILL
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XFILL_29_4_0 gnd vdd FILL
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XDFFPOSX1_6 DFFPOSX1_6/Q CLKBUF1_92/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XFILL_13_8_1 gnd vdd FILL
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 INVX2_4/A NOR2X1_9/B gnd INVX1_14/A vdd NOR2X1
XAOI21X1_19 MUX2X1_9/B NOR2X1_47/B NOR2X1_45/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI22X1_49 OAI22X1_49/A OAI22X1_49/B OAI22X1_49/C OAI22X1_49/D gnd OAI22X1_49/Y vdd
+ OAI22X1
XOAI22X1_16 NOR2X1_401/Y OAI22X1_16/B OAI22X1_16/C OAI22X1_16/D gnd OAI22X1_16/Y vdd
+ OAI22X1
XOAI22X1_27 NOR2X1_452/Y OAI22X1_27/B OAI22X1_27/C NOR2X1_451/Y gnd OAI22X1_27/Y vdd
+ OAI22X1
XOAI22X1_38 OAI22X1_38/A OAI22X1_38/B OAI22X1_38/C OAI22X1_38/D gnd OAI22X1_38/Y vdd
+ OAI22X1
XOAI21X1_400 NAND2X1_24/Y BUFX4_178/Y OAI21X1_399/Y gnd OAI21X1_400/Y vdd OAI21X1
XOAI21X1_422 OAI21X1_54/A BUFX4_209/Y OAI21X1_421/Y gnd OAI21X1_422/Y vdd OAI21X1
XOAI21X1_411 NOR2X1_39/A BUFX4_303/Y NOR2X1_608/A gnd OAI21X1_412/C vdd OAI21X1
XOAI21X1_444 AND2X2_1/Y NOR2X1_299/Y traffic_Street_1[3] gnd OR2X2_2/B vdd OAI21X1
XOAI21X1_433 BUFX4_190/Y BUFX4_462/Y AND2X2_46/A gnd OAI21X1_433/Y vdd OAI21X1
XOAI21X1_455 NOR3X1_4/C INVX2_15/Y traffic_Street_0[0] gnd NAND3X1_17/C vdd OAI21X1
XOAI21X1_466 NAND3X1_26/Y NOR3X1_6/A NOR2X1_309/Y gnd NOR3X1_9/C vdd OAI21X1
XOAI21X1_499 INVX1_205/A OR2X2_6/B NOR2X1_331/Y gnd AND2X2_10/B vdd OAI21X1
XOAI21X1_488 AND2X2_8/A INVX2_19/Y INVX1_201/Y gnd OAI21X1_488/Y vdd OAI21X1
XOAI21X1_477 INVX1_201/A NOR2X1_316/Y AOI22X1_9/C gnd OAI21X1_477/Y vdd OAI21X1
XDFFPOSX1_391 BUFX2_2/A CLKBUF1_59/Y NOR2X1_359/Y gnd vdd DFFPOSX1
XDFFPOSX1_380 INVX1_347/A CLKBUF1_65/Y MUX2X1_283/Y gnd vdd DFFPOSX1
XFILL_45_7_1 gnd vdd FILL
XFILL_44_2_0 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XFILL_36_7_1 gnd vdd FILL
XFILL_35_2_0 gnd vdd FILL
XOAI21X1_71 BUFX4_301/Y BUFX4_44/Y INVX1_398/A gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_60 MUX2X1_9/B OAI21X1_64/B OAI21X1_59/Y gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_82 NAND2X1_31/Y BUFX4_468/Y OAI21X1_81/Y gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_93 BUFX4_120/Y BUFX4_476/Y INVX1_289/A gnd OAI21X1_94/C vdd OAI21X1
XFILL_2_7_1 gnd vdd FILL
XFILL_27_7_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XOAI21X1_241 MUX2X1_97/B NAND2X1_68/Y OAI21X1_241/C gnd OAI21X1_241/Y vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XOAI21X1_230 BUFX4_383/Y BUFX4_141/Y INVX1_442/A gnd OAI21X1_231/C vdd OAI21X1
XOAI21X1_263 NAND2X1_70/Y MUX2X1_66/B OAI21X1_263/C gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_252 BUFX4_384/Y BUFX4_433/Y OAI21X1_252/C gnd OAI21X1_253/C vdd OAI21X1
XOAI21X1_274 BUFX4_135/Y BUFX4_160/Y OAI21X1_274/C gnd OAI21X1_274/Y vdd OAI21X1
XINVX1_316 INVX1_316/A gnd INVX1_316/Y vdd INVX1
XOAI21X1_296 BUFX4_386/Y BUFX4_458/Y OAI21X1_661/A gnd OAI21X1_296/Y vdd OAI21X1
XOAI21X1_285 MUX2X1_57/A NAND2X1_74/Y OAI21X1_285/C gnd OAI21X1_285/Y vdd OAI21X1
XINVX1_305 INVX1_305/A gnd INVX1_305/Y vdd INVX1
XAND2X2_30 BUFX4_232/Y AND2X2_30/B gnd AND2X2_30/Y vdd AND2X2
XINVX1_349 INVX1_349/A gnd INVX1_349/Y vdd INVX1
XINVX1_327 INVX1_327/A gnd INVX1_327/Y vdd INVX1
XINVX1_338 INVX1_338/A gnd INVX1_338/Y vdd INVX1
XAND2X2_41 AND2X2_41/A AND2X2_41/B gnd AND2X2_41/Y vdd AND2X2
XAND2X2_52 AND2X2_52/A AND2X2_52/B gnd AND2X2_52/Y vdd AND2X2
XFILL_9_3_0 gnd vdd FILL
XNAND2X1_280 NAND2X1_280/A NOR2X1_476/Y gnd NAND3X1_77/C vdd NAND2X1
XNAND2X1_291 BUFX4_222/Y NOR2X1_732/A gnd NAND2X1_291/Y vdd NAND2X1
XNOR2X1_707 NOR2X1_707/A NOR2X1_707/B gnd NOR2X1_707/Y vdd NOR2X1
XFILL_18_7_1 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XNOR2X1_718 NOR2X1_565/B NOR2X1_716/B gnd NOR2X1_718/Y vdd NOR2X1
XNOR2X1_729 NOR2X1_729/A NOR2X1_729/B gnd NOR2X1_729/Y vdd NOR2X1
XAOI21X1_309 BUFX4_414/Y MUX2X1_204/Y OAI21X1_697/Y gnd AOI21X1_310/C vdd AOI21X1
XOAI21X1_1504 NAND2X1_76/Y BUFX4_318/Y OAI21X1_1504/C gnd OAI21X1_1504/Y vdd OAI21X1
XOAI21X1_1537 BUFX4_194/Y BUFX4_312/Y NAND2X1_184/B gnd OAI21X1_1537/Y vdd OAI21X1
XOAI21X1_1548 NAND2X1_82/Y BUFX4_428/Y OAI21X1_1548/C gnd DFFPOSX1_568/D vdd OAI21X1
XDFFPOSX1_19 OAI21X1_876/A CLKBUF1_14/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XOAI21X1_1515 BUFX4_310/Y BUFX4_300/Y NAND2X1_244/A gnd OAI21X1_1516/C vdd OAI21X1
XOAI21X1_1526 NAND2X1_79/Y BUFX4_72/Y OAI21X1_1525/Y gnd OAI21X1_1526/Y vdd OAI21X1
XOAI21X1_1559 INVX4_5/A BUFX4_196/Y OAI21X1_1133/B gnd OAI21X1_1560/C vdd OAI21X1
XFILL_50_0_0 gnd vdd FILL
XCLKBUF1_50 BUFX4_10/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XCLKBUF1_61 BUFX4_9/Y gnd CLKBUF1_61/Y vdd CLKBUF1
XCLKBUF1_83 BUFX4_9/Y gnd CLKBUF1_83/Y vdd CLKBUF1
XCLKBUF1_72 BUFX4_1/Y gnd CLKBUF1_72/Y vdd CLKBUF1
XCLKBUF1_94 BUFX4_1/Y gnd CLKBUF1_94/Y vdd CLKBUF1
XFILL_41_0_0 gnd vdd FILL
XFILL_42_5_1 gnd vdd FILL
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_102 INVX1_102/A gnd MUX2X1_89/B vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XFILL_49_1_0 gnd vdd FILL
XBUFX4_400 address[5] gnd BUFX4_400/Y vdd BUFX4
XBUFX4_411 address[2] gnd BUFX4_411/Y vdd BUFX4
XBUFX4_422 INVX8_3/Y gnd BUFX4_422/Y vdd BUFX4
XBUFX4_433 INVX8_23/Y gnd BUFX4_433/Y vdd BUFX4
XBUFX4_455 INVX8_25/Y gnd BUFX4_455/Y vdd BUFX4
XBUFX4_444 INVX8_2/Y gnd BUFX4_444/Y vdd BUFX4
XBUFX4_466 INVX8_15/Y gnd BUFX4_466/Y vdd BUFX4
XNOR2X1_504 NOR2X1_503/Y NOR2X1_504/B gnd NOR2X1_504/Y vdd NOR2X1
XBUFX4_477 INVX8_16/Y gnd NOR2X1_74/B vdd BUFX4
XNOR2X1_515 NOR2X1_230/A BUFX4_155/Y gnd NOR2X1_515/Y vdd NOR2X1
XNOR2X1_526 BUFX4_37/Y NOR2X1_526/B gnd NOR2X1_526/Y vdd NOR2X1
XNOR2X1_559 INVX8_30/A NOR2X1_559/B gnd NOR2X1_559/Y vdd NOR2X1
XNOR2X1_548 address[6] OAI22X1_60/Y gnd NOR2X1_548/Y vdd NOR2X1
XNOR2X1_537 NOR2X1_692/A BUFX4_367/Y gnd NOR2X1_537/Y vdd NOR2X1
XFILL_27_3 gnd vdd FILL
XFILL_33_5_1 gnd vdd FILL
XAOI21X1_106 MUX2X1_97/B MUX2X1_102/S NOR2X1_174/Y gnd AOI21X1_106/Y vdd AOI21X1
XFILL_32_0_0 gnd vdd FILL
XAOI21X1_117 BUFX4_466/Y NOR2X1_188/B NOR2X1_190/Y gnd AOI21X1_117/Y vdd AOI21X1
XAOI21X1_139 BUFX4_465/Y NOR2X1_220/B NOR2X1_220/Y gnd AOI21X1_139/Y vdd AOI21X1
XAOI21X1_128 MUX2X1_59/B MUX2X1_369/S NOR2X1_206/Y gnd AOI21X1_128/Y vdd AOI21X1
XOAI21X1_1301 BUFX4_424/Y NAND2X1_37/Y OAI21X1_1300/Y gnd DFFPOSX1_207/D vdd OAI21X1
XOAI21X1_1323 BUFX4_57/Y BUFX4_398/Y NAND2X1_175/B gnd OAI21X1_1323/Y vdd OAI21X1
XOAI21X1_1312 BUFX4_58/Y BUFX4_52/Y DFFPOSX1_185/Q gnd OAI21X1_1312/Y vdd OAI21X1
XDFFPOSX1_924 INVX1_117/A CLKBUF1_27/Y MUX2X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_913 INVX1_114/A CLKBUF1_86/Y MUX2X1_101/Y gnd vdd DFFPOSX1
XDFFPOSX1_902 OAI21X1_222/C CLKBUF1_8/Y OAI21X1_223/Y gnd vdd DFFPOSX1
XOAI21X1_1345 BUFX4_428/Y NAND2X1_51/Y OAI21X1_1345/C gnd DFFPOSX1_323/D vdd OAI21X1
XOAI21X1_1356 NOR2X1_77/B BUFX4_183/Y OAI21X1_1119/B gnd OAI21X1_1356/Y vdd OAI21X1
XOAI21X1_1334 BUFX4_121/Y BUFX4_395/Y INVX1_298/A gnd OAI21X1_1334/Y vdd OAI21X1
XDFFPOSX1_946 OAI21X1_246/C CLKBUF1_49/Y OAI21X1_247/Y gnd vdd DFFPOSX1
XDFFPOSX1_957 NOR2X1_511/A CLKBUF1_82/Y AOI21X1_120/Y gnd vdd DFFPOSX1
XOAI21X1_1378 BUFX4_385/Y BUFX4_130/Y INVX1_351/A gnd OAI21X1_1379/C vdd OAI21X1
XOAI21X1_1367 NAND2X1_56/Y BUFX4_439/Y OAI21X1_1367/C gnd DFFPOSX1_286/D vdd OAI21X1
XOAI21X1_1389 BUFX4_321/Y NAND2X1_58/Y OAI21X1_1389/C gnd DFFPOSX1_249/D vdd OAI21X1
XDFFPOSX1_935 NOR2X1_181/A CLKBUF1_54/Y AOI21X1_111/Y gnd vdd DFFPOSX1
XDFFPOSX1_968 INVX1_128/A CLKBUF1_49/Y MUX2X1_115/Y gnd vdd DFFPOSX1
XDFFPOSX1_979 INVX1_133/A CLKBUF1_10/Y MUX2X1_120/Y gnd vdd DFFPOSX1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XINVX4_10 INVX4_10/A gnd INVX4_10/Y vdd INVX4
XFILL_7_6_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XDFFPOSX1_209 AOI21X1_467/B CLKBUF1_85/Y OAI21X1_1305/Y gnd vdd DFFPOSX1
XBUFX4_230 BUFX4_22/Y gnd BUFX4_230/Y vdd BUFX4
XNOR2X1_301 AND2X2_2/B AND2X2_2/A gnd NOR2X1_301/Y vdd NOR2X1
XBUFX4_263 BUFX4_24/Y gnd BUFX4_263/Y vdd BUFX4
XBUFX4_252 BUFX4_24/Y gnd BUFX4_252/Y vdd BUFX4
XBUFX4_241 BUFX4_20/Y gnd BUFX4_241/Y vdd BUFX4
XNOR2X1_334 NOR2X1_334/A NOR2X1_334/B gnd NOR2X1_334/Y vdd NOR2X1
XNOR2X1_312 INVX4_7/Y INVX4_6/Y gnd NOR2X1_312/Y vdd NOR2X1
XNOR2X1_323 INVX2_21/Y NOR3X1_10/Y gnd NOR2X1_341/B vdd NOR2X1
XBUFX4_296 INVX8_5/Y gnd NOR2X1_16/A vdd BUFX4
XBUFX4_274 BUFX4_24/Y gnd BUFX4_274/Y vdd BUFX4
XBUFX4_285 BUFX4_22/Y gnd BUFX4_285/Y vdd BUFX4
XNOR2X1_345 traffic_Street_1[3] NOR2X1_300/B gnd INVX2_26/A vdd NOR2X1
XNOR2X1_367 BUFX4_83/Y NOR2X1_367/B gnd NOR2X1_367/Y vdd NOR2X1
XNOR2X1_356 INVX1_192/Y BUFX4_307/Y gnd NOR2X1_356/Y vdd NOR2X1
XNOR2X1_389 NOR2X1_187/A BUFX4_344/Y gnd NOR2X1_389/Y vdd NOR2X1
XNOR2X1_378 BUFX4_34/Y MUX2X1_192/Y gnd NOR2X1_378/Y vdd NOR2X1
XOAI21X1_807 NOR2X1_41/A BUFX4_368/Y OAI21X1_807/C gnd OAI21X1_808/C vdd OAI21X1
XOAI21X1_818 OAI22X1_24/Y BUFX4_392/Y BUFX4_402/Y gnd OAI21X1_819/A vdd OAI21X1
XOAI21X1_829 OAI21X1_829/A NOR2X1_446/Y BUFX4_38/Y gnd OAI22X1_25/A vdd OAI21X1
XOAI21X1_1120 BUFX4_330/Y NOR2X1_669/A BUFX4_150/Y gnd OAI22X1_57/C vdd OAI21X1
XOAI21X1_1131 NOR2X1_549/Y OAI21X1_1130/Y OAI21X1_1131/C gnd NOR2X1_550/B vdd OAI21X1
XOAI21X1_1153 BUFX4_348/Y OAI21X1_1153/B BUFX4_147/Y gnd AOI21X1_483/C vdd OAI21X1
XDFFPOSX1_732 INVX1_57/A CLKBUF1_2/Y MUX2X1_47/Y gnd vdd DFFPOSX1
XOAI21X1_1142 INVX1_32/A BUFX4_332/Y AOI21X1_480/Y gnd OAI21X1_1142/Y vdd OAI21X1
XDFFPOSX1_710 OAI21X1_89/C CLKBUF1_24/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XMUX2X1_329 BUFX4_441/Y INVX1_244/Y MUX2X1_88/S gnd MUX2X1_329/Y vdd MUX2X1
XMUX2X1_307 INVX1_344/Y BUFX4_69/Y MUX2X1_70/S gnd MUX2X1_307/Y vdd MUX2X1
XDFFPOSX1_721 INVX1_51/A CLKBUF1_54/Y MUX2X1_41/Y gnd vdd DFFPOSX1
XMUX2X1_318 INVX1_453/Y BUFX4_316/Y MUX2X1_76/S gnd MUX2X1_318/Y vdd MUX2X1
XOAI21X1_1164 NOR2X1_563/Y OAI21X1_1163/Y OAI21X1_1164/C gnd MUX2X1_258/A vdd OAI21X1
XOAI21X1_1186 INVX1_48/Y BUFX4_266/Y BUFX4_148/Y gnd AOI21X1_495/C vdd OAI21X1
XDFFPOSX1_743 OAI21X1_101/C CLKBUF1_23/Y OAI21X1_102/Y gnd vdd DFFPOSX1
XOAI21X1_1175 MUX2X1_260/Y BUFX4_170/Y BUFX4_49/Y gnd OAI22X1_66/D vdd OAI21X1
XOAI21X1_1197 BUFX4_339/Y NOR2X1_109/A BUFX4_158/Y gnd OAI22X1_71/C vdd OAI21X1
XDFFPOSX1_765 NOR2X1_501/A CLKBUF1_15/Y OAI21X1_122/Y gnd vdd DFFPOSX1
XDFFPOSX1_754 OAI21X1_115/C CLKBUF1_58/Y OAI21X1_116/Y gnd vdd DFFPOSX1
XDFFPOSX1_776 INVX1_74/A CLKBUF1_68/Y MUX2X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_798 INVX1_89/A CLKBUF1_55/Y MUX2X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_787 INVX1_81/A CLKBUF1_77/Y MUX2X1_71/Y gnd vdd DFFPOSX1
XAOI21X1_470 BUFX4_276/Y AOI21X1_470/B AOI21X1_470/C gnd AOI21X1_470/Y vdd AOI21X1
XAOI21X1_492 BUFX4_258/Y INVX1_441/Y AOI21X1_492/C gnd AOI21X1_492/Y vdd AOI21X1
XAOI21X1_481 OAI21X1_41/C BUFX4_338/Y AND2X2_51/Y gnd AOI21X1_481/Y vdd AOI21X1
XNAND3X1_41 INVX4_7/Y NAND3X1_43/B NAND3X1_43/C gnd AOI22X1_5/D vdd NAND3X1
XNAND3X1_30 INVX4_6/A INVX1_190/Y NAND3X1_16/C gnd NAND3X1_30/Y vdd NAND3X1
XNAND3X1_52 INVX1_209/Y NAND3X1_58/A NAND3X1_58/C gnd NAND3X1_52/Y vdd NAND3X1
XNAND3X1_63 INVX4_9/A NAND3X1_62/Y NAND3X1_63/C gnd NAND3X1_63/Y vdd NAND3X1
XNAND3X1_74 BUFX4_153/Y NAND3X1_74/B NAND3X1_74/C gnd NAND3X1_74/Y vdd NAND3X1
XFILL_47_4_1 gnd vdd FILL
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B gnd NOR2X1_30/Y vdd NOR2X1
XNOR2X1_41 NOR2X1_41/A NOR2X1_43/B gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_63 NOR2X1_63/A NOR2X1_60/Y gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 INVX4_1/A INVX1_27/A gnd INVX2_10/A vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A NOR2X1_85/B gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_74 INVX4_2/A NOR2X1_74/B gnd NOR2X1_76/B vdd NOR2X1
XNOR2X1_96 BUFX4_52/Y NOR2X1_96/B gnd NOR2X1_97/B vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_109 traffic_Street_0[0] traffic_Street_0[1] gnd NAND3X1_14/B vdd NAND2X1
XNAND2X1_7 NAND2X1_7/A NAND2X1_6/B gnd NAND2X1_7/Y vdd NAND2X1
XFILL_38_4_1 gnd vdd FILL
XNOR2X1_131 BUFX4_131/Y BUFX4_57/Y gnd MUX2X1_88/S vdd NOR2X1
XNOR2X1_142 BUFX4_127/Y BUFX4_120/Y gnd MUX2X1_92/S vdd NOR2X1
XMUX2X1_81 INVX1_94/Y MUX2X1_49/A MUX2X1_81/S gnd MUX2X1_81/Y vdd MUX2X1
XNOR2X1_120 BUFX4_184/Y BUFX4_142/Y gnd MUX2X1_320/S vdd NOR2X1
XMUX2X1_70 INVX1_80/Y MUX2X1_58/A MUX2X1_70/S gnd MUX2X1_70/Y vdd MUX2X1
XNOR2X1_164 NOR2X1_164/A NOR2X1_167/B gnd AOI21X1_99/C vdd NOR2X1
XMUX2X1_92 BUFX4_217/Y MUX2X1_92/B MUX2X1_92/S gnd MUX2X1_92/Y vdd MUX2X1
XNOR2X1_153 BUFX4_405/Y BUFX4_56/Y gnd NOR2X1_155/B vdd NOR2X1
XNOR2X1_175 NOR2X1_175/A MUX2X1_102/S gnd NOR2X1_175/Y vdd NOR2X1
XNOR2X1_197 NOR2X1_197/A NOR2X1_703/B gnd NOR2X1_197/Y vdd NOR2X1
XNOR2X1_186 BUFX4_431/Y NOR2X1_39/B gnd NOR2X1_188/B vdd NOR2X1
XOAI21X1_615 AOI21X1_284/Y AOI21X1_285/Y BUFX4_41/Y gnd OAI21X1_615/Y vdd OAI21X1
XFILL_21_3_1 gnd vdd FILL
XOAI21X1_604 OAI21X1_604/A OAI21X1_604/B BUFX4_417/Y gnd OAI21X1_604/Y vdd OAI21X1
XOAI21X1_626 INVX1_28/Y BUFX4_220/Y NAND2X1_190/Y gnd MUX2X1_187/A vdd OAI21X1
XOAI21X1_637 INVX1_163/Y BUFX4_36/Y BUFX4_360/Y gnd OAI21X1_638/A vdd OAI21X1
XOAI21X1_648 INVX1_280/Y AND2X2_52/A OAI21X1_648/C gnd MUX2X1_195/B vdd OAI21X1
XOAI21X1_659 BUFX4_32/Y MUX2X1_198/Y NAND2X1_209/Y gnd OAI21X1_659/Y vdd OAI21X1
XMUX2X1_104 INVX1_117/Y MUX2X1_96/A MUX2X1_353/S gnd MUX2X1_104/Y vdd MUX2X1
XMUX2X1_115 INVX1_128/Y BUFX4_177/Y MUX2X1_366/S gnd MUX2X1_115/Y vdd MUX2X1
XMUX2X1_137 MUX2X1_86/B INVX1_150/Y MUX2X1_400/S gnd MUX2X1_137/Y vdd MUX2X1
XMUX2X1_126 BUFX4_381/Y INVX1_139/Y NOR2X1_232/Y gnd MUX2X1_126/Y vdd MUX2X1
XDFFPOSX1_540 INVX1_325/A CLKBUF1_60/Y MUX2X1_392/Y gnd vdd DFFPOSX1
XDFFPOSX1_573 NOR2X1_738/A CLKBUF1_53/Y AOI21X1_626/Y gnd vdd DFFPOSX1
XDFFPOSX1_562 NOR2X1_734/A CLKBUF1_19/Y AOI21X1_622/Y gnd vdd DFFPOSX1
XDFFPOSX1_551 INVX1_263/A CLKBUF1_90/Y MUX2X1_394/Y gnd vdd DFFPOSX1
XMUX2X1_148 INVX1_161/Y BUFX4_372/Y MUX2X1_6/S gnd MUX2X1_148/Y vdd MUX2X1
XMUX2X1_159 INVX1_172/Y BUFX4_178/Y MUX2X1_18/S gnd MUX2X1_159/Y vdd MUX2X1
XDFFPOSX1_584 OAI21X1_796/B CLKBUF1_35/Y OAI21X1_1556/Y gnd vdd DFFPOSX1
XDFFPOSX1_595 INVX1_4/A CLKBUF1_40/Y MUX2X1_1/Y gnd vdd DFFPOSX1
XINVX1_11 INVX1_11/A gnd MUX2X1_8/A vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XFILL_29_4_1 gnd vdd FILL
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XDFFPOSX1_7 DFFPOSX1_7/Q CLKBUF1_90/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XFILL_12_3_1 gnd vdd FILL
XOAI22X1_17 NOR2X1_404/Y OAI22X1_17/B OAI22X1_17/C OAI22X1_17/D gnd OAI22X1_17/Y vdd
+ OAI22X1
XOAI22X1_28 OAI22X1_28/A OAI22X1_28/B OAI22X1_28/C AND2X2_35/Y gnd OAI22X1_28/Y vdd
+ OAI22X1
XOAI22X1_39 OAI22X1_39/A OAI22X1_39/B OAI22X1_39/C OAI22X1_39/D gnd OAI22X1_39/Y vdd
+ OAI22X1
XOAI21X1_401 BUFX4_125/Y BUFX4_295/Y OAI21X1_401/C gnd OAI21X1_401/Y vdd OAI21X1
XOAI21X1_423 INVX4_4/A BUFX4_461/Y INVX1_338/A gnd OAI21X1_423/Y vdd OAI21X1
XOAI21X1_412 OAI21X1_40/A MUX2X1_58/A OAI21X1_412/C gnd OAI21X1_412/Y vdd OAI21X1
XOAI21X1_445 OR2X2_1/Y traffic_Street_1[0] AND2X2_3/A gnd OR2X2_2/A vdd OAI21X1
XOAI21X1_434 MUX2X1_61/B OAI21X1_64/B OAI21X1_433/Y gnd OAI21X1_434/Y vdd OAI21X1
XOAI21X1_456 AND2X2_4/Y NOR2X1_304/Y traffic_Street_0[3] gnd NAND3X1_18/C vdd OAI21X1
XOAI21X1_467 NOR3X1_9/C NOR3X1_3/Y INVX2_13/Y gnd OAI21X1_467/Y vdd OAI21X1
XOAI21X1_478 INVX4_7/Y INVX4_6/Y INVX2_14/Y gnd NAND2X1_129/A vdd OAI21X1
XOAI21X1_489 NOR2X1_326/Y OAI21X1_487/Y OAI21X1_488/Y gnd NAND3X1_64/C vdd OAI21X1
XDFFPOSX1_392 BUFX2_9/A CLKBUF1_59/Y AND2X2_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_370 NOR2X1_650/A CLKBUF1_61/Y AOI21X1_538/Y gnd vdd DFFPOSX1
XDFFPOSX1_381 INVX1_411/A CLKBUF1_29/Y MUX2X1_284/Y gnd vdd DFFPOSX1
XFILL_44_2_1 gnd vdd FILL
XOAI21X1_990 BUFX4_355/Y OAI21X1_47/C BUFX4_156/Y gnd OAI22X1_41/C vdd OAI21X1
XFILL_8_2 gnd vdd FILL
XFILL_35_2_1 gnd vdd FILL
XOAI21X1_72 NAND2X1_30/Y MUX2X1_82/B OAI21X1_71/Y gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_61 BUFX4_190/Y BUFX4_462/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_50 MUX2X1_29/B OAI21X1_48/B OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_83 BUFX4_124/Y BUFX4_46/Y OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_94 NAND2X1_36/Y BUFX4_217/Y OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XFILL_26_2_1 gnd vdd FILL
XOAI21X1_220 BUFX4_119/Y BUFX4_404/Y OAI21X1_220/C gnd OAI21X1_220/Y vdd OAI21X1
XOAI21X1_231 NAND2X1_64/Y BUFX4_466/Y OAI21X1_231/C gnd OAI21X1_231/Y vdd OAI21X1
XOAI21X1_242 BUFX4_60/Y BUFX4_432/Y OAI21X1_242/C gnd OAI21X1_242/Y vdd OAI21X1
XOAI21X1_253 NAND2X1_69/Y BUFX4_377/Y OAI21X1_253/C gnd OAI21X1_253/Y vdd OAI21X1
XOAI21X1_264 BUFX4_451/Y BUFX4_162/Y INVX1_284/A gnd OAI21X1_265/C vdd OAI21X1
XINVX1_317 INVX1_317/A gnd INVX1_317/Y vdd INVX1
XOAI21X1_297 NAND2X1_76/Y BUFX4_218/Y OAI21X1_296/Y gnd OAI21X1_297/Y vdd OAI21X1
XOAI21X1_275 MUX2X1_64/B NAND2X1_73/Y OAI21X1_274/Y gnd OAI21X1_275/Y vdd OAI21X1
XOAI21X1_286 BUFX4_192/Y BUFX4_163/Y NOR2X1_616/A gnd OAI21X1_286/Y vdd OAI21X1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XAND2X2_31 AND2X2_31/A BUFX4_97/Y gnd AND2X2_31/Y vdd AND2X2
XINVX1_339 INVX1_339/A gnd INVX1_339/Y vdd INVX1
XAND2X2_20 AND2X2_20/A INVX1_3/A gnd AND2X2_20/Y vdd AND2X2
XAND2X2_53 BUFX4_255/Y AND2X2_53/B gnd AND2X2_53/Y vdd AND2X2
XAND2X2_42 AND2X2_42/A BUFX4_91/Y gnd AND2X2_42/Y vdd AND2X2
XFILL_9_3_1 gnd vdd FILL
XNAND2X1_270 BUFX4_391/Y OAI22X1_36/Y gnd AOI21X1_391/A vdd NAND2X1
XNAND2X1_292 BUFX4_224/Y NAND2X1_292/B gnd NAND2X1_292/Y vdd NAND2X1
XNAND2X1_281 BUFX4_417/Y NAND2X1_281/B gnd NAND2X1_281/Y vdd NAND2X1
XNOR2X1_708 NOR2X1_428/B NOR2X1_707/B gnd NOR2X1_708/Y vdd NOR2X1
XFILL_17_2_1 gnd vdd FILL
XNOR2X1_719 NOR2X1_719/A NOR2X1_231/B gnd NOR2X1_719/Y vdd NOR2X1
XOAI21X1_1505 BUFX4_137/Y BUFX4_455/Y NAND2X1_187/B gnd OAI21X1_1506/C vdd OAI21X1
XOAI21X1_1538 BUFX4_440/Y NAND2X1_81/Y OAI21X1_1537/Y gnd DFFPOSX1_555/D vdd OAI21X1
XOAI21X1_1527 BUFX4_389/Y BUFX4_310/Y OAI21X1_1527/C gnd OAI21X1_1528/C vdd OAI21X1
XOAI21X1_1516 NAND2X1_78/Y BUFX4_429/Y OAI21X1_1516/C gnd DFFPOSX1_528/D vdd OAI21X1
XOAI21X1_1549 INVX4_3/A BUFX4_199/Y INVX1_390/A gnd OAI21X1_1549/Y vdd OAI21X1
XFILL_50_0_1 gnd vdd FILL
XFILL_20_9_0 gnd vdd FILL
XCLKBUF1_40 BUFX4_7/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XCLKBUF1_51 BUFX4_3/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XCLKBUF1_62 BUFX4_6/Y gnd CLKBUF1_62/Y vdd CLKBUF1
XCLKBUF1_84 BUFX4_7/Y gnd CLKBUF1_84/Y vdd CLKBUF1
XCLKBUF1_73 BUFX4_2/Y gnd CLKBUF1_73/Y vdd CLKBUF1
XCLKBUF1_95 BUFX4_10/Y gnd CLKBUF1_95/Y vdd CLKBUF1
XFILL_41_0_1 gnd vdd FILL
XFILL_11_9_0 gnd vdd FILL
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XFILL_49_1_1 gnd vdd FILL
XBUFX4_401 address[5] gnd BUFX4_401/Y vdd BUFX4
XBUFX4_412 address[2] gnd BUFX4_412/Y vdd BUFX4
XBUFX4_434 INVX8_23/Y gnd BUFX4_434/Y vdd BUFX4
XBUFX4_423 INVX8_3/Y gnd MUX2X1_6/B vdd BUFX4
XBUFX4_456 INVX8_25/Y gnd BUFX4_456/Y vdd BUFX4
XBUFX4_445 INVX8_2/Y gnd BUFX4_445/Y vdd BUFX4
XBUFX4_467 INVX8_15/Y gnd BUFX4_467/Y vdd BUFX4
XNOR2X1_505 NOR2X1_505/A BUFX4_288/Y gnd NOR2X1_505/Y vdd NOR2X1
XBUFX4_478 INVX8_16/Y gnd BUFX4_478/Y vdd BUFX4
XNOR2X1_516 NOR2X1_516/A BUFX4_81/Y gnd NOR2X1_516/Y vdd NOR2X1
XNOR2X1_549 NOR2X1_739/A BUFX4_363/Y gnd NOR2X1_549/Y vdd NOR2X1
XNOR2X1_538 BUFX4_393/Y NOR2X1_538/B gnd OAI22X1_60/D vdd NOR2X1
XNOR2X1_527 BUFX4_272/Y INVX1_448/A gnd NOR2X1_527/Y vdd NOR2X1
XFILL_32_0_1 gnd vdd FILL
XAOI21X1_118 MUX2X1_97/B MUX2X1_364/S NOR2X1_192/Y gnd AOI21X1_118/Y vdd AOI21X1
XAOI21X1_129 BUFX4_177/Y MUX2X1_369/S NOR2X1_207/Y gnd AOI21X1_129/Y vdd AOI21X1
XAOI21X1_107 MUX2X1_44/A MUX2X1_102/S NOR2X1_175/Y gnd AOI21X1_107/Y vdd AOI21X1
XOAI21X1_1302 BUFX4_193/Y BUFX4_478/Y AND2X2_38/B gnd OAI21X1_1302/Y vdd OAI21X1
XOAI21X1_1313 BUFX4_316/Y NAND2X1_39/Y OAI21X1_1312/Y gnd OAI21X1_1313/Y vdd OAI21X1
XDFFPOSX1_914 NOR2X1_172/A CLKBUF1_37/Y AOI21X1_105/Y gnd vdd DFFPOSX1
XDFFPOSX1_903 NOR2X1_164/A CLKBUF1_101/Y AOI21X1_99/Y gnd vdd DFFPOSX1
XOAI21X1_1324 MUX2X1_9/B NAND2X1_44/Y OAI21X1_1323/Y gnd OAI21X1_1324/Y vdd OAI21X1
XOAI21X1_1346 BUFX4_56/Y BUFX4_184/Y NAND2X1_282/B gnd OAI21X1_1347/C vdd OAI21X1
XOAI21X1_1335 NAND2X1_48/Y MUX2X1_18/B OAI21X1_1334/Y gnd OAI21X1_1335/Y vdd OAI21X1
XDFFPOSX1_936 INVX1_122/A CLKBUF1_101/Y MUX2X1_109/Y gnd vdd DFFPOSX1
XDFFPOSX1_947 OAI21X1_248/C CLKBUF1_9/Y OAI21X1_249/Y gnd vdd DFFPOSX1
XOAI21X1_1379 NAND2X1_57/Y BUFX4_65/Y OAI21X1_1379/C gnd DFFPOSX1_272/D vdd OAI21X1
XOAI21X1_1368 BUFX4_128/Y BUFX4_297/Y NOR2X1_424/B gnd OAI21X1_1369/C vdd OAI21X1
XOAI21X1_1357 NAND2X1_52/Y BUFX4_318/Y OAI21X1_1356/Y gnd DFFPOSX1_321/D vdd OAI21X1
XDFFPOSX1_925 INVX1_118/A CLKBUF1_54/Y MUX2X1_105/Y gnd vdd DFFPOSX1
XDFFPOSX1_958 NOR2X1_619/A CLKBUF1_9/Y AOI21X1_121/Y gnd vdd DFFPOSX1
XDFFPOSX1_969 INVX1_129/A CLKBUF1_9/Y MUX2X1_116/Y gnd vdd DFFPOSX1
XFILL_23_0_1 gnd vdd FILL
XINVX4_11 INVX4_11/A gnd INVX4_11/Y vdd INVX4
XFILL_6_1_1 gnd vdd FILL
XFILL_43_8_0 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XBUFX4_220 BUFX4_20/Y gnd BUFX4_220/Y vdd BUFX4
XBUFX4_242 BUFX4_20/Y gnd BUFX4_242/Y vdd BUFX4
XBUFX4_264 BUFX4_18/Y gnd AND2X2_23/A vdd BUFX4
XBUFX4_231 BUFX4_17/Y gnd BUFX4_231/Y vdd BUFX4
XBUFX4_253 BUFX4_19/Y gnd BUFX4_253/Y vdd BUFX4
XNOR2X1_324 INVX1_203/A OAI22X1_2/C gnd INVX4_12/A vdd NOR2X1
XNOR2X1_313 INVX4_7/A INVX4_6/A gnd NOR2X1_314/A vdd NOR2X1
XNOR2X1_302 NOR2X1_299/Y AND2X2_1/Y gnd AOI22X1_9/D vdd NOR2X1
XBUFX4_297 BUFX4_302/A gnd BUFX4_297/Y vdd BUFX4
XBUFX4_286 BUFX4_19/Y gnd AND2X2_36/B vdd BUFX4
XBUFX4_275 BUFX4_19/Y gnd BUFX4_275/Y vdd BUFX4
XNOR2X1_368 BUFX4_337/Y INVX1_235/Y gnd NOR2X1_368/Y vdd NOR2X1
XNOR2X1_346 NOR2X1_344/Y XNOR2X1_6/Y gnd NAND3X1_66/C vdd NOR2X1
XNOR2X1_335 NOR3X1_10/Y NAND3X1_65/C gnd NOR2X1_335/Y vdd NOR2X1
XNOR2X1_357 police_Interrupt NOR2X1_357/B gnd AND2X2_17/A vdd NOR2X1
XFILL_34_8_0 gnd vdd FILL
XFILL_25_1 gnd vdd FILL
XNOR2X1_379 NOR2X1_379/A BUFX4_252/Y gnd OAI22X1_7/D vdd NOR2X1
XOAI21X1_819 OAI21X1_819/A NOR2X1_437/Y OAI21X1_819/C gnd OAI21X1_820/A vdd OAI21X1
XOAI21X1_808 NOR2X1_438/Y OAI21X1_808/B OAI21X1_808/C gnd NOR2X1_439/B vdd OAI21X1
XOAI21X1_1121 BUFX4_291/Y INVX1_454/A BUFX4_102/Y gnd OAI22X1_57/B vdd OAI21X1
XOAI21X1_1110 BUFX4_282/Y INVX1_459/A AOI21X1_474/Y gnd OAI21X1_1110/Y vdd OAI21X1
XDFFPOSX1_722 INVX1_52/A CLKBUF1_41/Y MUX2X1_42/Y gnd vdd DFFPOSX1
XOAI21X1_1132 BUFX4_225/Y INVX1_461/A AOI21X1_479/Y gnd OAI21X1_1132/Y vdd OAI21X1
XOAI21X1_1143 NOR2X1_558/Y OAI21X1_1141/Y OAI21X1_1142/Y gnd NOR2X1_559/B vdd OAI21X1
XDFFPOSX1_711 NOR2X1_71/A CLKBUF1_80/Y AOI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_700 OAI21X1_77/C CLKBUF1_24/Y OAI21X1_78/Y gnd vdd DFFPOSX1
XMUX2X1_319 BUFX4_440/Y INVX1_249/Y MUX2X1_320/S gnd MUX2X1_319/Y vdd MUX2X1
XOAI21X1_1165 MUX2X1_258/Y BUFX4_170/Y BUFX4_393/Y gnd OAI22X1_66/A vdd OAI21X1
XMUX2X1_308 INVX1_417/Y BUFX4_316/Y MUX2X1_70/S gnd MUX2X1_308/Y vdd MUX2X1
XOAI21X1_1154 AND2X2_22/A OAI21X1_1452/C BUFX4_114/Y gnd AOI21X1_484/C vdd OAI21X1
XDFFPOSX1_755 INVX1_65/A CLKBUF1_1/Y MUX2X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_733 INVX1_58/A CLKBUF1_90/Y MUX2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_744 AOI21X1_362/A CLKBUF1_85/Y OAI21X1_104/Y gnd vdd DFFPOSX1
XOAI21X1_1176 NOR2X1_557/Y OAI21X1_1176/B NAND2X1_341/Y gnd OAI21X1_1177/A vdd OAI21X1
XOAI21X1_1198 OAI21X1_140/C BUFX4_278/Y BUFX4_88/Y gnd OAI22X1_71/B vdd OAI21X1
XDFFPOSX1_766 NOR2X1_579/A CLKBUF1_46/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XOAI21X1_1187 INVX1_55/Y BUFX4_268/Y BUFX4_85/Y gnd AOI21X1_496/C vdd OAI21X1
XDFFPOSX1_788 INVX1_82/A CLKBUF1_20/Y MUX2X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_777 INVX1_75/A CLKBUF1_20/Y MUX2X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_799 NOR2X1_107/A CLKBUF1_88/Y AOI21X1_59/Y gnd vdd DFFPOSX1
XFILL_0_8_0 gnd vdd FILL
XFILL_25_8_0 gnd vdd FILL
XAOI21X1_460 NOR2X1_248/A BUFX4_261/Y AOI21X1_460/C gnd NOR2X1_520/B vdd AOI21X1
XAOI21X1_482 INVX1_37/Y BUFX4_368/Y BUFX4_156/Y gnd AOI21X1_482/Y vdd AOI21X1
XAOI21X1_493 BUFX4_155/Y AOI21X1_493/B AOI21X1_492/Y gnd MUX2X1_260/A vdd AOI21X1
XAOI21X1_471 BUFX4_278/Y NOR2X1_654/A AOI21X1_471/C gnd AOI21X1_471/Y vdd AOI21X1
XFILL_8_9_0 gnd vdd FILL
XNAND3X1_20 NOR2X1_351/B AND2X2_6/A NAND3X1_20/C gnd NAND3X1_20/Y vdd NAND3X1
XNAND3X1_31 BUFX2_3/A NAND3X1_17/Y NAND3X1_31/C gnd NAND3X1_31/Y vdd NAND3X1
XNAND3X1_53 INVX4_9/Y NAND3X1_52/Y NAND3X1_53/C gnd NAND3X1_53/Y vdd NAND3X1
XNAND3X1_42 INVX4_11/A NAND3X1_43/B NAND3X1_43/C gnd XOR2X1_3/A vdd NAND3X1
XNAND3X1_64 XOR2X1_3/Y NAND3X1_64/B NAND3X1_64/C gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_75 BUFX4_48/Y NAND3X1_75/B NAND3X1_75/C gnd NAND3X1_75/Y vdd NAND3X1
XNOR2X1_20 NOR2X1_20/A NOR2X1_16/Y gnd AOI21X1_4/C vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A NOR2X1_60/Y gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_31 NOR2X1_31/A NOR2X1_30/B gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_53 INVX2_9/Y INVX2_10/Y gnd INVX8_12/A vdd NOR2X1
XNOR2X1_42 NOR2X1_42/A NOR2X1_43/B gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_86 BUFX4_479/Y BUFX4_137/Y gnd MUX2X1_50/S vdd NOR2X1
XFILL_16_8_0 gnd vdd FILL
XNOR2X1_75 NOR2X1_75/A NOR2X1_76/B gnd NOR2X1_75/Y vdd NOR2X1
XNAND2X1_8 NAND2X1_8/A NAND2X1_6/B gnd NAND2X1_8/Y vdd NAND2X1
XNOR2X1_132 NOR2X1_132/A MUX2X1_88/S gnd NOR2X1_132/Y vdd NOR2X1
XNOR2X1_121 NOR2X1_121/A MUX2X1_320/S gnd AOI21X1_68/C vdd NOR2X1
XNOR2X1_110 BUFX4_398/Y BUFX4_190/Y gnd AOI21X1_62/B vdd NOR2X1
XMUX2X1_60 INVX1_70/Y MUX2X1_64/B MUX2X1_59/S gnd MUX2X1_60/Y vdd MUX2X1
XMUX2X1_71 INVX1_81/Y MUX2X1_71/B MUX2X1_71/S gnd MUX2X1_71/Y vdd MUX2X1
XNOR2X1_154 NOR2X1_154/A NOR2X1_155/B gnd AOI21X1_91/C vdd NOR2X1
XNOR2X1_143 NOR2X1_143/A MUX2X1_92/S gnd NOR2X1_143/Y vdd NOR2X1
XMUX2X1_82 INVX1_95/Y MUX2X1_82/B MUX2X1_81/S gnd MUX2X1_82/Y vdd MUX2X1
XMUX2X1_93 MUX2X1_82/B INVX1_106/Y MUX2X1_92/S gnd MUX2X1_93/Y vdd MUX2X1
XNOR2X1_165 NOR2X1_165/A NOR2X1_167/B gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_176 NOR2X1_176/A MUX2X1_102/S gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_198 NOR2X1_198/A NOR2X1_703/B gnd NOR2X1_198/Y vdd NOR2X1
XNOR2X1_187 NOR2X1_187/A NOR2X1_188/B gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_605 INVX1_261/Y BUFX4_102/Y OAI21X1_605/C gnd OAI21X1_605/Y vdd OAI21X1
XOAI21X1_627 INVX1_273/Y BUFX4_222/Y NAND2X1_192/Y gnd MUX2X1_188/B vdd OAI21X1
XOAI21X1_616 BUFX4_154/Y OAI21X1_616/B BUFX4_351/Y gnd AOI21X1_286/C vdd OAI21X1
XOAI21X1_638 OAI21X1_638/A AND2X2_24/Y BUFX4_149/Y gnd OAI21X1_639/A vdd OAI21X1
XOAI21X1_649 INVX1_175/Y BUFX4_247/Y NAND2X1_204/Y gnd MUX2X1_195/A vdd OAI21X1
XMUX2X1_105 INVX1_118/Y MUX2X1_44/A MUX2X1_353/S gnd MUX2X1_105/Y vdd MUX2X1
XMUX2X1_116 INVX1_129/Y BUFX4_377/Y MUX2X1_366/S gnd MUX2X1_116/Y vdd MUX2X1
XMUX2X1_127 BUFX4_467/Y INVX1_140/Y NOR2X1_232/Y gnd MUX2X1_127/Y vdd MUX2X1
XMUX2X1_138 INVX1_151/Y MUX2X1_39/B MUX2X1_406/S gnd MUX2X1_138/Y vdd MUX2X1
XDFFPOSX1_530 NAND2X1_340/A CLKBUF1_64/Y DFFPOSX1_530/D gnd vdd DFFPOSX1
XDFFPOSX1_541 NOR2X1_729/A CLKBUF1_89/Y AOI21X1_617/Y gnd vdd DFFPOSX1
XDFFPOSX1_574 NOR2X1_739/A CLKBUF1_19/Y AOI21X1_627/Y gnd vdd DFFPOSX1
XDFFPOSX1_563 INVX1_269/A CLKBUF1_53/Y MUX2X1_401/Y gnd vdd DFFPOSX1
XMUX2X1_149 INVX1_162/Y BUFX4_470/Y MUX2X1_6/S gnd MUX2X1_149/Y vdd MUX2X1
XDFFPOSX1_552 INVX1_323/A CLKBUF1_17/Y MUX2X1_395/Y gnd vdd DFFPOSX1
XDFFPOSX1_596 INVX1_5/A CLKBUF1_98/Y MUX2X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_585 OAI21X1_974/B CLKBUF1_11/Y OAI21X1_1558/Y gnd vdd DFFPOSX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XDFFPOSX1_8 AND2X2_49/A CLKBUF1_90/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XFILL_40_6_0 gnd vdd FILL
XAOI21X1_290 NAND2X1_5/A BUFX4_343/Y BUFX4_159/Y gnd OAI21X1_622/C vdd AOI21X1
XFILL_48_7_0 gnd vdd FILL
XFILL_31_6_0 gnd vdd FILL
XFILL_39_7_0 gnd vdd FILL
XOAI22X1_29 NOR2X1_454/Y OAI22X1_29/B OAI22X1_29/C NOR2X1_453/Y gnd OAI22X1_29/Y vdd
+ OAI22X1
XOAI22X1_18 OAI22X1_18/A OAI22X1_18/B OAI22X1_18/C OAI22X1_18/D gnd OAI22X1_18/Y vdd
+ OAI22X1
XFILL_22_6_0 gnd vdd FILL
XOAI21X1_402 NAND2X1_24/Y BUFX4_375/Y OAI21X1_401/Y gnd OAI21X1_402/Y vdd OAI21X1
XOAI21X1_413 BUFX4_62/Y BUFX4_460/Y OAI21X1_413/C gnd OAI21X1_414/C vdd OAI21X1
XOAI21X1_446 AOI22X1_9/D AND2X2_3/B OR2X2_2/A gnd NAND3X1_12/B vdd OAI21X1
XOAI21X1_435 BUFX4_190/Y BUFX4_462/Y NOR2X1_611/A gnd OAI21X1_435/Y vdd OAI21X1
XOAI21X1_424 OAI21X1_54/A MUX2X1_77/B OAI21X1_423/Y gnd OAI21X1_424/Y vdd OAI21X1
XOAI21X1_457 OR2X2_3/Y traffic_Street_0[0] AND2X2_6/A gnd INVX1_214/A vdd OAI21X1
XOAI21X1_468 AOI22X1_1/Y INVX1_187/A INVX4_6/Y gnd OAI21X1_468/Y vdd OAI21X1
XOAI21X1_479 INVX2_18/Y INVX2_19/A INVX1_196/Y gnd XOR2X1_1/A vdd OAI21X1
XDFFPOSX1_382 NOR2X1_632/A CLKBUF1_80/Y AOI21X1_520/Y gnd vdd DFFPOSX1
XDFFPOSX1_360 INVX1_344/A CLKBUF1_98/Y MUX2X1_307/Y gnd vdd DFFPOSX1
XDFFPOSX1_371 NOR2X1_412/B CLKBUF1_15/Y AOI21X1_539/Y gnd vdd DFFPOSX1
XDFFPOSX1_393 BUFX2_10/A CLKBUF1_59/Y NOR2X1_358/Y gnd vdd DFFPOSX1
XFILL_5_7_0 gnd vdd FILL
XFILL_13_6_0 gnd vdd FILL
XOAI21X1_980 INVX1_6/Y BUFX4_347/Y OAI21X1_980/C gnd NAND3X1_78/C vdd OAI21X1
XOAI21X1_991 INVX1_36/A AND2X2_52/A BUFX4_88/Y gnd OAI22X1_41/B vdd OAI21X1
XOAI21X1_51 BUFX4_450/Y BUFX4_462/Y INVX1_275/A gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_62 MUX2X1_6/B OAI21X1_64/B OAI21X1_61/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_40 OAI21X1_40/A BUFX4_70/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_84 NAND2X1_32/Y BUFX4_213/Y OAI21X1_83/Y gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_73 BUFX4_301/Y BUFX4_44/Y OAI21X1_73/C gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_95 INVX4_5/A BUFX4_479/Y AND2X2_31/A gnd OAI21X1_96/C vdd OAI21X1
XOAI21X1_210 BUFX4_451/Y BUFX4_405/Y NOR2X1_447/A gnd OAI21X1_210/Y vdd OAI21X1
XOAI21X1_221 NAND2X1_62/Y MUX2X1_57/A OAI21X1_220/Y gnd OAI21X1_221/Y vdd OAI21X1
XOAI21X1_243 BUFX4_177/Y NAND2X1_68/Y OAI21X1_242/Y gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_254 BUFX4_384/Y BUFX4_434/Y OAI21X1_254/C gnd OAI21X1_255/C vdd OAI21X1
XOAI21X1_265 NAND2X1_72/Y BUFX4_216/Y OAI21X1_265/C gnd OAI21X1_265/Y vdd OAI21X1
XOAI21X1_232 BUFX4_123/Y BUFX4_139/Y INVX1_288/A gnd OAI21X1_232/Y vdd OAI21X1
XOAI21X1_298 BUFX4_389/Y BUFX4_458/Y OAI21X1_895/A gnd OAI21X1_299/C vdd OAI21X1
XOAI21X1_276 BUFX4_135/Y BUFX4_163/Y AOI21X1_455/A gnd OAI21X1_276/Y vdd OAI21X1
XOAI21X1_287 BUFX4_465/Y NAND2X1_74/Y OAI21X1_286/Y gnd OAI21X1_287/Y vdd OAI21X1
XINVX1_307 INVX1_307/A gnd INVX1_307/Y vdd INVX1
XAND2X2_10 AND2X2_10/A AND2X2_10/B gnd AND2X2_10/Y vdd AND2X2
XINVX1_329 INVX1_329/A gnd INVX1_329/Y vdd INVX1
XAND2X2_21 BUFX4_78/Y AND2X2_21/B gnd AND2X2_21/Y vdd AND2X2
XAND2X2_32 AND2X2_32/A AND2X2_32/B gnd AND2X2_32/Y vdd AND2X2
XINVX1_318 INVX1_318/A gnd INVX1_318/Y vdd INVX1
XAND2X2_54 AND2X2_54/A BUFX4_392/Y gnd AND2X2_54/Y vdd AND2X2
XAND2X2_43 AND2X2_43/A BUFX4_95/Y gnd AND2X2_43/Y vdd AND2X2
XDFFPOSX1_190 INVX1_227/A CLKBUF1_65/Y MUX2X1_290/Y gnd vdd DFFPOSX1
XNAND2X1_271 AND2X2_52/A NOR2X1_657/A gnd OAI21X1_911/C vdd NAND2X1
XNAND2X1_260 NOR2X1_295/A BUFX4_282/Y gnd OAI21X1_870/C vdd NAND2X1
XNAND2X1_293 BUFX4_226/Y NOR2X1_735/A gnd OAI21X1_971/C vdd NAND2X1
XNAND2X1_282 AND2X2_25/B NAND2X1_282/B gnd OAI21X1_946/C vdd NAND2X1
XFILL_45_5_0 gnd vdd FILL
XNOR2X1_709 NOR2X1_709/A NOR2X1_707/B gnd NOR2X1_709/Y vdd NOR2X1
XOAI21X1_1506 BUFX4_439/Y NAND2X1_77/Y OAI21X1_1506/C gnd DFFPOSX1_515/D vdd OAI21X1
XOAI21X1_1539 BUFX4_189/Y BUFX4_312/Y AND2X2_30/B gnd OAI21X1_1540/C vdd OAI21X1
XOAI21X1_1528 NAND2X1_79/Y AND2X2_6/B OAI21X1_1528/C gnd DFFPOSX1_538/D vdd OAI21X1
XOAI21X1_1517 BUFX4_313/Y BUFX4_300/Y INVX1_385/A gnd OAI21X1_1518/C vdd OAI21X1
XFILL_36_5_0 gnd vdd FILL
XFILL_20_9_1 gnd vdd FILL
XCLKBUF1_41 BUFX4_8/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XCLKBUF1_30 BUFX4_7/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XCLKBUF1_63 BUFX4_10/Y gnd CLKBUF1_63/Y vdd CLKBUF1
XCLKBUF1_52 BUFX4_6/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XCLKBUF1_74 BUFX4_4/Y gnd CLKBUF1_74/Y vdd CLKBUF1
XCLKBUF1_85 BUFX4_2/Y gnd CLKBUF1_85/Y vdd CLKBUF1
XCLKBUF1_96 BUFX4_3/Y gnd CLKBUF1_96/Y vdd CLKBUF1
XFILL_2_5_0 gnd vdd FILL
XFILL_27_5_0 gnd vdd FILL
XFILL_11_9_1 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd MUX2X1_91/B vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XBUFX4_413 address[2] gnd BUFX4_413/Y vdd BUFX4
XBUFX4_402 address[5] gnd BUFX4_402/Y vdd BUFX4
XBUFX4_435 INVX8_23/Y gnd BUFX4_435/Y vdd BUFX4
XBUFX4_424 INVX8_3/Y gnd BUFX4_424/Y vdd BUFX4
XBUFX4_446 INVX8_2/Y gnd MUX2X1_9/B vdd BUFX4
XBUFX4_468 INVX8_15/Y gnd BUFX4_468/Y vdd BUFX4
XNOR2X1_506 NOR2X1_288/A BUFX4_326/Y gnd NOR2X1_506/Y vdd NOR2X1
XBUFX4_479 INVX8_16/Y gnd BUFX4_479/Y vdd BUFX4
XFILL_18_5_0 gnd vdd FILL
XNOR2X1_517 NOR2X1_517/A BUFX4_155/Y gnd NOR2X1_517/Y vdd NOR2X1
XBUFX4_457 INVX8_25/Y gnd BUFX4_457/Y vdd BUFX4
XNOR2X1_539 BUFX4_288/Y NOR2X1_539/B gnd NOR2X1_539/Y vdd NOR2X1
XNOR2X1_528 NOR2X1_528/A BUFX4_353/Y gnd NOR2X1_528/Y vdd NOR2X1
XAOI21X1_119 BUFX4_177/Y MUX2X1_364/S NOR2X1_193/Y gnd AOI21X1_119/Y vdd AOI21X1
XAOI21X1_108 BUFX4_466/Y MUX2X1_102/S NOR2X1_176/Y gnd AOI21X1_108/Y vdd AOI21X1
XOAI21X1_1303 BUFX4_67/Y NAND2X1_37/Y OAI21X1_1302/Y gnd OAI21X1_1303/Y vdd OAI21X1
XOAI21X1_1314 BUFX4_449/Y BUFX4_53/Y NOR2X1_367/B gnd OAI21X1_1314/Y vdd OAI21X1
XOAI21X1_1347 BUFX4_63/Y NAND2X1_51/Y OAI21X1_1347/C gnd OAI21X1_1347/Y vdd OAI21X1
XOAI21X1_1325 BUFX4_57/Y BUFX4_398/Y AOI21X1_319/B gnd OAI21X1_1326/C vdd OAI21X1
XOAI21X1_1336 BUFX4_121/Y BUFX4_395/Y INVX1_343/A gnd OAI21X1_1336/Y vdd OAI21X1
XDFFPOSX1_904 NOR2X1_165/A CLKBUF1_71/Y AOI21X1_100/Y gnd vdd DFFPOSX1
XDFFPOSX1_915 OAI21X1_696/A CLKBUF1_39/Y OAI21X1_225/Y gnd vdd DFFPOSX1
XDFFPOSX1_948 OAI21X1_898/A CLKBUF1_61/Y OAI21X1_251/Y gnd vdd DFFPOSX1
XOAI21X1_1358 NOR2X1_84/B BUFX4_185/Y INVX1_250/A gnd OAI21X1_1358/Y vdd OAI21X1
XOAI21X1_1369 NAND2X1_56/Y BUFX4_428/Y OAI21X1_1369/C gnd DFFPOSX1_287/D vdd OAI21X1
XDFFPOSX1_937 NOR2X1_182/A CLKBUF1_54/Y AOI21X1_112/Y gnd vdd DFFPOSX1
XDFFPOSX1_926 INVX1_119/A CLKBUF1_29/Y MUX2X1_106/Y gnd vdd DFFPOSX1
XDFFPOSX1_959 NOR2X1_197/A CLKBUF1_37/Y AOI21X1_122/Y gnd vdd DFFPOSX1
XAOI21X1_620 BUFX4_67/Y NOR2X1_733/B NOR2X1_732/Y gnd AOI21X1_620/Y vdd AOI21X1
XINVX4_12 INVX4_12/A gnd INVX4_12/Y vdd INVX4
XFILL_43_8_1 gnd vdd FILL
XFILL_42_3_0 gnd vdd FILL
XBUFX4_221 BUFX4_21/Y gnd INVX8_31/A vdd BUFX4
XBUFX4_210 INVX8_11/Y gnd MUX2X1_97/B vdd BUFX4
XBUFX4_232 BUFX4_24/Y gnd BUFX4_232/Y vdd BUFX4
XBUFX4_254 BUFX4_23/Y gnd AND2X2_27/A vdd BUFX4
XBUFX4_243 BUFX4_22/Y gnd AND2X2_47/B vdd BUFX4
XNOR2X1_325 INVX1_200/Y OAI22X1_2/C gnd AOI22X1_6/A vdd NOR2X1
XNOR2X1_314 NOR2X1_314/A NOR2X1_312/Y gnd INVX2_20/A vdd NOR2X1
XBUFX4_276 BUFX4_24/Y gnd BUFX4_276/Y vdd BUFX4
XBUFX4_287 BUFX4_18/Y gnd BUFX4_287/Y vdd BUFX4
XBUFX4_265 BUFX4_18/Y gnd BUFX4_265/Y vdd BUFX4
XBUFX4_298 BUFX4_302/A gnd BUFX4_298/Y vdd BUFX4
XNOR2X1_303 XNOR2X1_1/B INVX1_188/Y gnd MUX2X1_174/B vdd NOR2X1
XNOR2X1_358 INVX4_9/A AND2X2_17/A gnd NOR2X1_358/Y vdd NOR2X1
XNOR2X1_347 AND2X2_2/B AOI22X1_5/D gnd NOR2X1_347/Y vdd NOR2X1
XNOR2X1_336 NOR2X1_336/A NOR2X1_336/B gnd AOI22X1_7/C vdd NOR2X1
XFILL_34_8_1 gnd vdd FILL
XNOR2X1_369 BUFX4_246/Y INVX1_238/Y gnd NOR2X1_369/Y vdd NOR2X1
XFILL_25_2 gnd vdd FILL
XFILL_33_3_0 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XOAI21X1_809 BUFX4_364/Y NOR2X1_46/A BUFX4_149/Y gnd OAI22X1_23/C vdd OAI21X1
XOAI21X1_1100 BUFX4_370/Y NOR2X1_652/A BUFX4_156/Y gnd OAI21X1_1102/B vdd OAI21X1
XOAI21X1_1122 OAI22X1_57/Y BUFX4_34/Y BUFX4_165/Y gnd OAI22X1_59/B vdd OAI21X1
XOAI21X1_1111 BUFX4_283/Y OAI21X1_1436/C BUFX4_98/Y gnd OAI21X1_1112/B vdd OAI21X1
XOAI21X1_1144 BUFX4_332/Y NOR2X1_31/A BUFX4_149/Y gnd OAI22X1_64/C vdd OAI21X1
XDFFPOSX1_712 INVX1_45/A CLKBUF1_19/Y MUX2X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_701 NOR2X1_499/A CLKBUF1_19/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XOAI21X1_1133 BUFX4_226/Y OAI21X1_1133/B BUFX4_108/Y gnd OAI21X1_1134/B vdd OAI21X1
XMUX2X1_309 INVX1_452/Y MUX2X1_9/B MUX2X1_71/S gnd MUX2X1_309/Y vdd MUX2X1
XDFFPOSX1_723 NOR2X1_78/A CLKBUF1_68/Y AOI21X1_40/Y gnd vdd DFFPOSX1
XOAI21X1_1155 AOI21X1_483/Y AOI21X1_484/Y BUFX4_33/Y gnd NAND2X1_337/A vdd OAI21X1
XOAI21X1_1166 INVX1_436/Y BUFX4_249/Y NAND2X1_338/Y gnd MUX2X1_259/B vdd OAI21X1
XDFFPOSX1_745 INVX1_399/A CLKBUF1_23/Y OAI21X1_106/Y gnd vdd DFFPOSX1
XDFFPOSX1_734 NOR2X1_85/A CLKBUF1_23/Y AOI21X1_45/Y gnd vdd DFFPOSX1
XOAI21X1_1177 OAI21X1_1177/A INVX4_14/Y INVX4_13/Y gnd OAI22X1_94/C vdd OAI21X1
XDFFPOSX1_756 INVX1_66/A CLKBUF1_18/Y MUX2X1_56/Y gnd vdd DFFPOSX1
XOAI21X1_1188 AOI21X1_495/Y AOI21X1_496/Y BUFX4_40/Y gnd NAND2X1_342/B vdd OAI21X1
XDFFPOSX1_778 INVX1_76/A CLKBUF1_95/Y MUX2X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_767 NOR2X1_97/A CLKBUF1_102/Y AOI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_789 INVX1_83/A CLKBUF1_6/Y MUX2X1_73/Y gnd vdd DFFPOSX1
XOAI21X1_1199 OAI22X1_71/Y BUFX4_37/Y BUFX4_206/Y gnd OAI22X1_72/A vdd OAI21X1
XFILL_0_8_1 gnd vdd FILL
XFILL_25_8_1 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XAOI21X1_461 address[6] MUX2X1_255/Y INVX4_13/Y gnd AOI22X1_33/B vdd AOI21X1
XAOI21X1_450 NOR2X1_292/A BUFX4_224/Y AOI21X1_450/C gnd NOR2X1_508/B vdd AOI21X1
XAOI21X1_483 BUFX4_340/Y INVX1_427/Y AOI21X1_483/C gnd AOI21X1_483/Y vdd AOI21X1
XAOI21X1_472 AOI21X1_472/A BUFX4_342/Y BUFX4_151/Y gnd AOI21X1_473/B vdd AOI21X1
XAOI21X1_494 BUFX4_259/Y INVX1_60/Y BUFX4_81/Y gnd AOI21X1_494/Y vdd AOI21X1
XFILL_8_9_1 gnd vdd FILL
XNAND3X1_10 NOR2X1_300/B AND2X2_3/A OR2X2_2/B gnd NAND3X1_10/Y vdd NAND3X1
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_32 INVX1_194/Y NAND3X1_32/B INVX1_195/Y gnd NAND3X1_32/Y vdd NAND3X1
XNAND3X1_21 INVX2_14/Y NAND3X1_21/B NAND3X1_20/Y gnd AND2X2_7/A vdd NAND3X1
XNAND3X1_65 INVX4_9/Y INVX1_211/Y NAND3X1_65/C gnd AND2X2_14/B vdd NAND3X1
XNAND3X1_43 INVX1_202/Y NAND3X1_43/B NAND3X1_43/C gnd XNOR2X1_4/A vdd NAND3X1
XNAND3X1_54 INVX2_19/Y INVX4_10/Y NAND3X1_54/C gnd NAND3X1_54/Y vdd NAND3X1
XNAND3X1_76 BUFX4_41/Y NAND3X1_76/B NAND3X1_76/C gnd NAND3X1_76/Y vdd NAND3X1
XNOR2X1_10 NOR2X1_2/A INVX1_14/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_21 INVX2_5/Y XNOR2X1_8/A gnd INVX8_7/A vdd NOR2X1
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_54 BUFX4_42/Y BUFX4_57/Y gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_32 INVX1_23/Y XNOR2X1_8/A gnd INVX8_9/A vdd NOR2X1
XNOR2X1_65 BUFX4_46/Y BUFX4_133/Y gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_87 NOR2X1_87/A MUX2X1_50/S gnd NOR2X1_87/Y vdd NOR2X1
XFILL_16_8_1 gnd vdd FILL
XNOR2X1_76 NOR2X1_76/A NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNOR2X1_98 NOR2X1_98/A NOR2X1_97/B gnd NOR2X1_98/Y vdd NOR2X1
XNAND2X1_9 NOR2X1_10/Y NOR2X1_6/Y gnd MUX2X1_9/S vdd NAND2X1
XNOR2X1_100 NOR2X1_100/A NOR2X1_97/B gnd NOR2X1_100/Y vdd NOR2X1
XNOR2X1_133 AND2X2_44/A MUX2X1_88/S gnd NOR2X1_133/Y vdd NOR2X1
XNOR2X1_111 INVX1_290/A AOI21X1_62/B gnd NOR2X1_111/Y vdd NOR2X1
XNOR2X1_122 NOR2X1_122/A MUX2X1_320/S gnd NOR2X1_122/Y vdd NOR2X1
XMUX2X1_50 BUFX4_469/Y INVX1_60/Y MUX2X1_50/S gnd MUX2X1_50/Y vdd MUX2X1
XMUX2X1_72 INVX1_82/Y MUX2X1_77/B MUX2X1_71/S gnd MUX2X1_72/Y vdd MUX2X1
XMUX2X1_61 INVX1_71/Y MUX2X1_61/B MUX2X1_59/S gnd MUX2X1_61/Y vdd MUX2X1
XNOR2X1_155 NOR2X1_155/A NOR2X1_155/B gnd AOI21X1_92/C vdd NOR2X1
XMUX2X1_94 MUX2X1_49/A MUX2X1_94/B MUX2X1_94/S gnd MUX2X1_94/Y vdd MUX2X1
XNOR2X1_144 NOR2X1_144/A MUX2X1_92/S gnd AOI21X1_85/C vdd NOR2X1
XMUX2X1_83 INVX1_96/Y MUX2X1_83/B MUX2X1_81/S gnd MUX2X1_83/Y vdd MUX2X1
XNOR2X1_166 NOR2X1_166/A NOR2X1_167/B gnd NOR2X1_166/Y vdd NOR2X1
XNOR2X1_199 NOR2X1_199/A NOR2X1_703/B gnd NOR2X1_199/Y vdd NOR2X1
XNOR2X1_188 NOR2X1_188/A NOR2X1_188/B gnd NOR2X1_188/Y vdd NOR2X1
XNOR2X1_177 BUFX4_139/Y NOR2X1_96/B gnd MUX2X1_108/S vdd NOR2X1
XOAI21X1_606 BUFX4_272/Y MUX2X1_182/Y AOI21X1_281/Y gnd AOI22X1_15/B vdd OAI21X1
XOAI21X1_628 INVX1_274/Y BUFX4_224/Y NAND2X1_193/Y gnd MUX2X1_188/A vdd OAI21X1
XOAI21X1_617 BUFX4_146/Y OAI21X1_617/B AND2X2_36/B gnd OAI21X1_617/Y vdd OAI21X1
XOAI21X1_639 OAI21X1_639/A OAI21X1_639/B BUFX4_205/Y gnd AOI21X1_297/C vdd OAI21X1
XMUX2X1_117 INVX1_130/Y BUFX4_466/Y MUX2X1_366/S gnd MUX2X1_117/Y vdd MUX2X1
XDFFPOSX1_520 INVX1_321/A CLKBUF1_34/Y MUX2X1_386/Y gnd vdd DFFPOSX1
XMUX2X1_128 BUFX4_217/Y INVX1_141/Y NOR2X1_233/Y gnd MUX2X1_128/Y vdd MUX2X1
XDFFPOSX1_531 INVX1_261/A CLKBUF1_36/Y MUX2X1_389/Y gnd vdd DFFPOSX1
XMUX2X1_106 INVX1_119/Y BUFX4_465/Y MUX2X1_353/S gnd MUX2X1_106/Y vdd MUX2X1
XDFFPOSX1_553 INVX1_388/A CLKBUF1_57/Y MUX2X1_396/Y gnd vdd DFFPOSX1
XDFFPOSX1_564 INVX1_327/A CLKBUF1_73/Y MUX2X1_402/Y gnd vdd DFFPOSX1
XMUX2X1_139 INVX1_152/Y MUX2X1_40/B MUX2X1_406/S gnd MUX2X1_139/Y vdd MUX2X1
XDFFPOSX1_542 INVX1_441/A CLKBUF1_64/Y MUX2X1_393/Y gnd vdd DFFPOSX1
XDFFPOSX1_575 INVX1_270/A CLKBUF1_70/Y MUX2X1_404/Y gnd vdd DFFPOSX1
XDFFPOSX1_586 OAI21X1_1133/B CLKBUF1_25/Y OAI21X1_1560/Y gnd vdd DFFPOSX1
XDFFPOSX1_597 INVX1_6/A CLKBUF1_78/Y MUX2X1_3/Y gnd vdd DFFPOSX1
XINVX1_13 NOR2X1_1/B gnd NOR2X1_9/B vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XDFFPOSX1_9 DFFPOSX1_9/Q CLKBUF1_92/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XFILL_40_6_1 gnd vdd FILL
XAOI21X1_291 NAND2X1_361/A BUFX4_346/Y AND2X2_33/B gnd AOI21X1_291/Y vdd AOI21X1
XAOI21X1_280 INVX8_29/A MUX2X1_181/Y AOI21X1_280/C gnd NAND2X1_181/B vdd AOI21X1
XFILL_48_7_1 gnd vdd FILL
XFILL_47_2_0 gnd vdd FILL
XFILL_31_6_1 gnd vdd FILL
XFILL_30_1_0 gnd vdd FILL
XFILL_39_7_1 gnd vdd FILL
XFILL_38_2_0 gnd vdd FILL
XOAI22X1_19 OAI22X1_19/A OAI22X1_19/B OAI22X1_19/C OAI22X1_19/D gnd OAI22X1_19/Y vdd
+ OAI22X1
XFILL_22_6_1 gnd vdd FILL
XOAI21X1_403 BUFX4_125/Y BUFX4_294/Y OAI21X1_403/C gnd OAI21X1_404/C vdd OAI21X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 MUX2X1_71/B OAI21X1_48/B OAI21X1_414/C gnd OAI21X1_414/Y vdd OAI21X1
XOAI21X1_447 AND2X2_1/Y traffic_Street_1[2] traffic_Street_1[3] gnd NAND3X1_28/C vdd
+ OAI21X1
XOAI21X1_436 BUFX4_470/Y OAI21X1_64/B OAI21X1_435/Y gnd OAI21X1_436/Y vdd OAI21X1
XOAI21X1_425 INVX4_4/A BUFX4_464/Y INVX1_401/A gnd OAI21X1_425/Y vdd OAI21X1
XOAI21X1_458 AOI22X1_10/D BUFX4_320/Y INVX1_214/A gnd NAND3X1_21/B vdd OAI21X1
XOAI21X1_469 AND2X2_3/Y NOR3X1_1/B INVX4_8/A gnd NAND3X1_29/A vdd OAI21X1
XDFFPOSX1_383 NOR2X1_633/A CLKBUF1_24/Y AOI21X1_521/Y gnd vdd DFFPOSX1
XDFFPOSX1_350 INVX1_452/A CLKBUF1_99/Y MUX2X1_309/Y gnd vdd DFFPOSX1
XDFFPOSX1_361 INVX1_417/A CLKBUF1_58/Y MUX2X1_308/Y gnd vdd DFFPOSX1
XDFFPOSX1_372 INVX1_363/A CLKBUF1_83/Y DFFPOSX1_372/D gnd vdd DFFPOSX1
XDFFPOSX1_394 BUFX2_3/A CLKBUF1_3/Y INVX4_9/A gnd vdd DFFPOSX1
XFILL_5_7_1 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_970 INVX1_388/Y BUFX4_225/Y NAND2X1_292/Y gnd MUX2X1_238/A vdd OAI21X1
XOAI21X1_981 AOI21X1_427/Y OAI21X1_981/B NAND3X1_78/Y gnd AOI22X1_27/C vdd OAI21X1
XOAI21X1_992 BUFX4_31/Y MUX2X1_240/Y OAI21X1_992/C gnd NAND2X1_299/B vdd OAI21X1
XOAI21X1_30 NAND2X1_24/Y BUFX4_421/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 OAI21X1_54/A MUX2X1_9/B OAI21X1_51/Y gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_63 BUFX4_190/Y BUFX4_462/Y OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_41 NOR2X1_39/A INVX4_2/A OAI21X1_41/C gnd OAI21X1_42/C vdd OAI21X1
XOAI21X1_85 BUFX4_124/Y BUFX4_42/Y OAI21X1_85/C gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_74 NAND2X1_30/Y BUFX4_473/Y OAI21X1_73/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 NAND2X1_36/Y MUX2X1_49/A OAI21X1_96/C gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_211 NAND2X1_61/Y BUFX4_174/Y OAI21X1_210/Y gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_200 BUFX4_143/Y BUFX4_404/Y NAND2X1_219/A gnd OAI21X1_201/C vdd OAI21X1
XOAI21X1_222 BUFX4_119/Y BUFX4_408/Y OAI21X1_222/C gnd OAI21X1_222/Y vdd OAI21X1
XOAI21X1_244 BUFX4_60/Y BUFX4_435/Y OAI21X1_244/C gnd OAI21X1_244/Y vdd OAI21X1
XOAI21X1_255 NAND2X1_69/Y BUFX4_466/Y OAI21X1_255/C gnd OAI21X1_255/Y vdd OAI21X1
XOAI21X1_233 NAND2X1_66/Y MUX2X1_97/B OAI21X1_232/Y gnd OAI21X1_233/Y vdd OAI21X1
XOAI21X1_288 BUFX4_458/Y BUFX4_300/Y NOR2X1_383/A gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_299 NAND2X1_76/Y BUFX4_176/Y OAI21X1_299/C gnd OAI21X1_299/Y vdd OAI21X1
XOAI21X1_266 BUFX4_452/Y BUFX4_162/Y NOR2X1_469/A gnd OAI21X1_267/C vdd OAI21X1
XOAI21X1_277 MUX2X1_57/A NAND2X1_73/Y OAI21X1_276/Y gnd OAI21X1_277/Y vdd OAI21X1
XINVX1_308 INVX1_308/A gnd INVX1_308/Y vdd INVX1
XAND2X2_11 AND2X2_11/A AOI22X1_5/Y gnd AND2X2_11/Y vdd AND2X2
XAND2X2_22 AND2X2_22/A AND2X2_22/B gnd AND2X2_22/Y vdd AND2X2
XINVX1_319 INVX1_319/A gnd INVX1_319/Y vdd INVX1
XAND2X2_44 AND2X2_44/A BUFX4_250/Y gnd AND2X2_44/Y vdd AND2X2
XAND2X2_55 AND2X2_55/A BUFX4_258/Y gnd AND2X2_55/Y vdd AND2X2
XAND2X2_33 AND2X2_33/A AND2X2_33/B gnd AND2X2_33/Y vdd AND2X2
XDFFPOSX1_180 INVX1_346/A CLKBUF1_38/Y MUX2X1_277/Y gnd vdd DFFPOSX1
XDFFPOSX1_191 INVX1_291/A CLKBUF1_22/Y MUX2X1_291/Y gnd vdd DFFPOSX1
XNAND2X1_250 NOR2X1_93/A BUFX4_257/Y gnd OAI21X1_834/C vdd NAND2X1
XNAND2X1_261 NAND2X1_261/A BUFX4_284/Y gnd OAI21X1_871/C vdd NAND2X1
XNAND2X1_283 BUFX4_273/Y NOR2X1_668/A gnd NAND2X1_283/Y vdd NAND2X1
XNAND2X1_294 AND2X2_37/B NOR2X1_738/A gnd NAND2X1_294/Y vdd NAND2X1
XNAND2X1_272 BUFX4_247/Y NOR2X1_660/A gnd NAND2X1_272/Y vdd NAND2X1
XFILL_45_5_1 gnd vdd FILL
XFILL_44_0_0 gnd vdd FILL
XOAI21X1_1529 NOR2X1_84/B BUFX4_309/Y INVX1_262/A gnd OAI21X1_1530/C vdd OAI21X1
XOAI21X1_1507 BUFX4_132/Y BUFX4_459/Y NAND2X1_242/B gnd OAI21X1_1508/C vdd OAI21X1
XOAI21X1_1518 NAND2X1_78/Y BUFX4_73/Y OAI21X1_1518/C gnd OAI21X1_1518/Y vdd OAI21X1
XFILL_48_1 gnd vdd FILL
XFILL_36_5_1 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XCLKBUF1_31 BUFX4_1/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_42 BUFX4_5/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_20 BUFX4_2/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_53 BUFX4_1/Y gnd CLKBUF1_53/Y vdd CLKBUF1
XCLKBUF1_75 BUFX4_5/Y gnd CLKBUF1_75/Y vdd CLKBUF1
XCLKBUF1_64 BUFX4_5/Y gnd CLKBUF1_64/Y vdd CLKBUF1
XCLKBUF1_86 BUFX4_8/Y gnd CLKBUF1_86/Y vdd CLKBUF1
XCLKBUF1_97 BUFX4_6/Y gnd CLKBUF1_97/Y vdd CLKBUF1
XFILL_2_5_1 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_10_4_1 gnd vdd FILL
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XINVX1_105 INVX1_105/A gnd MUX2X1_92/B vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XBUFX4_403 INVX8_21/Y gnd BUFX4_403/Y vdd BUFX4
XBUFX4_414 address[2] gnd BUFX4_414/Y vdd BUFX4
XBUFX4_447 BUFX4_449/A gnd INVX4_4/A vdd BUFX4
XBUFX4_425 INVX8_3/Y gnd MUX2X1_27/B vdd BUFX4
XBUFX4_436 INVX8_2/Y gnd AND2X2_5/B vdd BUFX4
XNOR2X1_507 BUFX4_201/Y NOR2X1_507/B gnd NOR2X1_507/Y vdd NOR2X1
XFILL_18_5_1 gnd vdd FILL
XBUFX4_469 INVX8_15/Y gnd BUFX4_469/Y vdd BUFX4
XBUFX4_458 INVX8_25/Y gnd BUFX4_458/Y vdd BUFX4
XFILL_17_0_0 gnd vdd FILL
XNOR2X1_518 NOR2X1_518/A BUFX4_82/Y gnd NOR2X1_518/Y vdd NOR2X1
XNOR2X1_529 BUFX4_413/Y OAI22X1_51/Y gnd NOR2X1_529/Y vdd NOR2X1
XAOI21X1_109 MUX2X1_97/B MUX2X1_108/S NOR2X1_178/Y gnd AOI21X1_109/Y vdd AOI21X1
XOAI21X1_1304 BUFX4_193/Y BUFX4_479/Y AOI21X1_467/B gnd OAI21X1_1305/C vdd OAI21X1
XOAI21X1_1326 MUX2X1_18/B NAND2X1_44/Y OAI21X1_1326/C gnd DFFPOSX1_355/D vdd OAI21X1
XOAI21X1_1337 NAND2X1_48/Y BUFX4_69/Y OAI21X1_1336/Y gnd OAI21X1_1337/Y vdd OAI21X1
XDFFPOSX1_905 NOR2X1_166/A CLKBUF1_74/Y AOI21X1_101/Y gnd vdd DFFPOSX1
XOAI21X1_1315 NAND2X1_40/Y BUFX4_443/Y OAI21X1_1314/Y gnd DFFPOSX1_374/D vdd OAI21X1
XDFFPOSX1_938 NOR2X1_183/A CLKBUF1_41/Y AOI21X1_113/Y gnd vdd DFFPOSX1
XDFFPOSX1_927 NOR2X1_178/A CLKBUF1_27/Y AOI21X1_109/Y gnd vdd DFFPOSX1
XOAI21X1_1359 NAND2X1_53/Y BUFX4_439/Y OAI21X1_1358/Y gnd DFFPOSX1_306/D vdd OAI21X1
XOAI21X1_1348 BUFX4_59/Y BUFX4_184/Y OAI21X1_1348/C gnd OAI21X1_1348/Y vdd OAI21X1
XDFFPOSX1_916 AND2X2_32/A CLKBUF1_29/Y OAI21X1_227/Y gnd vdd DFFPOSX1
XDFFPOSX1_949 OAI21X1_252/C CLKBUF1_9/Y OAI21X1_253/Y gnd vdd DFFPOSX1
XAOI21X1_610 BUFX4_318/Y NOR2X1_231/B NOR2X1_722/Y gnd AOI21X1_610/Y vdd AOI21X1
XAOI21X1_621 BUFX4_322/Y NOR2X1_733/B NOR2X1_733/Y gnd AOI21X1_621/Y vdd AOI21X1
XINVX4_13 street gnd INVX4_13/Y vdd INVX4
XFILL_42_3_1 gnd vdd FILL
XBUFX4_211 INVX8_11/Y gnd MUX2X1_39/B vdd BUFX4
XBUFX4_200 address[3] gnd INVX8_29/A vdd BUFX4
XBUFX4_233 BUFX4_24/Y gnd BUFX4_233/Y vdd BUFX4
XBUFX4_255 BUFX4_24/Y gnd BUFX4_255/Y vdd BUFX4
XBUFX4_222 BUFX4_17/Y gnd BUFX4_222/Y vdd BUFX4
XBUFX4_244 BUFX4_22/Y gnd BUFX4_244/Y vdd BUFX4
XBUFX4_266 BUFX4_18/Y gnd BUFX4_266/Y vdd BUFX4
XBUFX4_277 BUFX4_17/Y gnd BUFX4_277/Y vdd BUFX4
XBUFX4_288 BUFX4_22/Y gnd BUFX4_288/Y vdd BUFX4
XNOR2X1_304 traffic_Street_0[0] traffic_Street_0[1] gnd NOR2X1_304/Y vdd NOR2X1
XNOR2X1_315 INVX2_19/A INVX2_18/Y gnd INVX1_201/A vdd NOR2X1
XNOR2X1_359 INVX4_9/Y AND2X2_18/Y gnd NOR2X1_359/Y vdd NOR2X1
XNOR2X1_348 INVX2_17/Y BUFX4_306/Y gnd NAND3X1_68/A vdd NOR2X1
XNOR2X1_337 INVX2_13/Y XNOR2X1_4/A gnd AOI22X1_7/B vdd NOR2X1
XBUFX4_299 BUFX4_302/A gnd BUFX4_299/Y vdd BUFX4
XNOR2X1_326 INVX2_19/A AND2X2_8/A gnd NOR2X1_326/Y vdd NOR2X1
XFILL_33_3_1 gnd vdd FILL
XOAI21X1_1101 BUFX4_370/Y INVX1_451/A AOI21X1_469/Y gnd OAI21X1_1102/C vdd OAI21X1
XOAI21X1_1112 NOR2X1_532/Y OAI21X1_1112/B OAI21X1_1110/Y gnd AOI21X1_475/B vdd OAI21X1
XOAI21X1_1156 BUFX4_362/Y NOR2X1_706/A BUFX4_156/Y gnd AOI21X1_485/C vdd OAI21X1
XOAI21X1_1145 OAI21X1_33/C BUFX4_233/Y BUFX4_111/Y gnd OAI22X1_64/B vdd OAI21X1
XOAI21X1_1134 NOR2X1_551/Y OAI21X1_1134/B OAI21X1_1132/Y gnd OAI21X1_1134/Y vdd OAI21X1
XDFFPOSX1_713 INVX1_46/A CLKBUF1_19/Y MUX2X1_38/Y gnd vdd DFFPOSX1
XOAI21X1_1123 BUFX4_354/Y DFFPOSX1_249/Q BUFX4_150/Y gnd OAI22X1_58/C vdd OAI21X1
XDFFPOSX1_702 NOR2X1_574/A CLKBUF1_24/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XOAI21X1_1167 INVX1_437/Y BUFX4_251/Y NAND2X1_339/Y gnd MUX2X1_259/A vdd OAI21X1
XDFFPOSX1_735 NOR2X1_87/A CLKBUF1_57/Y AOI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_746 NOR2X1_569/A CLKBUF1_23/Y OAI21X1_108/Y gnd vdd DFFPOSX1
XOAI21X1_1178 NOR2X1_85/A BUFX4_260/Y AOI21X1_494/Y gnd OAI21X1_1178/Y vdd OAI21X1
XDFFPOSX1_724 INVX1_53/A CLKBUF1_38/Y MUX2X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_757 INVX1_67/A CLKBUF1_18/Y MUX2X1_57/Y gnd vdd DFFPOSX1
XOAI21X1_1189 BUFX4_358/Y OAI21X1_131/C BUFX4_158/Y gnd OAI21X1_1189/Y vdd OAI21X1
XDFFPOSX1_768 NOR2X1_98/A CLKBUF1_38/Y AOI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_779 INVX1_77/A CLKBUF1_63/Y MUX2X1_67/Y gnd vdd DFFPOSX1
XFILL_24_3_1 gnd vdd FILL
XAOI21X1_440 NOR2X1_88/A BUFX4_150/Y BUFX4_329/Y gnd AOI21X1_440/Y vdd AOI21X1
XAOI21X1_451 INVX1_161/Y BUFX4_227/Y AOI21X1_451/C gnd AOI21X1_451/Y vdd AOI21X1
XAOI21X1_495 INVX1_52/A AND2X2_29/A AOI21X1_495/C gnd AOI21X1_495/Y vdd AOI21X1
XAOI21X1_462 NOR2X1_639/A BUFX4_152/Y BUFX4_262/Y gnd AOI21X1_462/Y vdd AOI21X1
XAOI21X1_484 BUFX4_240/Y INVX1_428/Y AOI21X1_484/C gnd AOI21X1_484/Y vdd AOI21X1
XAOI21X1_473 AOI21X1_473/A AOI21X1_473/B AOI21X1_473/C gnd AOI21X1_475/C vdd AOI21X1
XNAND3X1_11 INVX2_14/A NAND3X1_10/Y NAND3X1_11/C gnd NAND3X1_13/A vdd NAND3X1
XFILL_7_4_1 gnd vdd FILL
XNAND3X1_22 traffic_Street_0[3] INVX1_189/A NAND3X1_22/C gnd NAND3X1_23/C vdd NAND3X1
XNAND3X1_33 INVX2_20/A NAND3X1_43/B NAND3X1_43/C gnd AND2X2_8/A vdd NAND3X1
XNAND3X1_55 INVX4_9/A NAND3X1_54/Y NAND3X1_55/C gnd NAND3X1_55/Y vdd NAND3X1
XNAND3X1_44 INVX4_9/A NAND3X1_40/Y NAND3X1_44/C gnd NAND3X1_44/Y vdd NAND3X1
XNAND3X1_66 NAND3X1_66/A AOI22X1_9/Y NAND3X1_66/C gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_77 BUFX4_390/Y NAND3X1_76/Y NAND3X1_77/C gnd NAND3X1_77/Y vdd NAND3X1
XNOR2X1_11 INVX2_4/Y NOR2X1_9/B gnd INVX1_23/A vdd NOR2X1
XNOR2X1_33 NOR2X1_16/A BUFX4_191/Y gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_22 BUFX4_294/Y BUFX4_144/Y gnd AOI21X1_7/B vdd NOR2X1
XNOR2X1_55 NOR2X1_55/A NOR2X1_54/Y gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_44 BUFX4_461/Y NOR2X1_96/B gnd NOR2X1_47/B vdd NOR2X1
XNOR2X1_66 NOR2X1_66/A NOR2X1_65/Y gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_88 NOR2X1_88/A MUX2X1_50/S gnd NOR2X1_88/Y vdd NOR2X1
XNOR2X1_77 NOR2X1_74/B NOR2X1_77/B gnd MUX2X1_45/S vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_99 NOR2X1_99/A NOR2X1_97/B gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_123 NOR2X1_123/A MUX2X1_320/S gnd AOI21X1_70/C vdd NOR2X1
XNOR2X1_101 INVX2_9/Y INVX2_8/Y gnd INVX8_18/A vdd NOR2X1
XMUX2X1_40 INVX1_50/Y MUX2X1_40/B MUX2X1_42/S gnd MUX2X1_40/Y vdd MUX2X1
XNOR2X1_112 NOR2X1_112/A AOI21X1_62/B gnd AOI21X1_63/C vdd NOR2X1
XMUX2X1_51 INVX1_61/Y MUX2X1_59/B MUX2X1_51/S gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_62 INVX1_72/Y MUX2X1_66/B MUX2X1_59/S gnd MUX2X1_62/Y vdd MUX2X1
XMUX2X1_95 AND2X2_2/B MUX2X1_95/B MUX2X1_96/S gnd MUX2X1_95/Y vdd MUX2X1
XNOR2X1_167 NOR2X1_589/A NOR2X1_167/B gnd NOR2X1_167/Y vdd NOR2X1
XNOR2X1_134 NOR2X1_134/A MUX2X1_88/S gnd AOI21X1_78/C vdd NOR2X1
XNOR2X1_145 BUFX4_130/Y BUFX4_193/Y gnd MUX2X1_94/S vdd NOR2X1
XMUX2X1_84 INVX1_97/Y MUX2X1_39/B MUX2X1_84/S gnd MUX2X1_84/Y vdd MUX2X1
XMUX2X1_73 INVX1_83/Y MUX2X1_61/B MUX2X1_71/S gnd MUX2X1_73/Y vdd MUX2X1
XNOR2X1_156 MUX2X1_247/B NOR2X1_155/B gnd AOI21X1_93/C vdd NOR2X1
XNOR2X1_189 NOR2X1_514/A NOR2X1_188/B gnd NOR2X1_189/Y vdd NOR2X1
XNOR2X1_178 NOR2X1_178/A MUX2X1_108/S gnd NOR2X1_178/Y vdd NOR2X1
XOAI21X1_618 AOI21X1_286/Y AOI21X1_287/Y BUFX4_410/Y gnd OAI21X1_618/Y vdd OAI21X1
XOAI21X1_607 INVX1_262/Y BUFX4_274/Y NAND2X1_183/Y gnd MUX2X1_183/B vdd OAI21X1
XOAI21X1_629 INVX1_275/Y BUFX4_226/Y OAI21X1_629/C gnd MUX2X1_189/B vdd OAI21X1
XDFFPOSX1_521 INVX1_384/A CLKBUF1_57/Y MUX2X1_387/Y gnd vdd DFFPOSX1
XMUX2X1_129 BUFX4_180/Y INVX1_142/Y NOR2X1_233/Y gnd MUX2X1_129/Y vdd MUX2X1
XDFFPOSX1_510 NOR2X1_564/A CLKBUF1_18/Y AOI21X1_610/Y gnd vdd DFFPOSX1
XDFFPOSX1_532 INVX1_324/A CLKBUF1_64/Y MUX2X1_390/Y gnd vdd DFFPOSX1
XMUX2X1_107 MUX2X1_44/A INVX1_120/Y MUX2X1_108/S gnd MUX2X1_107/Y vdd MUX2X1
XMUX2X1_118 MUX2X1_59/B INVX1_131/Y NOR2X1_707/B gnd MUX2X1_118/Y vdd MUX2X1
XDFFPOSX1_543 INVX1_262/A CLKBUF1_92/Y DFFPOSX1_543/D gnd vdd DFFPOSX1
XDFFPOSX1_565 NOR2X1_735/A CLKBUF1_14/Y AOI21X1_623/Y gnd vdd DFFPOSX1
XDFFPOSX1_554 INVX1_439/A CLKBUF1_42/Y MUX2X1_397/Y gnd vdd DFFPOSX1
XDFFPOSX1_587 OAI21X1_617/B CLKBUF1_53/Y DFFPOSX1_587/D gnd vdd DFFPOSX1
XDFFPOSX1_576 INVX1_328/A CLKBUF1_94/Y MUX2X1_405/Y gnd vdd DFFPOSX1
XDFFPOSX1_598 INVX1_7/A CLKBUF1_76/Y MUX2X1_4/Y gnd vdd DFFPOSX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XNOR2X1_690 NOR2X1_690/A NOR2X1_167/B gnd NOR2X1_690/Y vdd NOR2X1
XAOI21X1_270 BUFX4_257/Y INVX1_249/Y AOI21X1_270/C gnd AOI21X1_270/Y vdd AOI21X1
XAOI21X1_292 BUFX4_202/Y AOI21X1_292/B AOI21X1_288/Y gnd MUX2X1_190/A vdd AOI21X1
XAOI21X1_281 BUFX4_271/Y OAI21X1_605/Y BUFX4_418/Y gnd AOI21X1_281/Y vdd AOI21X1
XFILL_47_2_1 gnd vdd FILL
XFILL_30_1_1 gnd vdd FILL
XDFFPOSX1_1050 NOR2X1_249/A CLKBUF1_64/Y AOI21X1_159/Y gnd vdd DFFPOSX1
XFILL_38_2_1 gnd vdd FILL
XFILL_50_9_0 gnd vdd FILL
XOAI21X1_404 NAND2X1_24/Y BUFX4_468/Y OAI21X1_404/C gnd OAI21X1_404/Y vdd OAI21X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_437 traffic_Street_1[0] traffic_Street_1[1] traffic_Street_1[2] gnd AND2X2_3/A
+ vdd OAI21X1
XOAI21X1_426 OAI21X1_54/A MUX2X1_61/B OAI21X1_425/Y gnd OAI21X1_426/Y vdd OAI21X1
XOAI21X1_448 traffic_Street_0[0] traffic_Street_0[1] traffic_Street_0[2] gnd AND2X2_6/A
+ vdd OAI21X1
XOAI21X1_415 BUFX4_62/Y BUFX4_460/Y AND2X2_36/A gnd OAI21X1_415/Y vdd OAI21X1
XOAI21X1_459 AND2X2_4/Y traffic_Street_0[2] traffic_Street_0[3] gnd OAI21X1_473/B
+ vdd OAI21X1
XDFFPOSX1_340 NOR2X1_657/A CLKBUF1_100/Y AOI21X1_545/Y gnd vdd DFFPOSX1
XDFFPOSX1_362 INVX1_229/A CLKBUF1_27/Y MUX2X1_301/Y gnd vdd DFFPOSX1
XDFFPOSX1_373 NOR2X1_652/A CLKBUF1_102/Y AOI21X1_540/Y gnd vdd DFFPOSX1
XDFFPOSX1_351 INVX1_296/A CLKBUF1_47/Y MUX2X1_310/Y gnd vdd DFFPOSX1
XDFFPOSX1_395 BUFX2_4/A CLKBUF1_59/Y INVX4_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_384 NOR2X1_634/A CLKBUF1_76/Y AOI21X1_522/Y gnd vdd DFFPOSX1
XFILL_4_2_1 gnd vdd FILL
XFILL_29_2_1 gnd vdd FILL
XFILL_41_9_0 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_960 BUFX4_340/Y NOR2X1_705/A BUFX4_147/Y gnd AOI21X1_418/C vdd OAI21X1
XOAI21X1_971 INVX1_389/Y BUFX4_227/Y OAI21X1_971/C gnd MUX2X1_239/B vdd OAI21X1
XOAI21X1_982 OAI21X1_14/C BUFX4_84/Y AOI21X1_430/Y gnd OAI21X1_982/Y vdd OAI21X1
XOAI21X1_993 NOR2X1_491/Y OAI21X1_987/Y OAI21X1_993/C gnd OAI21X1_993/Y vdd OAI21X1
XOAI21X1_20 OAI21X1_24/A MUX2X1_1/B OAI21X1_19/Y gnd OAI21X1_20/Y vdd OAI21X1
XFILL_32_9_0 gnd vdd FILL
XOAI21X1_31 BUFX4_125/Y BUFX4_292/Y OAI21X1_31/C gnd OAI21X1_32/C vdd OAI21X1
XOAI21X1_53 INVX4_4/A BUFX4_464/Y NOR2X1_440/A gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_42 OAI21X1_40/A BUFX4_316/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_86 NAND2X1_32/Y BUFX4_173/Y OAI21X1_85/Y gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_75 BUFX4_448/Y BUFX4_43/Y NOR2X1_403/A gnd OAI21X1_76/C vdd OAI21X1
XOAI21X1_64 BUFX4_69/Y OAI21X1_64/B OAI21X1_63/Y gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_97 BUFX4_120/Y BUFX4_476/Y AND2X2_45/A gnd OAI21X1_98/C vdd OAI21X1
XFILL_23_9_0 gnd vdd FILL
XOAI21X1_212 BUFX4_452/Y BUFX4_404/Y MUX2X1_246/A gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_201 BUFX4_216/Y NAND2X1_60/Y OAI21X1_201/C gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_256 BUFX4_126/Y BUFX4_432/Y NAND2X1_210/A gnd OAI21X1_256/Y vdd OAI21X1
XOAI21X1_245 BUFX4_377/Y NAND2X1_68/Y OAI21X1_244/Y gnd OAI21X1_245/Y vdd OAI21X1
XOAI21X1_223 NAND2X1_62/Y AND2X2_3/B OAI21X1_222/Y gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_234 BUFX4_123/Y BUFX4_138/Y AND2X2_33/A gnd OAI21X1_235/C vdd OAI21X1
XOAI21X1_289 NAND2X1_75/Y BUFX4_218/Y OAI21X1_288/Y gnd OAI21X1_289/Y vdd OAI21X1
XOAI21X1_267 NAND2X1_72/Y BUFX4_174/Y OAI21X1_267/C gnd OAI21X1_267/Y vdd OAI21X1
XOAI21X1_278 BUFX4_135/Y BUFX4_163/Y OAI21X1_278/C gnd OAI21X1_279/C vdd OAI21X1
XAND2X2_12 AND2X2_12/A OR2X2_6/Y gnd AND2X2_12/Y vdd AND2X2
XINVX1_309 INVX1_309/A gnd INVX1_309/Y vdd INVX1
XAND2X2_45 AND2X2_45/A AND2X2_32/B gnd AND2X2_45/Y vdd AND2X2
XAND2X2_34 BUFX4_34/Y AND2X2_34/B gnd AND2X2_34/Y vdd AND2X2
XAND2X2_23 AND2X2_23/A AND2X2_23/B gnd AND2X2_23/Y vdd AND2X2
XDFFPOSX1_181 INVX1_447/A CLKBUF1_27/Y MUX2X1_278/Y gnd vdd DFFPOSX1
XDFFPOSX1_170 INVX1_226/A CLKBUF1_23/Y MUX2X1_288/Y gnd vdd DFFPOSX1
XDFFPOSX1_192 INVX1_364/A CLKBUF1_83/Y MUX2X1_292/Y gnd vdd DFFPOSX1
XNAND2X1_262 INVX8_28/A OAI22X1_28/Y gnd AOI21X1_388/B vdd NAND2X1
XNAND2X1_251 BUFX4_38/Y MUX2X1_219/Y gnd AOI22X1_21/A vdd NAND2X1
XNAND2X1_240 BUFX4_291/Y NOR2X1_702/A gnd NAND2X1_240/Y vdd NAND2X1
XNAND2X1_284 BUFX4_275/Y INVX1_457/A gnd NAND2X1_284/Y vdd NAND2X1
XNAND2X1_295 BUFX4_34/Y MUX2X1_239/Y gnd AOI22X1_27/A vdd NAND2X1
XNAND2X1_273 BUFX4_410/Y MUX2X1_228/Y gnd NAND2X1_276/A vdd NAND2X1
XFILL_44_0_1 gnd vdd FILL
XFILL_14_9_0 gnd vdd FILL
XOAI21X1_1508 BUFX4_429/Y NAND2X1_77/Y OAI21X1_1508/C gnd DFFPOSX1_516/D vdd OAI21X1
XOAI21X1_1519 BUFX4_310/Y BUFX4_300/Y NAND2X1_340/A gnd OAI21X1_1520/C vdd OAI21X1
XOAI21X1_790 BUFX4_336/Y INVX1_324/Y NAND2X1_244/Y gnd OAI21X1_790/Y vdd OAI21X1
XMUX2X1_290 INVX1_227/Y BUFX4_443/Y MUX2X1_51/S gnd MUX2X1_290/Y vdd MUX2X1
XFILL_48_2 gnd vdd FILL
XFILL_35_0_1 gnd vdd FILL
XCLKBUF1_10 BUFX4_9/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XCLKBUF1_32 BUFX4_6/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_21 BUFX4_7/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_43 BUFX4_1/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XCLKBUF1_54 BUFX4_9/Y gnd CLKBUF1_54/Y vdd CLKBUF1
XCLKBUF1_65 BUFX4_9/Y gnd CLKBUF1_65/Y vdd CLKBUF1
XCLKBUF1_76 BUFX4_7/Y gnd CLKBUF1_76/Y vdd CLKBUF1
XCLKBUF1_98 BUFX4_3/Y gnd CLKBUF1_98/Y vdd CLKBUF1
XCLKBUF1_87 BUFX4_3/Y gnd CLKBUF1_87/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_26_0_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XBUFX4_404 INVX8_21/Y gnd BUFX4_404/Y vdd BUFX4
XBUFX4_426 INVX8_3/Y gnd BUFX4_426/Y vdd BUFX4
XBUFX4_415 address[2] gnd BUFX4_415/Y vdd BUFX4
XBUFX4_437 INVX8_2/Y gnd BUFX4_437/Y vdd BUFX4
XFILL_46_8_0 gnd vdd FILL
XBUFX4_448 BUFX4_449/A gnd BUFX4_448/Y vdd BUFX4
XBUFX4_459 INVX8_25/Y gnd BUFX4_459/Y vdd BUFX4
XNOR2X1_508 NOR2X1_508/A NOR2X1_508/B gnd NOR2X1_508/Y vdd NOR2X1
XFILL_17_0_1 gnd vdd FILL
XNOR2X1_519 BUFX4_204/Y NOR2X1_519/B gnd OAI22X1_48/D vdd NOR2X1
XOAI21X1_1305 BUFX4_318/Y NAND2X1_37/Y OAI21X1_1305/C gnd OAI21X1_1305/Y vdd OAI21X1
XDFFPOSX1_906 NOR2X1_589/A CLKBUF1_101/Y AOI21X1_102/Y gnd vdd DFFPOSX1
XOAI21X1_1327 BUFX4_57/Y BUFX4_398/Y NAND2X1_274/B gnd OAI21X1_1328/C vdd OAI21X1
XOAI21X1_1316 INVX4_4/A BUFX4_52/Y NOR2X1_414/B gnd OAI21X1_1316/Y vdd OAI21X1
XOAI21X1_1338 BUFX4_123/Y BUFX4_396/Y OAI21X1_1096/B gnd OAI21X1_1338/Y vdd OAI21X1
XDFFPOSX1_928 NOR2X1_179/A CLKBUF1_41/Y AOI21X1_110/Y gnd vdd DFFPOSX1
XDFFPOSX1_939 INVX1_123/A CLKBUF1_61/Y MUX2X1_110/Y gnd vdd DFFPOSX1
XOAI21X1_1349 BUFX4_318/Y NAND2X1_51/Y OAI21X1_1348/Y gnd DFFPOSX1_325/D vdd OAI21X1
XDFFPOSX1_917 AND2X2_42/A CLKBUF1_39/Y OAI21X1_229/Y gnd vdd DFFPOSX1
XFILL_37_8_0 gnd vdd FILL
XAOI21X1_600 MUX2X1_27/B MUX2X1_120/S NOR2X1_712/Y gnd AOI21X1_600/Y vdd AOI21X1
XAOI21X1_622 MUX2X1_4/B MUX2X1_400/S NOR2X1_734/Y gnd AOI21X1_622/Y vdd AOI21X1
XAOI21X1_611 BUFX4_439/Y NOR2X1_234/Y NOR2X1_723/Y gnd AOI21X1_611/Y vdd AOI21X1
XFILL_20_7_0 gnd vdd FILL
XINVX4_14 address[6] gnd INVX4_14/Y vdd INVX4
XFILL_3_8_0 gnd vdd FILL
XFILL_28_8_0 gnd vdd FILL
XFILL_11_7_0 gnd vdd FILL
XBUFX4_201 address[3] gnd BUFX4_201/Y vdd BUFX4
XBUFX4_212 INVX8_11/Y gnd MUX2X1_71/B vdd BUFX4
XFILL_19_8_0 gnd vdd FILL
XBUFX4_234 BUFX4_18/Y gnd BUFX4_234/Y vdd BUFX4
XBUFX4_245 BUFX4_17/Y gnd AND2X2_52/A vdd BUFX4
XBUFX4_223 BUFX4_17/Y gnd BUFX4_223/Y vdd BUFX4
XBUFX4_278 BUFX4_18/Y gnd BUFX4_278/Y vdd BUFX4
XBUFX4_256 BUFX4_20/Y gnd BUFX4_256/Y vdd BUFX4
XBUFX4_267 BUFX4_20/Y gnd AND2X2_29/A vdd BUFX4
XBUFX4_289 BUFX4_17/Y gnd BUFX4_289/Y vdd BUFX4
XNOR2X1_305 BUFX4_320/Y NOR2X1_351/B gnd INVX1_190/A vdd NOR2X1
XNOR2X1_316 INVX2_18/A INVX2_19/Y gnd NOR2X1_316/Y vdd NOR2X1
XNOR2X1_349 NOR2X1_349/A NOR2X1_349/B gnd NAND3X1_68/B vdd NOR2X1
XNOR2X1_338 INVX4_12/A NAND3X1_65/C gnd NOR2X1_338/Y vdd NOR2X1
XNOR2X1_327 OAI22X1_1/Y NOR2X1_327/B gnd NOR2X1_327/Y vdd NOR2X1
XOAI21X1_1113 BUFX4_342/Y NOR2X1_686/A BUFX4_148/Y gnd OAI22X1_53/C vdd OAI21X1
XOAI21X1_1102 NOR2X1_530/Y OAI21X1_1102/B OAI21X1_1102/C gnd OAI21X1_1103/A vdd OAI21X1
XOAI21X1_1135 OAI21X1_1134/Y BUFX4_41/Y BUFX4_169/Y gnd OAI22X1_63/C vdd OAI21X1
XOAI21X1_1124 BUFX4_220/Y NOR2X1_677/A BUFX4_103/Y gnd OAI22X1_58/B vdd OAI21X1
XDFFPOSX1_703 NOR2X1_66/A CLKBUF1_24/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_714 NOR2X1_72/A CLKBUF1_80/Y AOI21X1_37/Y gnd vdd DFFPOSX1
XOAI21X1_1146 OAI22X1_64/Y BUFX4_36/Y BUFX4_169/Y gnd OAI22X1_65/B vdd OAI21X1
XOAI21X1_1179 OAI21X1_99/C BUFX4_261/Y BUFX4_82/Y gnd OAI21X1_1180/B vdd OAI21X1
XDFFPOSX1_736 INVX1_59/A CLKBUF1_11/Y MUX2X1_49/Y gnd vdd DFFPOSX1
XOAI21X1_1168 NOR2X1_564/Y NOR2X1_565/Y BUFX4_252/Y gnd AOI21X1_489/A vdd OAI21X1
XDFFPOSX1_725 INVX1_54/A CLKBUF1_12/Y MUX2X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_747 INVX1_61/A CLKBUF1_46/Y MUX2X1_51/Y gnd vdd DFFPOSX1
XOAI21X1_1157 BUFX4_241/Y OAI21X1_1157/B BUFX4_115/Y gnd AOI21X1_486/C vdd OAI21X1
XDFFPOSX1_769 NOR2X1_99/A CLKBUF1_20/Y AOI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_758 INVX1_68/A CLKBUF1_1/Y MUX2X1_58/Y gnd vdd DFFPOSX1
XAOI21X1_452 INVX1_165/Y BUFX4_349/Y AOI21X1_452/C gnd AOI21X1_452/Y vdd AOI21X1
XAOI21X1_430 BUFX4_83/Y INVX1_30/Y BUFX4_236/Y gnd AOI21X1_430/Y vdd AOI21X1
XAOI21X1_441 BUFX4_414/Y AOI21X1_441/B BUFX4_167/Y gnd AOI22X1_29/B vdd AOI21X1
XAOI21X1_485 BUFX4_362/Y INVX1_429/Y AOI21X1_485/C gnd AOI21X1_485/Y vdd AOI21X1
XAOI21X1_463 INVX1_447/A BUFX4_151/Y BUFX4_344/Y gnd AOI21X1_463/Y vdd AOI21X1
XAOI21X1_474 BUFX4_281/Y INVX1_421/Y BUFX4_97/Y gnd AOI21X1_474/Y vdd AOI21X1
XAOI21X1_496 NOR2X1_83/A AND2X2_25/B AOI21X1_496/C gnd AOI21X1_496/Y vdd AOI21X1
XNAND3X1_12 INVX2_14/Y NAND3X1_12/B OR2X2_2/Y gnd NAND3X1_13/B vdd NAND3X1
XNAND3X1_23 BUFX2_3/A NAND3X1_23/B NAND3X1_23/C gnd NOR3X1_5/C vdd NAND3X1
XNAND3X1_56 NAND3X1_56/A XNOR2X1_4/Y NAND3X1_56/C gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_45 AOI22X1_6/B INVX1_203/Y NOR3X1_7/Y gnd AOI22X1_6/D vdd NAND3X1
XNAND3X1_34 INVX4_7/A NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_34/Y vdd NAND3X1
XNAND3X1_67 police_Interrupt INVX4_9/A AND2X2_18/A gnd XNOR2X1_7/A vdd NAND3X1
XNAND3X1_78 BUFX4_41/Y NAND3X1_78/B NAND3X1_78/C gnd NAND3X1_78/Y vdd NAND3X1
XNOR2X1_12 NOR2X1_2/A INVX1_23/Y gnd NOR2X1_12/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A AOI21X1_7/B gnd AOI21X1_5/C vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_33/Y gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_45 NOR2X1_45/A NOR2X1_47/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_56 NOR2X1_56/A NOR2X1_54/Y gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_65/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A MUX2X1_45/S gnd NOR2X1_78/Y vdd NOR2X1
XFILL_43_6_0 gnd vdd FILL
XNOR2X1_89 INVX2_9/Y INVX2_7/Y gnd INVX8_17/A vdd NOR2X1
XMUX2X1_63 INVX1_73/Y MUX2X1_59/B MUX2X1_66/S gnd MUX2X1_63/Y vdd MUX2X1
XNOR2X1_124 NOR2X1_124/A MUX2X1_320/S gnd AOI21X1_71/C vdd NOR2X1
XMUX2X1_30 MUX2X1_9/B INVX1_38/Y MUX2X1_31/S gnd MUX2X1_30/Y vdd MUX2X1
XNOR2X1_102 BUFX4_395/Y BUFX4_144/Y gnd MUX2X1_75/S vdd NOR2X1
XNOR2X1_113 NOR2X1_113/A AOI21X1_62/B gnd NOR2X1_113/Y vdd NOR2X1
XMUX2X1_41 INVX1_51/Y MUX2X1_44/A MUX2X1_42/S gnd MUX2X1_41/Y vdd MUX2X1
XMUX2X1_52 INVX1_62/Y MUX2X1_64/B MUX2X1_51/S gnd MUX2X1_52/Y vdd MUX2X1
XMUX2X1_96 MUX2X1_96/A INVX1_109/Y MUX2X1_96/S gnd MUX2X1_96/Y vdd MUX2X1
XNOR2X1_135 BUFX4_131/Y BUFX4_144/Y gnd NOR2X1_137/B vdd NOR2X1
XNOR2X1_146 NOR2X1_146/A MUX2X1_94/S gnd AOI21X1_86/C vdd NOR2X1
XMUX2X1_85 INVX1_98/Y BUFX4_176/Y MUX2X1_84/S gnd MUX2X1_85/Y vdd MUX2X1
XFILL_34_6_0 gnd vdd FILL
XMUX2X1_74 INVX1_84/Y MUX2X1_58/A MUX2X1_71/S gnd MUX2X1_74/Y vdd MUX2X1
XNOR2X1_157 NOR2X1_157/A NOR2X1_155/B gnd AOI21X1_94/C vdd NOR2X1
XNOR2X1_179 NOR2X1_179/A MUX2X1_108/S gnd NOR2X1_179/Y vdd NOR2X1
XNOR2X1_168 INVX2_11/Y INVX2_8/Y gnd INVX8_22/A vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XOAI21X1_619 INVX1_22/Y BUFX4_287/Y BUFX4_106/Y gnd OAI21X1_619/Y vdd OAI21X1
XOAI21X1_608 INVX1_263/Y BUFX4_276/Y OAI21X1_608/C gnd MUX2X1_183/A vdd OAI21X1
XMUX2X1_108 BUFX4_466/Y INVX1_121/Y MUX2X1_108/S gnd MUX2X1_108/Y vdd MUX2X1
XDFFPOSX1_511 INVX1_266/A CLKBUF1_32/Y MUX2X1_381/Y gnd vdd DFFPOSX1
XDFFPOSX1_522 INVX1_437/A CLKBUF1_52/Y MUX2X1_388/Y gnd vdd DFFPOSX1
XDFFPOSX1_500 NOR2X1_716/A CLKBUF1_89/Y AOI21X1_604/Y gnd vdd DFFPOSX1
XMUX2X1_119 BUFX4_371/Y INVX1_132/Y NOR2X1_707/B gnd MUX2X1_119/Y vdd MUX2X1
XDFFPOSX1_544 INVX1_322/A CLKBUF1_90/Y DFFPOSX1_544/D gnd vdd DFFPOSX1
XDFFPOSX1_555 NAND2X1_184/B CLKBUF1_23/Y DFFPOSX1_555/D gnd vdd DFFPOSX1
XDFFPOSX1_533 NOR2X1_727/A CLKBUF1_67/Y AOI21X1_615/Y gnd vdd DFFPOSX1
XDFFPOSX1_588 OAI21X1_797/B CLKBUF1_35/Y OAI21X1_1564/Y gnd vdd DFFPOSX1
XDFFPOSX1_599 NAND2X1_5/A CLKBUF1_84/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_566 INVX1_424/A CLKBUF1_72/Y MUX2X1_403/Y gnd vdd DFFPOSX1
XDFFPOSX1_577 INVX1_460/A CLKBUF1_11/Y MUX2X1_406/Y gnd vdd DFFPOSX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XFILL_0_6_0 gnd vdd FILL
XFILL_25_6_0 gnd vdd FILL
XNOR2X1_680 NOR2X1_680/A MUX2X1_94/S gnd NOR2X1_680/Y vdd NOR2X1
XNOR2X1_691 NOR2X1_691/A NOR2X1_167/B gnd NOR2X1_691/Y vdd NOR2X1
XAOI21X1_260 BUFX4_242/Y NOR2X1_694/A AOI21X1_260/C gnd OAI22X1_4/B vdd AOI21X1
XAOI21X1_293 BUFX4_412/Y MUX2X1_188/Y AND2X2_48/B gnd AOI22X1_16/B vdd AOI21X1
XAOI21X1_271 BUFX4_153/Y OAI21X1_589/Y AOI21X1_270/Y gnd AOI21X1_271/Y vdd AOI21X1
XAOI21X1_282 BUFX4_419/Y MUX2X1_183/Y BUFX4_165/Y gnd AOI22X1_15/A vdd AOI21X1
XFILL_8_7_0 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XDFFPOSX1_1051 INVX1_282/A CLKBUF1_52/Y OAI21X1_329/Y gnd vdd DFFPOSX1
XDFFPOSX1_1040 AND2X2_37/A CLKBUF1_42/Y AOI21X1_153/Y gnd vdd DFFPOSX1
XFILL_50_9_1 gnd vdd FILL
XOAI21X1_405 BUFX4_460/Y BUFX4_303/Y NOR2X1_379/A gnd OAI21X1_406/C vdd OAI21X1
XOAI21X1_438 NOR2X1_299/Y AND2X2_1/Y AOI21X1_212/B gnd AOI22X1_1/C vdd OAI21X1
XOAI21X1_427 INVX4_4/A BUFX4_462/Y NOR2X1_610/A gnd OAI21X1_427/Y vdd OAI21X1
XOAI21X1_416 BUFX4_177/Y OAI21X1_48/B OAI21X1_415/Y gnd OAI21X1_416/Y vdd OAI21X1
XOAI21X1_449 traffic_Street_0[1] traffic_Street_0[2] traffic_Street_0[3] gnd INVX2_15/A
+ vdd OAI21X1
XDFFPOSX1_330 AND2X2_22/B CLKBUF1_100/Y AOI21X1_546/Y gnd vdd DFFPOSX1
XDFFPOSX1_352 INVX1_345/A CLKBUF1_78/Y MUX2X1_311/Y gnd vdd DFFPOSX1
XDFFPOSX1_363 INVX1_293/A CLKBUF1_20/Y MUX2X1_302/Y gnd vdd DFFPOSX1
XDFFPOSX1_374 NOR2X1_367/B CLKBUF1_22/Y DFFPOSX1_374/D gnd vdd DFFPOSX1
XDFFPOSX1_341 INVX1_415/A CLKBUF1_46/Y OAI21X1_1331/Y gnd vdd DFFPOSX1
XDFFPOSX1_385 NOR2X1_635/A CLKBUF1_28/Y AOI21X1_523/Y gnd vdd DFFPOSX1
XDFFPOSX1_396 NOR2X1_625/A CLKBUF1_43/Y AOI21X1_513/Y gnd vdd DFFPOSX1
XFILL_41_9_1 gnd vdd FILL
XFILL_40_4_0 gnd vdd FILL
XOAI21X1_950 AOI22X1_25/Y AND2X2_48/B INVX4_14/Y gnd OAI22X1_42/B vdd OAI21X1
XOAI21X1_961 BUFX4_284/Y OAI21X1_961/B BUFX4_117/Y gnd AOI21X1_419/C vdd OAI21X1
XOAI21X1_972 INVX1_390/Y BUFX4_229/Y NAND2X1_294/Y gnd MUX2X1_239/A vdd OAI21X1
XOAI21X1_983 BUFX4_149/Y NOR2X1_25/A BUFX4_237/Y gnd OAI21X1_984/B vdd OAI21X1
XOAI21X1_994 BUFX4_49/Y AOI22X1_27/Y NAND2X1_300/Y gnd AOI22X1_28/C vdd OAI21X1
XFILL_48_5_0 gnd vdd FILL
XOAI21X1_10 BUFX4_292/Y BUFX4_303/Y INVX1_272/A gnd OAI21X1_11/C vdd OAI21X1
XFILL_32_9_1 gnd vdd FILL
XOAI21X1_54 OAI21X1_54/A MUX2X1_27/B OAI21X1_53/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_32 NAND2X1_24/Y BUFX4_64/Y OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_21 BUFX4_450/Y BUFX4_292/Y NOR2X1_443/A gnd OAI21X1_22/C vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XOAI21X1_43 BUFX4_62/Y BUFX4_460/Y OAI21X1_43/C gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_87 BUFX4_124/Y BUFX4_45/Y OAI21X1_87/C gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_76 NAND2X1_31/Y BUFX4_213/Y OAI21X1_76/C gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_65 BUFX4_190/Y BUFX4_464/Y OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_98 NAND2X1_36/Y BUFX4_381/Y OAI21X1_98/C gnd OAI21X1_98/Y vdd OAI21X1
XFILL_39_5_0 gnd vdd FILL
XFILL_23_9_1 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_213 NAND2X1_61/Y MUX2X1_57/A OAI21X1_212/Y gnd OAI21X1_213/Y vdd OAI21X1
XOAI21X1_202 BUFX4_143/Y BUFX4_407/Y INVX1_335/A gnd OAI21X1_203/C vdd OAI21X1
XOAI21X1_246 BUFX4_60/Y BUFX4_432/Y OAI21X1_246/C gnd OAI21X1_246/Y vdd OAI21X1
XOAI21X1_224 BUFX4_383/Y BUFX4_139/Y OAI21X1_696/A gnd OAI21X1_224/Y vdd OAI21X1
XOAI21X1_235 NAND2X1_66/Y MUX2X1_96/A OAI21X1_235/C gnd OAI21X1_235/Y vdd OAI21X1
XOAI21X1_257 NAND2X1_70/Y MUX2X1_59/B OAI21X1_256/Y gnd OAI21X1_257/Y vdd OAI21X1
XOAI21X1_268 BUFX4_451/Y BUFX4_164/Y INVX1_405/A gnd OAI21X1_269/C vdd OAI21X1
XOAI21X1_279 BUFX4_465/Y NAND2X1_73/Y OAI21X1_279/C gnd OAI21X1_279/Y vdd OAI21X1
XAND2X2_13 AND2X2_13/A XOR2X1_2/B gnd AND2X2_13/Y vdd AND2X2
XAND2X2_24 BUFX4_36/Y AND2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XAND2X2_35 AND2X2_35/A BUFX4_414/Y gnd AND2X2_35/Y vdd AND2X2
XAND2X2_46 AND2X2_46/A AND2X2_46/B gnd AND2X2_46/Y vdd AND2X2
XDFFPOSX1_171 NOR2X1_643/A CLKBUF1_57/Y AOI21X1_531/Y gnd vdd DFFPOSX1
XDFFPOSX1_182 NAND2X1_172/B CLKBUF1_65/Y DFFPOSX1_182/D gnd vdd DFFPOSX1
XDFFPOSX1_160 INVX1_356/A CLKBUF1_22/Y MUX2X1_347/Y gnd vdd DFFPOSX1
XDFFPOSX1_193 INVX1_448/A CLKBUF1_15/Y MUX2X1_293/Y gnd vdd DFFPOSX1
XNAND2X1_230 BUFX4_205/Y NAND2X1_230/B gnd AOI21X1_325/C vdd NAND2X1
XNAND2X1_252 NOR2X1_98/A BUFX4_259/Y gnd OAI21X1_835/C vdd NAND2X1
XNAND2X1_241 BUFX4_166/Y MUX2X1_213/Y gnd OAI21X1_782/C vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XNAND2X1_263 BUFX4_34/Y OAI22X1_29/Y gnd NAND2X1_263/Y vdd NAND2X1
XNAND2X1_274 BUFX4_249/Y NAND2X1_274/B gnd NAND2X1_274/Y vdd NAND2X1
XNAND2X1_285 BUFX4_391/Y NAND2X1_285/B gnd AOI22X1_28/A vdd NAND2X1
XNAND2X1_296 NOR2X1_47/A BUFX4_240/Y gnd OAI21X1_988/C vdd NAND2X1
XFILL_14_9_1 gnd vdd FILL
XFILL_13_4_0 gnd vdd FILL
XOAI21X1_1509 BUFX4_132/Y BUFX4_459/Y NAND2X1_286/B gnd OAI21X1_1510/C vdd OAI21X1
XOAI21X1_791 BUFX4_234/Y OAI21X1_791/B BUFX4_85/Y gnd AOI21X1_344/C vdd OAI21X1
XOAI21X1_780 NOR2X1_431/Y OAI21X1_779/Y OAI21X1_778/Y gnd OAI21X1_780/Y vdd OAI21X1
XMUX2X1_280 BUFX4_430/Y INVX1_302/Y MUX2X1_45/S gnd MUX2X1_280/Y vdd MUX2X1
XMUX2X1_291 INVX1_291/Y BUFX4_430/Y MUX2X1_51/S gnd MUX2X1_291/Y vdd MUX2X1
XFILL_48_3 gnd vdd FILL
XCLKBUF1_11 BUFX4_2/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XCLKBUF1_22 BUFX4_9/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_33 BUFX4_4/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_66 BUFX4_3/Y gnd CLKBUF1_66/Y vdd CLKBUF1
XCLKBUF1_55 BUFX4_3/Y gnd CLKBUF1_55/Y vdd CLKBUF1
XCLKBUF1_44 BUFX4_4/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XCLKBUF1_88 BUFX4_10/Y gnd CLKBUF1_88/Y vdd CLKBUF1
XCLKBUF1_99 BUFX4_3/Y gnd CLKBUF1_99/Y vdd CLKBUF1
XCLKBUF1_77 BUFX4_3/Y gnd CLKBUF1_77/Y vdd CLKBUF1
XINVX1_107 INVX1_107/A gnd MUX2X1_94/B vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XBUFX4_438 INVX8_2/Y gnd MUX2X1_1/B vdd BUFX4
XBUFX4_427 INVX8_3/Y gnd MUX2X1_18/B vdd BUFX4
XBUFX4_416 address[2] gnd BUFX4_416/Y vdd BUFX4
XBUFX4_405 INVX8_21/Y gnd BUFX4_405/Y vdd BUFX4
XFILL_46_8_1 gnd vdd FILL
XBUFX4_449 BUFX4_449/A gnd BUFX4_449/Y vdd BUFX4
XFILL_45_3_0 gnd vdd FILL
XNOR2X1_509 NOR2X1_509/A BUFX4_225/Y gnd NOR2X1_509/Y vdd NOR2X1
XOAI21X1_1328 BUFX4_69/Y NAND2X1_44/Y OAI21X1_1328/C gnd DFFPOSX1_356/D vdd OAI21X1
XOAI21X1_1317 NAND2X1_40/Y MUX2X1_27/B OAI21X1_1316/Y gnd DFFPOSX1_375/D vdd OAI21X1
XOAI21X1_1306 BUFX4_61/Y BUFX4_52/Y NAND2X1_172/B gnd OAI21X1_1307/C vdd OAI21X1
XDFFPOSX1_907 INVX1_110/A CLKBUF1_29/Y MUX2X1_97/Y gnd vdd DFFPOSX1
XOAI21X1_1339 NAND2X1_48/Y BUFX4_316/Y OAI21X1_1338/Y gnd OAI21X1_1339/Y vdd OAI21X1
XDFFPOSX1_929 INVX1_120/A CLKBUF1_54/Y MUX2X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_918 INVX1_442/A CLKBUF1_29/Y OAI21X1_231/Y gnd vdd DFFPOSX1
XFILL_37_8_1 gnd vdd FILL
XFILL_36_3_0 gnd vdd FILL
XAOI21X1_601 MUX2X1_27/B MUX2X1_376/S NOR2X1_713/Y gnd AOI21X1_601/Y vdd AOI21X1
XAOI21X1_612 BUFX4_424/Y NOR2X1_234/Y NOR2X1_724/Y gnd AOI21X1_612/Y vdd AOI21X1
XAOI21X1_623 BUFX4_63/Y NOR2X1_261/B NOR2X1_735/Y gnd AOI21X1_623/Y vdd AOI21X1
XFILL_20_7_1 gnd vdd FILL
XFILL_3_8_1 gnd vdd FILL
XFILL_28_8_1 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XBUFX4_202 address[3] gnd BUFX4_202/Y vdd BUFX4
XBUFX4_246 BUFX4_21/Y gnd BUFX4_246/Y vdd BUFX4
XBUFX4_213 INVX8_11/Y gnd BUFX4_213/Y vdd BUFX4
XBUFX4_235 BUFX4_23/Y gnd BUFX4_235/Y vdd BUFX4
XFILL_19_8_1 gnd vdd FILL
XBUFX4_224 BUFX4_22/Y gnd BUFX4_224/Y vdd BUFX4
XBUFX4_257 BUFX4_21/Y gnd BUFX4_257/Y vdd BUFX4
XFILL_18_3_0 gnd vdd FILL
XBUFX4_279 BUFX4_23/Y gnd AND2X2_41/A vdd BUFX4
XBUFX4_268 BUFX4_22/Y gnd BUFX4_268/Y vdd BUFX4
XNOR2X1_306 AND2X2_5/B AND2X2_5/A gnd NOR2X1_306/Y vdd NOR2X1
XNOR2X1_328 INVX2_22/A XOR2X1_3/A gnd NOR2X1_328/Y vdd NOR2X1
XNOR2X1_339 AND2X2_6/B AND2X2_6/A gnd NOR2X1_339/Y vdd NOR2X1
XNOR2X1_317 INVX1_201/A NOR2X1_316/Y gnd AND2X2_8/B vdd NOR2X1
XOAI21X1_1103 OAI21X1_1103/A BUFX4_33/Y BUFX4_166/Y gnd OAI22X1_52/B vdd OAI21X1
XOAI21X1_1125 BUFX4_354/Y NOR2X1_674/A AOI21X1_477/Y gnd OAI21X1_1125/Y vdd OAI21X1
XDFFPOSX1_704 NOR2X1_67/A CLKBUF1_80/Y AOI21X1_33/Y gnd vdd DFFPOSX1
XOAI21X1_1136 BUFX4_333/Y INVX1_7/A BUFX4_146/Y gnd OAI22X1_61/C vdd OAI21X1
XOAI21X1_1147 INVX1_426/Y BUFX4_235/Y NAND2X1_335/Y gnd MUX2X1_257/B vdd OAI21X1
XOAI21X1_1114 BUFX4_285/Y OAI21X1_1396/C BUFX4_99/Y gnd OAI22X1_53/B vdd OAI21X1
XDFFPOSX1_737 NOR2X1_88/A CLKBUF1_93/Y AOI21X1_47/Y gnd vdd DFFPOSX1
XOAI21X1_1169 NOR2X1_566/Y NOR2X1_567/Y BUFX4_357/Y gnd AOI21X1_489/B vdd OAI21X1
XDFFPOSX1_715 NOR2X1_75/A CLKBUF1_38/Y AOI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_748 INVX1_62/A CLKBUF1_68/Y MUX2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_726 INVX1_55/A CLKBUF1_86/Y MUX2X1_45/Y gnd vdd DFFPOSX1
XOAI21X1_1158 AOI21X1_485/Y AOI21X1_486/Y BUFX4_412/Y gnd NAND2X1_337/B vdd OAI21X1
XINVX1_460 INVX1_460/A gnd INVX1_460/Y vdd INVX1
XDFFPOSX1_759 NOR2X1_92/A CLKBUF1_1/Y AOI21X1_48/Y gnd vdd DFFPOSX1
XAOI21X1_442 INVX1_63/Y BUFX4_365/Y AOI21X1_442/C gnd AOI21X1_443/C vdd AOI21X1
XAOI21X1_431 NOR2X1_175/A BUFX4_90/Y AOI21X1_431/C gnd OAI22X1_43/B vdd AOI21X1
XAOI21X1_420 AOI21X1_420/A AOI21X1_420/B BUFX4_204/Y gnd AOI21X1_421/C vdd AOI21X1
XAOI21X1_453 BUFX4_117/Y AOI21X1_453/B AOI21X1_452/Y gnd AOI21X1_453/Y vdd AOI21X1
XAOI21X1_464 AOI21X1_464/A AOI21X1_464/B BUFX4_411/Y gnd OAI22X1_50/D vdd AOI21X1
XAOI21X1_475 BUFX4_414/Y AOI21X1_475/B AOI21X1_475/C gnd OAI22X1_55/C vdd AOI21X1
XAOI21X1_486 BUFX4_242/Y INVX1_430/Y AOI21X1_486/C gnd AOI21X1_486/Y vdd AOI21X1
XAOI21X1_497 INVX1_84/Y BUFX4_358/Y BUFX4_158/Y gnd AOI21X1_497/Y vdd AOI21X1
XNAND3X1_13 NAND3X1_13/A NAND3X1_13/B NOR3X1_2/Y gnd NOR3X1_3/C vdd NAND3X1
XNAND3X1_46 INVX4_11/A NAND3X1_46/B NOR3X1_7/Y gnd NAND3X1_46/Y vdd NAND3X1
XNAND3X1_35 NAND3X1_35/A NAND3X1_35/B NOR3X1_8/Y gnd NAND3X1_38/B vdd NAND3X1
XNAND3X1_24 AND2X2_7/B AND2X2_7/A NOR3X1_5/Y gnd NOR3X1_6/C vdd NAND3X1
XNAND3X1_57 INVX2_18/Y INVX1_196/Y INVX2_19/Y gnd XOR2X1_2/B vdd NAND3X1
XNAND3X1_68 NAND3X1_68/A NAND3X1_68/B AND2X2_18/A gnd AND2X2_15/B vdd NAND3X1
XNAND3X1_79 BUFX4_38/Y NAND3X1_79/B NAND3X1_79/C gnd AOI22X1_29/A vdd NAND3X1
XNOR2X1_35 NOR2X1_35/A NOR2X1_33/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A AOI21X1_7/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_13 INVX4_1/A INVX1_27/Y gnd INVX2_7/A vdd NOR2X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_47/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_68 NOR2X1_68/A NOR2X1_65/Y gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_57 BUFX4_44/Y BUFX4_385/Y gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_79 NOR2X1_74/B BUFX4_142/Y gnd NOR2X1_83/B vdd NOR2X1
XFILL_43_6_1 gnd vdd FILL
XFILL_42_1_0 gnd vdd FILL
XMUX2X1_20 INVX1_26/Y MUX2X1_8/B MUX2X1_18/S gnd MUX2X1_20/Y vdd MUX2X1
XMUX2X1_42 INVX1_52/Y AND2X2_3/B MUX2X1_42/S gnd MUX2X1_42/Y vdd MUX2X1
XMUX2X1_31 BUFX4_69/Y INVX1_39/Y MUX2X1_31/S gnd MUX2X1_31/Y vdd MUX2X1
XMUX2X1_53 INVX1_63/Y MUX2X1_44/A MUX2X1_51/S gnd MUX2X1_53/Y vdd MUX2X1
XNOR2X1_114 NOR2X1_582/A AOI21X1_62/B gnd NOR2X1_114/Y vdd NOR2X1
XNOR2X1_103 NOR2X1_410/A MUX2X1_75/S gnd NOR2X1_103/Y vdd NOR2X1
XMUX2X1_97 INVX1_110/Y MUX2X1_97/B MUX2X1_97/S gnd MUX2X1_97/Y vdd MUX2X1
XNOR2X1_125 BUFX4_185/Y BUFX4_136/Y gnd AOI21X1_72/B vdd NOR2X1
XMUX2X1_86 INVX1_99/Y MUX2X1_86/B MUX2X1_84/S gnd MUX2X1_86/Y vdd MUX2X1
XNOR2X1_136 NOR2X1_397/A NOR2X1_137/B gnd NOR2X1_136/Y vdd NOR2X1
XNOR2X1_147 NOR2X1_147/A MUX2X1_94/S gnd AOI21X1_87/C vdd NOR2X1
XMUX2X1_75 MUX2X1_77/B INVX1_85/Y MUX2X1_75/S gnd MUX2X1_75/Y vdd MUX2X1
XMUX2X1_64 INVX1_74/Y MUX2X1_64/B MUX2X1_66/S gnd MUX2X1_64/Y vdd MUX2X1
XFILL_34_6_1 gnd vdd FILL
XNOR2X1_158 BUFX4_406/Y NOR2X1_96/B gnd MUX2X1_340/S vdd NOR2X1
XFILL_33_1_0 gnd vdd FILL
XNOR2X1_169 BUFX4_140/Y BUFX4_56/Y gnd NOR2X1_172/B vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XOAI21X1_609 INVX1_264/Y BUFX4_278/Y OAI21X1_609/C gnd MUX2X1_184/B vdd OAI21X1
XMUX2X1_109 MUX2X1_96/A INVX1_122/Y INVX1_219/A gnd MUX2X1_109/Y vdd MUX2X1
XDFFPOSX1_523 NOR2X1_723/A CLKBUF1_52/Y AOI21X1_611/Y gnd vdd DFFPOSX1
XDFFPOSX1_512 INVX1_320/A CLKBUF1_17/Y MUX2X1_382/Y gnd vdd DFFPOSX1
XDFFPOSX1_501 NOR2X1_483/B CLKBUF1_68/Y AOI21X1_605/Y gnd vdd DFFPOSX1
XDFFPOSX1_545 INVX1_387/A CLKBUF1_97/Y DFFPOSX1_545/D gnd vdd DFFPOSX1
XDFFPOSX1_556 AND2X2_30/B CLKBUF1_23/Y OAI21X1_1540/Y gnd vdd DFFPOSX1
XDFFPOSX1_534 INVX1_440/A CLKBUF1_64/Y MUX2X1_391/Y gnd vdd DFFPOSX1
XDFFPOSX1_578 INVX1_461/A CLKBUF1_35/Y MUX2X1_407/Y gnd vdd DFFPOSX1
XDFFPOSX1_567 OAI21X1_613/B CLKBUF1_5/Y DFFPOSX1_567/D gnd vdd DFFPOSX1
XDFFPOSX1_589 NOR2X1_486/A CLKBUF1_25/Y DFFPOSX1_589/D gnd vdd DFFPOSX1
XINVX1_290 INVX1_290/A gnd INVX1_290/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XNAND2X1_90 NAND2X1_90/A NAND2X1_6/B gnd NAND2X1_90/Y vdd NAND2X1
XFILL_0_6_1 gnd vdd FILL
XFILL_25_6_1 gnd vdd FILL
XNOR2X1_670 NOR2X1_670/A MUX2X1_88/S gnd NOR2X1_670/Y vdd NOR2X1
XFILL_24_1_0 gnd vdd FILL
XNOR2X1_681 NOR2X1_545/A MUX2X1_94/S gnd NOR2X1_681/Y vdd NOR2X1
XNOR2X1_692 NOR2X1_692/A NOR2X1_167/B gnd NOR2X1_692/Y vdd NOR2X1
XAOI21X1_261 AND2X2_52/A NOR2X1_698/A AOI21X1_261/C gnd OAI22X1_4/D vdd AOI21X1
XAOI21X1_250 BUFX4_349/Y INVX1_223/Y AOI21X1_250/C gnd AOI21X1_250/Y vdd AOI21X1
XAOI21X1_294 NAND2X1_94/A BUFX4_413/Y BUFX4_333/Y gnd AOI21X1_294/Y vdd AOI21X1
XAOI21X1_272 BUFX4_416/Y MUX2X1_179/Y BUFX4_205/Y gnd AOI22X1_13/A vdd AOI21X1
XAOI21X1_283 BUFX4_49/Y AOI22X1_15/Y BUFX4_401/Y gnd AOI22X1_17/B vdd AOI21X1
XFILL_8_7_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XDFFPOSX1_1052 INVX1_340/A CLKBUF1_52/Y OAI21X1_331/Y gnd vdd DFFPOSX1
XDFFPOSX1_1030 INVX1_144/A CLKBUF1_34/Y MUX2X1_131/Y gnd vdd DFFPOSX1
XDFFPOSX1_1041 NOR2X1_243/A CLKBUF1_42/Y AOI21X1_154/Y gnd vdd DFFPOSX1
XOAI21X1_439 traffic_Street_1[1] traffic_Street_1[2] traffic_Street_1[3] gnd NAND3X1_5/A
+ vdd OAI21X1
XOAI21X1_417 BUFX4_58/Y BUFX4_464/Y AOI21X1_449/A gnd OAI21X1_417/Y vdd OAI21X1
XOAI21X1_406 OAI21X1_40/A MUX2X1_71/B OAI21X1_406/C gnd OAI21X1_406/Y vdd OAI21X1
XOAI21X1_428 OAI21X1_54/A BUFX4_470/Y OAI21X1_427/Y gnd OAI21X1_428/Y vdd OAI21X1
XDFFPOSX1_331 AND2X2_27/B CLKBUF1_6/Y AOI21X1_547/Y gnd vdd DFFPOSX1
XDFFPOSX1_320 OAI21X1_947/B CLKBUF1_16/Y DFFPOSX1_320/D gnd vdd DFFPOSX1
XDFFPOSX1_364 INVX1_366/A CLKBUF1_61/Y MUX2X1_303/Y gnd vdd DFFPOSX1
XDFFPOSX1_353 INVX1_418/A CLKBUF1_55/Y MUX2X1_312/Y gnd vdd DFFPOSX1
XDFFPOSX1_342 INVX1_232/A CLKBUF1_51/Y MUX2X1_315/Y gnd vdd DFFPOSX1
XDFFPOSX1_397 INVX1_304/A CLKBUF1_24/Y MUX2X1_267/Y gnd vdd DFFPOSX1
XDFFPOSX1_375 NOR2X1_414/B CLKBUF1_58/Y DFFPOSX1_375/D gnd vdd DFFPOSX1
XDFFPOSX1_386 INVX1_221/A CLKBUF1_8/Y MUX2X1_279/Y gnd vdd DFFPOSX1
XFILL_40_4_1 gnd vdd FILL
XOAI21X1_940 BUFX4_33/Y INVX1_368/Y BUFX4_340/Y gnd OAI21X1_941/A vdd OAI21X1
XOAI21X1_951 BUFX4_278/Y INVX1_374/Y OAI21X1_951/C gnd OAI21X1_951/Y vdd OAI21X1
XOAI21X1_984 NOR2X1_490/Y OAI21X1_984/B OAI21X1_982/Y gnd NOR2X1_491/B vdd OAI21X1
XOAI21X1_973 BUFX4_231/Y INVX1_460/A OAI21X1_973/C gnd OAI21X1_975/C vdd OAI21X1
XOAI21X1_962 OAI21X1_962/A OAI21X1_962/B BUFX4_410/Y gnd AOI21X1_420/B vdd OAI21X1
XOAI21X1_995 INVX1_114/Y BUFX4_89/Y BUFX4_246/Y gnd AOI21X1_431/C vdd OAI21X1
XFILL_48_5_1 gnd vdd FILL
XFILL_47_0_0 gnd vdd FILL
XOAI21X1_11 OAI21X1_11/A MUX2X1_9/B OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_33 BUFX4_125/Y BUFX4_293/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_22 OAI21X1_24/A MUX2X1_6/B OAI21X1_22/C gnd OAI21X1_22/Y vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XOAI21X1_44 BUFX4_443/Y OAI21X1_48/B OAI21X1_43/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_77 BUFX4_448/Y BUFX4_43/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_66 BUFX4_316/Y OAI21X1_64/B OAI21X1_65/Y gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_55 INVX4_4/A BUFX4_462/Y INVX1_392/A gnd OAI21X1_56/C vdd OAI21X1
XOAI21X1_88 NAND2X1_32/Y BUFX4_372/Y OAI21X1_87/Y gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_99 BUFX4_120/Y BUFX4_479/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XFILL_39_5_1 gnd vdd FILL
XFILL_38_0_0 gnd vdd FILL
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_203 BUFX4_174/Y NAND2X1_60/Y OAI21X1_203/C gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_247 BUFX4_466/Y NAND2X1_68/Y OAI21X1_246/Y gnd OAI21X1_247/Y vdd OAI21X1
XOAI21X1_236 BUFX4_123/Y BUFX4_139/Y AND2X2_43/A gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_225 NAND2X1_64/Y BUFX4_216/Y OAI21X1_224/Y gnd OAI21X1_225/Y vdd OAI21X1
XOAI21X1_214 BUFX4_452/Y BUFX4_408/Y NOR2X1_588/A gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_258 BUFX4_126/Y BUFX4_433/Y OAI21X1_900/A gnd OAI21X1_259/C vdd OAI21X1
XOAI21X1_269 NAND2X1_72/Y BUFX4_380/Y OAI21X1_269/C gnd OAI21X1_269/Y vdd OAI21X1
XAND2X2_14 AND2X2_14/A AND2X2_14/B gnd AND2X2_14/Y vdd AND2X2
XAND2X2_25 AND2X2_25/A AND2X2_25/B gnd AND2X2_25/Y vdd AND2X2
XAND2X2_47 AND2X2_47/A AND2X2_47/B gnd AND2X2_47/Y vdd AND2X2
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XDFFPOSX1_161 INVX1_419/A CLKBUF1_41/Y MUX2X1_348/Y gnd vdd DFFPOSX1
XDFFPOSX1_150 NOR2X1_694/A CLKBUF1_27/Y AOI21X1_582/Y gnd vdd DFFPOSX1
XDFFPOSX1_172 NOR2X1_644/A CLKBUF1_34/Y AOI21X1_532/Y gnd vdd DFFPOSX1
XDFFPOSX1_183 NAND2X1_228/B CLKBUF1_15/Y DFFPOSX1_183/D gnd vdd DFFPOSX1
XDFFPOSX1_194 OAI21X1_581/B CLKBUF1_45/Y OAI21X1_1391/Y gnd vdd DFFPOSX1
XNAND2X1_220 NOR2X1_178/A BUFX4_220/Y gnd NAND2X1_220/Y vdd NAND2X1
XNAND2X1_242 BUFX4_225/Y NAND2X1_242/B gnd OAI21X1_783/C vdd NAND2X1
XNAND2X1_253 NOR2X1_112/A BUFX4_263/Y gnd NAND2X1_253/Y vdd NAND2X1
XNAND2X1_231 BUFX4_411/Y NAND2X1_231/B gnd AOI22X1_20/B vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_286 AND2X2_36/B NAND2X1_286/B gnd OAI21X1_963/C vdd NAND2X1
XNAND2X1_264 INVX1_168/A BUFX4_291/Y gnd NAND2X1_264/Y vdd NAND2X1
XNAND2X1_275 BUFX4_251/Y NOR2X1_653/A gnd OAI21X1_914/C vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_297 OAI21X1_63/C BUFX4_242/Y gnd OAI21X1_989/C vdd NAND2X1
XFILL_29_0_0 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XOAI21X1_770 NOR2X1_426/Y OAI21X1_769/Y OAI21X1_770/C gnd OAI21X1_770/Y vdd OAI21X1
XOAI21X1_792 BUFX4_48/Y OAI21X1_792/B AOI21X1_346/Y gnd OAI21X1_819/C vdd OAI21X1
XOAI21X1_781 OAI21X1_780/Y BUFX4_37/Y INVX8_29/A gnd OAI21X1_781/Y vdd OAI21X1
XMUX2X1_270 BUFX4_65/Y INVX1_362/Y NOR2X1_57/Y gnd MUX2X1_270/Y vdd MUX2X1
XMUX2X1_281 BUFX4_66/Y INVX1_348/Y MUX2X1_45/S gnd MUX2X1_281/Y vdd MUX2X1
XMUX2X1_292 INVX1_364/Y BUFX4_68/Y MUX2X1_51/S gnd MUX2X1_292/Y vdd MUX2X1
XCLKBUF1_12 BUFX4_8/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_23 BUFX4_5/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_45 BUFX4_8/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_56 BUFX4_6/Y gnd CLKBUF1_56/Y vdd CLKBUF1
XCLKBUF1_34 BUFX4_6/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XCLKBUF1_78 BUFX4_2/Y gnd CLKBUF1_78/Y vdd CLKBUF1
XCLKBUF1_67 BUFX4_4/Y gnd CLKBUF1_67/Y vdd CLKBUF1
XCLKBUF1_89 BUFX4_4/Y gnd CLKBUF1_89/Y vdd CLKBUF1
XINVX1_108 INVX1_108/A gnd MUX2X1_95/B vdd INVX1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XBUFX4_428 INVX8_3/Y gnd BUFX4_428/Y vdd BUFX4
XBUFX4_417 address[2] gnd BUFX4_417/Y vdd BUFX4
XBUFX4_406 INVX8_21/Y gnd BUFX4_406/Y vdd BUFX4
XBUFX4_439 INVX8_2/Y gnd BUFX4_439/Y vdd BUFX4
XFILL_45_3_1 gnd vdd FILL
XOAI21X1_1329 BUFX4_58/Y BUFX4_396/Y AOI21X1_470/B gnd OAI21X1_1329/Y vdd OAI21X1
XOAI21X1_1307 BUFX4_443/Y NAND2X1_39/Y OAI21X1_1307/C gnd DFFPOSX1_182/D vdd OAI21X1
XOAI21X1_1318 BUFX4_449/Y BUFX4_53/Y INVX1_365/A gnd OAI21X1_1318/Y vdd OAI21X1
XDFFPOSX1_919 NOR2X1_399/A CLKBUF1_27/Y AOI21X1_106/Y gnd vdd DFFPOSX1
XDFFPOSX1_908 INVX1_111/A CLKBUF1_83/Y MUX2X1_98/Y gnd vdd DFFPOSX1
XFILL_36_3_1 gnd vdd FILL
XAOI21X1_624 BUFX4_441/Y NOR2X1_737/B NOR2X1_736/Y gnd AOI21X1_624/Y vdd AOI21X1
XAOI21X1_613 BUFX4_67/Y NOR2X1_234/Y NOR2X1_725/Y gnd AOI21X1_613/Y vdd AOI21X1
XAOI21X1_602 BUFX4_422/Y NOR2X1_220/B NOR2X1_714/Y gnd AOI21X1_602/Y vdd AOI21X1
XFILL_2_3_1 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XBUFX4_203 address[3] gnd AND2X2_48/B vdd BUFX4
XBUFX4_214 INVX8_11/Y gnd BUFX4_214/Y vdd BUFX4
XBUFX4_236 BUFX4_20/Y gnd BUFX4_236/Y vdd BUFX4
XBUFX4_225 BUFX4_20/Y gnd BUFX4_225/Y vdd BUFX4
XBUFX4_269 BUFX4_21/Y gnd AND2X2_25/B vdd BUFX4
XFILL_18_3_1 gnd vdd FILL
XBUFX4_247 BUFX4_23/Y gnd BUFX4_247/Y vdd BUFX4
XBUFX4_258 BUFX4_20/Y gnd BUFX4_258/Y vdd BUFX4
XNOR2X1_307 NOR2X1_304/Y AND2X2_4/Y gnd AOI22X1_10/D vdd NOR2X1
XNOR2X1_329 INVX2_24/A INVX1_209/A gnd INVX1_205/A vdd NOR2X1
XNOR2X1_318 NOR2X1_311/B NAND3X1_36/Y gnd NOR2X1_318/Y vdd NOR2X1
XOAI21X1_1104 INVX1_417/Y BUFX4_275/Y BUFX4_158/Y gnd AOI21X1_470/C vdd OAI21X1
XOAI21X1_1137 NAND2X1_8/A AND2X2_37/B BUFX4_109/Y gnd OAI22X1_61/B vdd OAI21X1
XDFFPOSX1_705 NOR2X1_68/A CLKBUF1_19/Y AOI21X1_34/Y gnd vdd DFFPOSX1
XOAI21X1_1126 BUFX4_104/Y AOI21X1_476/Y OAI21X1_1125/Y gnd OAI21X1_1126/Y vdd OAI21X1
XOAI21X1_1115 BUFX4_367/Y NOR2X1_689/A BUFX4_148/Y gnd OAI22X1_54/C vdd OAI21X1
XDFFPOSX1_738 INVX1_60/A CLKBUF1_23/Y MUX2X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_716 INVX1_47/A CLKBUF1_38/Y OAI21X1_91/Y gnd vdd DFFPOSX1
XOAI21X1_1148 INVX1_40/Y BUFX4_237/Y NAND2X1_336/Y gnd MUX2X1_257/A vdd OAI21X1
XDFFPOSX1_727 NOR2X1_80/A CLKBUF1_68/Y AOI21X1_41/Y gnd vdd DFFPOSX1
XOAI21X1_1159 BUFX4_244/Y INVX1_431/Y AOI21X1_487/Y gnd OAI21X1_1159/Y vdd OAI21X1
XINVX1_461 INVX1_461/A gnd INVX1_461/Y vdd INVX1
XDFFPOSX1_749 INVX1_63/A CLKBUF1_54/Y MUX2X1_53/Y gnd vdd DFFPOSX1
XINVX1_450 INVX1_450/A gnd INVX1_450/Y vdd INVX1
XAOI21X1_410 BUFX4_345/Y AOI21X1_410/B AOI21X1_410/C gnd NOR2X1_480/B vdd AOI21X1
XAOI21X1_443 BUFX4_108/Y AOI21X1_443/B AOI21X1_443/C gnd AOI21X1_443/Y vdd AOI21X1
XAOI21X1_421 BUFX4_205/Y MUX2X1_235/Y AOI21X1_421/C gnd NAND2X1_285/B vdd AOI21X1
XAOI21X1_432 NOR2X1_182/A BUFX4_94/Y AOI21X1_432/C gnd OAI22X1_43/C vdd AOI21X1
XAOI21X1_454 INVX8_32/A AOI21X1_454/B NOR2X1_512/Y gnd AOI21X1_454/Y vdd AOI21X1
XAOI21X1_465 BUFX4_263/Y INVX1_412/Y BUFX4_86/Y gnd AOI21X1_465/Y vdd AOI21X1
XAOI21X1_476 BUFX4_354/Y AOI21X1_476/B NOR2X1_547/Y gnd AOI21X1_476/Y vdd AOI21X1
XAOI21X1_487 AND2X2_47/B AOI21X1_487/B BUFX4_116/Y gnd AOI21X1_487/Y vdd AOI21X1
XAOI21X1_498 AND2X2_41/A INVX1_121/Y BUFX4_89/Y gnd AOI21X1_498/Y vdd AOI21X1
XNAND3X1_14 INVX2_15/A NAND3X1_14/B OR2X2_4/Y gnd AOI22X1_3/D vdd NAND3X1
XNAND3X1_47 INVX1_202/Y XNOR2X1_4/B NOR3X1_7/Y gnd NAND3X1_47/Y vdd NAND3X1
XNAND3X1_36 INVX1_194/Y NAND3X1_36/B INVX1_195/Y gnd NAND3X1_36/Y vdd NAND3X1
XNAND3X1_25 INVX4_7/A NAND3X1_17/B NAND3X1_17/C gnd NAND3X1_25/Y vdd NAND3X1
XNAND3X1_58 NAND3X1_58/A NAND3X1_58/B NAND3X1_58/C gnd NAND3X1_59/B vdd NAND3X1
XNAND3X1_69 INVX1_218/Y INVX1_217/A AND2X2_16/Y gnd NAND3X1_69/Y vdd NAND3X1
XNOR2X1_25 NOR2X1_25/A AOI21X1_7/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_36 NOR2X1_36/A NOR2X1_33/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_14 INVX2_7/Y INVX2_6/Y gnd INVX8_5/A vdd NOR2X1
XNOR2X1_58 NOR2X1_58/A NOR2X1_57/Y gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_65/Y gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XFILL_42_1_1 gnd vdd FILL
XMUX2X1_10 INVX1_15/Y MUX2X1_18/B MUX2X1_9/S gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_21 INVX1_28/Y MUX2X1_9/B MUX2X1_21/S gnd MUX2X1_21/Y vdd MUX2X1
XNOR2X1_115 INVX2_3/A INVX1_3/Y gnd INVX2_11/A vdd NOR2X1
XMUX2X1_32 BUFX4_316/Y INVX1_40/Y MUX2X1_31/S gnd MUX2X1_32/Y vdd MUX2X1
XMUX2X1_43 MUX2X1_64/B INVX1_53/Y MUX2X1_45/S gnd MUX2X1_43/Y vdd MUX2X1
XNOR2X1_104 NOR2X1_104/A MUX2X1_75/S gnd AOI21X1_57/C vdd NOR2X1
XMUX2X1_54 INVX1_64/Y MUX2X1_58/A MUX2X1_51/S gnd MUX2X1_54/Y vdd MUX2X1
XNOR2X1_137 NOR2X1_137/A NOR2X1_137/B gnd AOI21X1_80/C vdd NOR2X1
XMUX2X1_87 INVX1_100/Y MUX2X1_83/B MUX2X1_84/S gnd MUX2X1_87/Y vdd MUX2X1
XNOR2X1_148 NOR2X1_599/A MUX2X1_94/S gnd AOI21X1_88/C vdd NOR2X1
XNOR2X1_126 NOR2X1_394/A AOI21X1_72/B gnd NOR2X1_126/Y vdd NOR2X1
XMUX2X1_65 INVX1_75/Y BUFX4_371/Y MUX2X1_66/S gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_76 INVX1_86/Y MUX2X1_71/B MUX2X1_76/S gnd MUX2X1_76/Y vdd MUX2X1
XFILL_33_1_1 gnd vdd FILL
XNOR2X1_159 NOR2X1_159/A MUX2X1_340/S gnd AOI21X1_95/C vdd NOR2X1
XMUX2X1_98 INVX1_111/Y MUX2X1_96/A MUX2X1_97/S gnd MUX2X1_98/Y vdd MUX2X1
XDFFPOSX1_513 INVX1_383/A CLKBUF1_48/Y MUX2X1_383/Y gnd vdd DFFPOSX1
XDFFPOSX1_502 NOR2X1_565/B CLKBUF1_18/Y AOI21X1_606/Y gnd vdd DFFPOSX1
XDFFPOSX1_524 NOR2X1_724/A CLKBUF1_56/Y AOI21X1_612/Y gnd vdd DFFPOSX1
XDFFPOSX1_546 INVX1_438/A CLKBUF1_92/Y DFFPOSX1_546/D gnd vdd DFFPOSX1
XDFFPOSX1_535 MUX2X1_182/A CLKBUF1_36/Y DFFPOSX1_535/D gnd vdd DFFPOSX1
XDFFPOSX1_557 NAND2X1_292/B CLKBUF1_97/Y DFFPOSX1_557/D gnd vdd DFFPOSX1
XDFFPOSX1_579 INVX1_271/A CLKBUF1_53/Y MUX2X1_408/Y gnd vdd DFFPOSX1
XDFFPOSX1_568 OAI21X1_793/B CLKBUF1_14/Y DFFPOSX1_568/D gnd vdd DFFPOSX1
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XNAND2X1_91 NAND2X1_91/A NAND2X1_6/B gnd NAND2X1_91/Y vdd NAND2X1
XNAND2X1_80 INVX8_26/A INVX4_4/Y gnd NAND2X1_80/Y vdd NAND2X1
XNOR2X1_671 NOR2X1_671/A NOR2X1_137/B gnd NOR2X1_671/Y vdd NOR2X1
XNOR2X1_660 NOR2X1_660/A AOI21X1_62/B gnd NOR2X1_660/Y vdd NOR2X1
XFILL_24_1_1 gnd vdd FILL
XNOR2X1_693 NOR2X1_693/A NOR2X1_172/B gnd NOR2X1_693/Y vdd NOR2X1
XNOR2X1_682 NOR2X1_421/B MUX2X1_96/S gnd NOR2X1_682/Y vdd NOR2X1
XAOI21X1_240 INVX1_210/A NAND3X1_65/C INVX4_9/A gnd AOI22X1_8/A vdd AOI21X1
XAOI21X1_251 BUFX4_226/Y INVX1_224/Y OAI21X1_557/Y gnd AOI21X1_251/Y vdd AOI21X1
XAOI21X1_284 BUFX4_154/Y INVX1_268/Y OAI21X1_613/Y gnd AOI21X1_284/Y vdd AOI21X1
XAOI21X1_273 BUFX4_262/Y AOI21X1_273/B BUFX4_94/Y gnd AOI21X1_273/Y vdd AOI21X1
XAOI21X1_262 BUFX4_148/Y INVX1_240/Y OAI21X1_579/Y gnd OAI21X1_580/A vdd AOI21X1
XAOI21X1_295 NAND2X1_90/A BUFX4_36/Y AOI21X1_295/C gnd NOR2X1_377/B vdd AOI21X1
XOAI21X1_1490 NAND2X1_75/Y BUFX4_445/Y OAI21X1_1489/Y gnd OAI21X1_1490/Y vdd OAI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_44_9_0 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XDFFPOSX1_1020 INVX1_138/A CLKBUF1_56/Y MUX2X1_125/Y gnd vdd DFFPOSX1
XDFFPOSX1_1053 INVX1_406/A CLKBUF1_97/Y OAI21X1_333/Y gnd vdd DFFPOSX1
XDFFPOSX1_1031 NOR2X1_235/A CLKBUF1_57/Y AOI21X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_1042 AND2X2_55/A CLKBUF1_42/Y AOI21X1_155/Y gnd vdd DFFPOSX1
XFILL_35_9_0 gnd vdd FILL
XOAI21X1_429 BUFX4_191/Y BUFX4_461/Y OAI21X1_429/C gnd OAI21X1_429/Y vdd OAI21X1
XOAI21X1_418 MUX2X1_61/B OAI21X1_48/B OAI21X1_417/Y gnd OAI21X1_418/Y vdd OAI21X1
XOAI21X1_407 NOR2X1_39/A INVX4_2/A AOI21X1_382/A gnd OAI21X1_407/Y vdd OAI21X1
XDFFPOSX1_310 INVX1_249/A CLKBUF1_42/Y MUX2X1_319/Y gnd vdd DFFPOSX1
XDFFPOSX1_321 OAI21X1_1119/B CLKBUF1_75/Y DFFPOSX1_321/D gnd vdd DFFPOSX1
XDFFPOSX1_365 INVX1_451/A CLKBUF1_95/Y MUX2X1_304/Y gnd vdd DFFPOSX1
XDFFPOSX1_354 NAND2X1_175/B CLKBUF1_99/Y OAI21X1_1324/Y gnd vdd DFFPOSX1
XDFFPOSX1_332 NOR2X1_660/A CLKBUF1_99/Y AOI21X1_548/Y gnd vdd DFFPOSX1
XDFFPOSX1_343 INVX1_297/A CLKBUF1_6/Y MUX2X1_316/Y gnd vdd DFFPOSX1
XDFFPOSX1_398 NOR2X1_626/A CLKBUF1_70/Y AOI21X1_514/Y gnd vdd DFFPOSX1
XDFFPOSX1_387 INVX1_302/A CLKBUF1_13/Y MUX2X1_280/Y gnd vdd DFFPOSX1
XDFFPOSX1_376 INVX1_365/A CLKBUF1_22/Y OAI21X1_1319/Y gnd vdd DFFPOSX1
XFILL_1_9_0 gnd vdd FILL
XFILL_26_9_0 gnd vdd FILL
XNOR2X1_490 NOR2X1_19/A BUFX4_85/Y gnd NOR2X1_490/Y vdd NOR2X1
XOAI21X1_941 OAI21X1_941/A NOR2X1_478/Y BUFX4_108/Y gnd OAI22X1_39/D vdd OAI21X1
XOAI21X1_952 INVX1_375/Y BUFX4_280/Y BUFX4_113/Y gnd OAI21X1_953/A vdd OAI21X1
XOAI21X1_930 INVX1_359/Y BUFX4_100/Y BUFX4_328/Y gnd OAI21X1_931/A vdd OAI21X1
XOAI21X1_963 INVX1_383/Y BUFX4_287/Y OAI21X1_963/C gnd MUX2X1_236/B vdd OAI21X1
XOAI21X1_985 BUFX4_360/Y NOR2X1_30/A BUFX4_149/Y gnd OAI22X1_40/C vdd OAI21X1
XOAI21X1_974 BUFX4_232/Y OAI21X1_974/B BUFX4_80/Y gnd OAI21X1_974/Y vdd OAI21X1
XOAI21X1_996 MUX2X1_99/A BUFX4_92/Y BUFX4_328/Y gnd OAI21X1_997/A vdd OAI21X1
XFILL_47_0_1 gnd vdd FILL
XFILL_17_9_0 gnd vdd FILL
XOAI21X1_45 BUFX4_62/Y BUFX4_460/Y OAI21X1_45/C gnd OAI21X1_46/C vdd OAI21X1
XOAI21X1_34 NAND2X1_24/Y MUX2X1_8/B OAI21X1_33/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_12 BUFX4_295/Y BUFX4_299/Y OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_23 BUFX4_450/Y BUFX4_292/Y NOR2X1_492/A gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_67 BUFX4_301/Y BUFX4_45/Y NOR2X1_400/A gnd OAI21X1_68/C vdd OAI21X1
XOAI21X1_78 NAND2X1_31/Y BUFX4_173/Y OAI21X1_77/Y gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_56 OAI21X1_54/A BUFX4_69/Y OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_89 BUFX4_124/Y BUFX4_45/Y OAI21X1_89/C gnd OAI21X1_90/C vdd OAI21X1
XFILL_38_0_1 gnd vdd FILL
XFILL_50_7_0 gnd vdd FILL
XOAI21X1_204 BUFX4_142/Y BUFX4_405/Y MUX2X1_245/B gnd OAI21X1_204/Y vdd OAI21X1
XOAI21X1_237 NAND2X1_66/Y BUFX4_377/Y OAI21X1_236/Y gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_215 NAND2X1_61/Y BUFX4_465/Y OAI21X1_214/Y gnd OAI21X1_215/Y vdd OAI21X1
XOAI21X1_226 BUFX4_383/Y BUFX4_138/Y AND2X2_32/A gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_259 NAND2X1_70/Y BUFX4_177/Y OAI21X1_259/C gnd OAI21X1_259/Y vdd OAI21X1
XOAI21X1_248 BUFX4_384/Y BUFX4_434/Y OAI21X1_248/C gnd OAI21X1_248/Y vdd OAI21X1
XAND2X2_15 AND2X2_15/A AND2X2_15/B gnd AND2X2_15/Y vdd AND2X2
XAND2X2_37 AND2X2_37/A AND2X2_37/B gnd AND2X2_37/Y vdd AND2X2
XAND2X2_26 AND2X2_26/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XDFFPOSX1_140 INVX1_398/A CLKBUF1_94/Y OAI21X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 INVX1_222/A CLKBUF1_43/Y MUX2X1_269/Y gnd vdd DFFPOSX1
XDFFPOSX1_173 INVX1_414/A CLKBUF1_85/Y MUX2X1_289/Y gnd vdd DFFPOSX1
XDFFPOSX1_151 INVX1_308/A CLKBUF1_22/Y MUX2X1_349/Y gnd vdd DFFPOSX1
XAND2X2_48 AND2X2_48/A AND2X2_48/B gnd AND2X2_48/Y vdd AND2X2
XNAND2X1_210 NAND2X1_210/A BUFX4_369/Y gnd OAI21X1_666/C vdd NAND2X1
XDFFPOSX1_184 AOI21X1_407/B CLKBUF1_83/Y DFFPOSX1_184/D gnd vdd DFFPOSX1
XDFFPOSX1_195 INVX1_311/A CLKBUF1_8/Y OAI21X1_1393/Y gnd vdd DFFPOSX1
XNAND2X1_243 BUFX4_227/Y NOR2X1_724/A gnd NAND2X1_243/Y vdd NAND2X1
XNAND2X1_221 NOR2X1_181/A BUFX4_222/Y gnd NAND2X1_221/Y vdd NAND2X1
XNAND2X1_232 AND2X2_25/B NOR2X1_693/A gnd OAI21X1_751/C vdd NAND2X1
XNAND2X1_254 NOR2X1_155/A AND2X2_29/A gnd OAI21X1_843/C vdd NAND2X1
XNAND2X1_287 BUFX4_288/Y NOR2X1_725/A gnd NAND2X1_287/Y vdd NAND2X1
XNAND2X1_265 NAND2X1_95/A BUFX4_220/Y gnd NAND2X1_265/Y vdd NAND2X1
XNAND2X1_276 NAND2X1_276/A AOI21X1_393/Y gnd AOI22X1_24/A vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XNAND2X1_298 BUFX4_37/Y OAI22X1_41/Y gnd OAI21X1_992/C vdd NAND2X1
XFILL_41_7_0 gnd vdd FILL
XOAI21X1_760 AND2X2_41/A OAI21X1_760/B BUFX4_117/Y gnd OAI22X1_20/B vdd OAI21X1
XOAI21X1_793 BUFX4_153/Y OAI21X1_793/B BUFX4_350/Y gnd OAI21X1_793/Y vdd OAI21X1
XOAI21X1_771 OAI21X1_770/Y BUFX4_50/Y BUFX4_400/Y gnd OAI21X1_771/Y vdd OAI21X1
XOAI21X1_782 NOR2X1_430/Y OAI21X1_781/Y OAI21X1_782/C gnd OAI21X1_792/B vdd OAI21X1
XMUX2X1_271 BUFX4_65/Y INVX1_361/Y NOR2X1_60/Y gnd MUX2X1_271/Y vdd MUX2X1
XMUX2X1_260 MUX2X1_260/A MUX2X1_260/B BUFX4_32/Y gnd MUX2X1_260/Y vdd MUX2X1
XMUX2X1_282 BUFX4_324/Y INVX1_410/Y MUX2X1_45/S gnd MUX2X1_282/Y vdd MUX2X1
XMUX2X1_293 INVX1_448/Y BUFX4_324/Y MUX2X1_51/S gnd MUX2X1_293/Y vdd MUX2X1
XFILL_49_8_0 gnd vdd FILL
XFILL_32_7_0 gnd vdd FILL
XCLKBUF1_24 BUFX4_7/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_13 BUFX4_9/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_35 BUFX4_1/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_57 BUFX4_6/Y gnd CLKBUF1_57/Y vdd CLKBUF1
XCLKBUF1_46 BUFX4_10/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XCLKBUF1_79 BUFX4_5/Y gnd CLKBUF1_79/Y vdd CLKBUF1
XCLKBUF1_68 BUFX4_2/Y gnd CLKBUF1_68/Y vdd CLKBUF1
XFILL_23_7_0 gnd vdd FILL
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XFILL_6_8_0 gnd vdd FILL
XBUFX4_418 address[2] gnd BUFX4_418/Y vdd BUFX4
XBUFX4_429 INVX8_3/Y gnd BUFX4_429/Y vdd BUFX4
XBUFX4_407 INVX8_21/Y gnd BUFX4_407/Y vdd BUFX4
XFILL_14_7_0 gnd vdd FILL
XOAI21X1_1319 NAND2X1_40/Y BUFX4_66/Y OAI21X1_1318/Y gnd OAI21X1_1319/Y vdd OAI21X1
XOAI21X1_1308 BUFX4_61/Y BUFX4_54/Y NAND2X1_228/B gnd OAI21X1_1308/Y vdd OAI21X1
XOAI21X1_590 BUFX4_256/Y OAI21X1_590/B BUFX4_92/Y gnd AOI21X1_270/C vdd OAI21X1
XDFFPOSX1_909 INVX1_112/A CLKBUF1_13/Y MUX2X1_99/Y gnd vdd DFFPOSX1
XFILL_39_1 gnd vdd FILL
XAOI21X1_614 BUFX4_322/Y NOR2X1_234/Y NOR2X1_726/Y gnd AOI21X1_614/Y vdd AOI21X1
XAOI21X1_625 MUX2X1_18/B NOR2X1_737/B NOR2X1_737/Y gnd AOI21X1_625/Y vdd AOI21X1
XAOI21X1_603 BUFX4_445/Y NOR2X1_716/B NOR2X1_715/Y gnd AOI21X1_603/Y vdd AOI21X1
XBUFX4_215 INVX8_11/Y gnd MUX2X1_59/B vdd BUFX4
XBUFX4_226 BUFX4_23/Y gnd BUFX4_226/Y vdd BUFX4
XBUFX4_237 BUFX4_19/Y gnd BUFX4_237/Y vdd BUFX4
XBUFX4_204 address[3] gnd BUFX4_204/Y vdd BUFX4
XFILL_46_6_0 gnd vdd FILL
XBUFX4_248 BUFX4_21/Y gnd BUFX4_248/Y vdd BUFX4
XBUFX4_259 BUFX4_22/Y gnd BUFX4_259/Y vdd BUFX4
XNOR2X1_319 INVX4_7/A BUFX4_307/Y gnd NOR2X1_319/Y vdd NOR2X1
XNOR2X1_308 AND2X2_6/B NOR2X1_308/B gnd NOR3X1_4/B vdd NOR2X1
XOAI21X1_1138 BUFX4_334/Y INVX1_21/A BUFX4_157/Y gnd OAI22X1_62/C vdd OAI21X1
XOAI21X1_1127 OAI21X1_1126/Y BUFX4_417/Y INVX8_29/A gnd OAI22X1_59/C vdd OAI21X1
XOAI21X1_1105 INVX1_418/Y BUFX4_277/Y BUFX4_96/Y gnd AOI21X1_471/C vdd OAI21X1
XOAI21X1_1116 BUFX4_287/Y OAI21X1_1116/B BUFX4_100/Y gnd OAI22X1_54/B vdd OAI21X1
XOAI21X1_1149 NOR2X1_43/A BUFX4_368/Y AOI21X1_482/Y gnd OAI21X1_1150/C vdd OAI21X1
XDFFPOSX1_706 NOR2X1_69/A CLKBUF1_80/Y AOI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_739 INVX1_289/A CLKBUF1_92/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_728 NOR2X1_81/A CLKBUF1_38/Y AOI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_717 NOR2X1_76/A CLKBUF1_54/Y AOI21X1_39/Y gnd vdd DFFPOSX1
XINVX1_451 INVX1_451/A gnd INVX1_451/Y vdd INVX1
XINVX1_440 INVX1_440/A gnd INVX1_440/Y vdd INVX1
XFILL_37_6_0 gnd vdd FILL
XAOI21X1_400 BUFX4_92/Y OAI21X1_925/Y AOI21X1_399/Y gnd OAI22X1_37/C vdd AOI21X1
XAOI21X1_433 NOR2X1_138/A BUFX4_249/Y AOI21X1_433/C gnd OAI22X1_44/B vdd AOI21X1
XFILL_20_5_0 gnd vdd FILL
XAOI21X1_411 BUFX4_272/Y INVX1_371/Y AOI21X1_411/C gnd AOI21X1_411/Y vdd AOI21X1
XAOI21X1_422 OAI21X1_965/Y AOI21X1_422/B BUFX4_411/Y gnd AOI21X1_423/C vdd AOI21X1
XAOI21X1_477 BUFX4_354/Y INVX1_423/Y BUFX4_150/Y gnd AOI21X1_477/Y vdd AOI21X1
XAOI21X1_466 BUFX4_90/Y AOI21X1_466/B AOI21X1_466/C gnd AOI21X1_466/Y vdd AOI21X1
XAOI21X1_444 INVX1_75/Y BUFX4_280/Y AOI21X1_444/C gnd AOI21X1_444/Y vdd AOI21X1
XAOI21X1_455 AOI21X1_455/A BUFX4_241/Y BUFX4_77/Y gnd AOI21X1_455/Y vdd AOI21X1
XAOI21X1_499 NOR2X1_172/A BUFX4_287/Y AOI21X1_499/C gnd AOI21X1_499/Y vdd AOI21X1
XAOI21X1_488 NOR2X1_710/A BUFX4_328/Y BUFX4_118/Y gnd AOI21X1_488/Y vdd AOI21X1
XNAND3X1_48 INVX2_24/A NAND3X1_58/A NAND3X1_58/C gnd NAND3X1_48/Y vdd NAND3X1
XNAND3X1_15 AND2X2_5/B INVX2_15/A NAND3X1_15/C gnd NAND3X1_17/B vdd NAND3X1
XNAND3X1_26 NOR3X1_5/Y NAND3X1_26/B AND2X2_7/Y gnd NAND3X1_26/Y vdd NAND3X1
XNAND3X1_37 NAND3X1_37/A NAND3X1_26/B NOR2X1_318/Y gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_59 INVX4_9/Y NAND3X1_59/B NAND3X1_59/C gnd NAND3X1_59/Y vdd NAND3X1
XFILL_3_6_0 gnd vdd FILL
XNOR2X1_26 INVX1_14/Y XNOR2X1_8/A gnd INVX8_8/A vdd NOR2X1
XNOR2X1_15 INVX1_1/Y XNOR2X1_8/A gnd INVX8_6/A vdd NOR2X1
XNOR2X1_37 INVX4_1/Y INVX1_27/Y gnd INVX2_8/A vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNOR2X1_59 NOR2X1_59/A NOR2X1_57/Y gnd NOR2X1_59/Y vdd NOR2X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_47/B gnd NOR2X1_48/Y vdd NOR2X1
XFILL_11_5_0 gnd vdd FILL
XMUX2X1_11 INVX1_16/Y BUFX4_71/Y MUX2X1_9/S gnd MUX2X1_11/Y vdd MUX2X1
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_33 BUFX4_173/Y INVX1_41/Y NOR2X1_54/Y gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_22 INVX1_29/Y BUFX4_421/Y MUX2X1_21/S gnd MUX2X1_22/Y vdd MUX2X1
XNOR2X1_105 NOR2X1_105/A MUX2X1_75/S gnd AOI21X1_58/C vdd NOR2X1
XMUX2X1_44 MUX2X1_44/A INVX1_54/Y MUX2X1_45/S gnd MUX2X1_44/Y vdd MUX2X1
XMUX2X1_66 INVX1_76/Y MUX2X1_66/B MUX2X1_66/S gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_88 MUX2X1_40/B MUX2X1_88/B MUX2X1_88/S gnd MUX2X1_88/Y vdd MUX2X1
XNOR2X1_138 NOR2X1_138/A NOR2X1_137/B gnd NOR2X1_138/Y vdd NOR2X1
XNOR2X1_127 NOR2X1_127/A AOI21X1_72/B gnd NOR2X1_127/Y vdd NOR2X1
XNOR2X1_116 INVX2_10/Y INVX2_11/Y gnd INVX8_19/A vdd NOR2X1
XNOR2X1_149 INVX2_7/Y INVX2_11/Y gnd INVX8_21/A vdd NOR2X1
XMUX2X1_77 INVX1_87/Y MUX2X1_77/B MUX2X1_76/S gnd MUX2X1_77/Y vdd MUX2X1
XMUX2X1_55 MUX2X1_59/B INVX1_65/Y MUX2X1_55/S gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_99 MUX2X1_99/A BUFX4_377/Y MUX2X1_97/S gnd MUX2X1_99/Y vdd MUX2X1
XDFFPOSX1_514 INVX1_436/A CLKBUF1_2/Y MUX2X1_384/Y gnd vdd DFFPOSX1
XDFFPOSX1_503 INVX1_265/A CLKBUF1_79/Y OAI21X1_1498/Y gnd vdd DFFPOSX1
XDFFPOSX1_547 NOR2X1_730/A CLKBUF1_56/Y AOI21X1_618/Y gnd vdd DFFPOSX1
XDFFPOSX1_525 NOR2X1_725/A CLKBUF1_32/Y AOI21X1_613/Y gnd vdd DFFPOSX1
XDFFPOSX1_536 OAI21X1_791/B CLKBUF1_60/Y OAI21X1_1524/Y gnd vdd DFFPOSX1
XINVX1_270 INVX1_270/A gnd INVX1_270/Y vdd INVX1
XDFFPOSX1_569 INVX1_390/A CLKBUF1_14/Y OAI21X1_1550/Y gnd vdd DFFPOSX1
XDFFPOSX1_558 AND2X2_53/B CLKBUF1_92/Y DFFPOSX1_558/D gnd vdd DFFPOSX1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XINVX1_292 INVX1_292/A gnd INVX1_292/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_70 INVX8_23/A INVX4_5/Y gnd NAND2X1_70/Y vdd NAND2X1
XNAND2X1_92 NAND2X1_92/A NAND2X1_6/B gnd NAND2X1_92/Y vdd NAND2X1
XNAND2X1_81 INVX8_26/A INVX8_9/A gnd NAND2X1_81/Y vdd NAND2X1
XNOR2X1_650 NOR2X1_650/A NOR2X1_97/B gnd NOR2X1_650/Y vdd NOR2X1
XNOR2X1_661 NOR2X1_525/A AOI21X1_62/B gnd NOR2X1_661/Y vdd NOR2X1
XNOR2X1_694 NOR2X1_694/A MUX2X1_102/S gnd NOR2X1_694/Y vdd NOR2X1
XNOR2X1_672 NOR2X1_425/A NOR2X1_137/B gnd NOR2X1_672/Y vdd NOR2X1
XNOR2X1_683 NOR2X1_683/A MUX2X1_96/S gnd NOR2X1_683/Y vdd NOR2X1
XAOI21X1_230 INVX2_20/A NOR3X1_7/Y INVX2_25/A gnd AOI21X1_230/Y vdd AOI21X1
XAOI21X1_241 AOI21X1_225/Y NAND3X1_64/Y AOI21X1_241/C gnd NOR3X1_13/C vdd AOI21X1
XAOI21X1_252 NOR2X1_642/A BUFX4_150/Y BUFX4_227/Y gnd AOI21X1_252/Y vdd AOI21X1
XAOI21X1_274 NOR2X1_707/A BUFX4_341/Y BUFX4_96/Y gnd OAI21X1_596/C vdd AOI21X1
XAOI21X1_263 BUFX4_148/Y INVX1_241/Y AOI21X1_263/C gnd OAI21X1_583/A vdd AOI21X1
XAOI21X1_285 BUFX4_154/Y INVX1_269/Y OAI21X1_614/Y gnd AOI21X1_285/Y vdd AOI21X1
XAOI21X1_296 INVX1_155/A BUFX4_31/Y AOI21X1_296/C gnd OAI21X1_639/B vdd AOI21X1
XOAI21X1_1491 BUFX4_456/Y BUFX4_298/Y NOR2X1_435/B gnd OAI21X1_1492/C vdd OAI21X1
XOAI21X1_1480 BUFX4_318/Y NAND2X1_73/Y OAI21X1_1479/Y gnd OAI21X1_1480/Y vdd OAI21X1
XFILL_44_9_1 gnd vdd FILL
XFILL_43_4_0 gnd vdd FILL
XDFFPOSX1_1010 NOR2X1_226/A CLKBUF1_18/Y AOI21X1_143/Y gnd vdd DFFPOSX1
XDFFPOSX1_1054 INVX1_444/A CLKBUF1_52/Y OAI21X1_335/Y gnd vdd DFFPOSX1
XDFFPOSX1_1032 NOR2X1_236/A CLKBUF1_56/Y AOI21X1_149/Y gnd vdd DFFPOSX1
XDFFPOSX1_1021 INVX1_139/A CLKBUF1_79/Y MUX2X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_1043 OAI21X1_320/C CLKBUF1_36/Y OAI21X1_321/Y gnd vdd DFFPOSX1
XFILL_35_9_1 gnd vdd FILL
XFILL_34_4_0 gnd vdd FILL
XFILL_21_1 gnd vdd FILL
XOAI21X1_408 OAI21X1_40/A MUX2X1_77/B OAI21X1_407/Y gnd OAI21X1_408/Y vdd OAI21X1
XOAI21X1_419 BUFX4_62/Y NOR2X1_39/A OAI21X1_419/C gnd OAI21X1_419/Y vdd OAI21X1
XDFFPOSX1_300 INVX1_373/A CLKBUF1_23/Y MUX2X1_323/Y gnd vdd DFFPOSX1
XDFFPOSX1_311 NOR2X1_423/A CLKBUF1_85/Y AOI21X1_552/Y gnd vdd DFFPOSX1
XDFFPOSX1_322 NAND2X1_177/B CLKBUF1_17/Y OAI21X1_1343/Y gnd vdd DFFPOSX1
XDFFPOSX1_355 AOI21X1_319/B CLKBUF1_6/Y DFFPOSX1_355/D gnd vdd DFFPOSX1
XDFFPOSX1_344 INVX1_342/A CLKBUF1_51/Y MUX2X1_317/Y gnd vdd DFFPOSX1
XDFFPOSX1_333 NOR2X1_525/A CLKBUF1_77/Y AOI21X1_549/Y gnd vdd DFFPOSX1
XDFFPOSX1_366 INVX1_449/A CLKBUF1_37/Y MUX2X1_297/Y gnd vdd DFFPOSX1
XDFFPOSX1_388 INVX1_348/A CLKBUF1_38/Y MUX2X1_281/Y gnd vdd DFFPOSX1
XDFFPOSX1_377 NOR2X1_530/B CLKBUF1_10/Y OAI21X1_1321/Y gnd vdd DFFPOSX1
XDFFPOSX1_399 INVX1_412/A CLKBUF1_94/Y MUX2X1_268/Y gnd vdd DFFPOSX1
XFILL_26_9_1 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XFILL_1_9_1 gnd vdd FILL
XFILL_25_4_0 gnd vdd FILL
XNOR2X1_480 BUFX4_394/Y NOR2X1_480/B gnd NOR2X1_480/Y vdd NOR2X1
XNOR2X1_491 BUFX4_415/Y NOR2X1_491/B gnd NOR2X1_491/Y vdd NOR2X1
XOAI21X1_920 OAI21X1_920/A AND2X2_38/Y OAI21X1_918/Y gnd OAI21X1_920/Y vdd OAI21X1
XOAI21X1_942 MUX2X1_231/Y BUFX4_366/Y BUFX4_109/Y gnd OAI21X1_942/Y vdd OAI21X1
XOAI21X1_931 OAI21X1_931/A AND2X2_40/Y BUFX4_412/Y gnd OAI22X1_38/D vdd OAI21X1
XOAI21X1_964 INVX1_384/Y BUFX4_289/Y NAND2X1_287/Y gnd MUX2X1_236/A vdd OAI21X1
XOAI21X1_975 NOR2X1_486/Y OAI21X1_974/Y OAI21X1_975/C gnd NOR2X1_487/B vdd OAI21X1
XOAI21X1_953 OAI21X1_953/A AND2X2_41/Y OAI21X1_951/Y gnd MUX2X1_235/B vdd OAI21X1
XOAI21X1_986 OAI21X1_31/C AND2X2_22/A BUFX4_86/Y gnd OAI22X1_40/B vdd OAI21X1
XOAI21X1_997 OAI21X1_997/A AND2X2_42/Y BUFX4_35/Y gnd OAI22X1_43/A vdd OAI21X1
XFILL_8_5_0 gnd vdd FILL
XFILL_16_4_0 gnd vdd FILL
XFILL_17_9_1 gnd vdd FILL
XOAI21X1_13 OAI21X1_11/A BUFX4_421/Y OAI21X1_12/Y gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_24 OAI21X1_24/A BUFX4_64/Y OAI21X1_23/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_35 BUFX4_464/Y BUFX4_303/Y OAI21X1_35/C gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_68 NAND2X1_30/Y BUFX4_214/Y OAI21X1_68/C gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_57 INVX4_4/A BUFX4_464/Y INVX1_426/A gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_46 MUX2X1_27/B OAI21X1_48/B OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_79 BUFX4_448/Y BUFX4_42/Y NOR2X1_499/A gnd OAI21X1_79/Y vdd OAI21X1
XFILL_50_7_1 gnd vdd FILL
XOAI21X1_216 BUFX4_119/Y BUFX4_408/Y INVX1_286/A gnd OAI21X1_217/C vdd OAI21X1
XOAI21X1_205 MUX2X1_57/A NAND2X1_60/Y OAI21X1_204/Y gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_238 BUFX4_123/Y BUFX4_138/Y OAI21X1_238/C gnd OAI21X1_239/C vdd OAI21X1
XOAI21X1_227 NAND2X1_64/Y MUX2X1_96/A OAI21X1_226/Y gnd OAI21X1_227/Y vdd OAI21X1
XOAI21X1_249 NAND2X1_69/Y MUX2X1_97/B OAI21X1_248/Y gnd OAI21X1_249/Y vdd OAI21X1
XAND2X2_38 BUFX4_256/Y AND2X2_38/B gnd AND2X2_38/Y vdd AND2X2
XDFFPOSX1_130 INVX1_184/A CLKBUF1_96/Y MUX2X1_170/Y gnd vdd DFFPOSX1
XAND2X2_27 AND2X2_27/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XAND2X2_16 AND2X2_16/A INVX1_215/Y gnd AND2X2_16/Y vdd AND2X2
XAND2X2_49 AND2X2_49/A BUFX4_256/Y gnd AND2X2_49/Y vdd AND2X2
XDFFPOSX1_141 OAI21X1_73/C CLKBUF1_70/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_163 NOR2X1_627/A CLKBUF1_43/Y AOI21X1_515/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 NOR2X1_695/A CLKBUF1_65/Y AOI21X1_583/Y gnd vdd DFFPOSX1
XNAND2X1_211 BUFX4_35/Y OAI22X1_11/Y gnd OAI21X1_669/C vdd NAND2X1
XNAND2X1_200 NOR2X1_266/A AND2X2_51/B gnd OAI21X1_643/C vdd NAND2X1
XDFFPOSX1_185 DFFPOSX1_185/Q CLKBUF1_58/Y OAI21X1_1313/Y gnd vdd DFFPOSX1
XDFFPOSX1_174 NOR2X1_370/B CLKBUF1_45/Y DFFPOSX1_174/D gnd vdd DFFPOSX1
XDFFPOSX1_196 MUX2X1_230/B CLKBUF1_8/Y DFFPOSX1_196/D gnd vdd DFFPOSX1
XNAND2X1_222 NOR2X1_87/A BUFX4_230/Y gnd NAND2X1_222/Y vdd NAND2X1
XNAND2X1_244 NAND2X1_244/A BUFX4_336/Y gnd NAND2X1_244/Y vdd NAND2X1
XNAND2X1_233 BUFX4_273/Y NOR2X1_687/A gnd NAND2X1_233/Y vdd NAND2X1
XNAND2X1_266 NOR2X1_252/A BUFX4_224/Y gnd NAND2X1_266/Y vdd NAND2X1
XNAND2X1_277 BUFX4_38/Y NAND2X1_277/B gnd AOI21X1_397/B vdd NAND2X1
XNAND2X1_255 BUFX4_416/Y OAI22X1_26/Y gnd NAND2X1_255/Y vdd NAND2X1
XNAND2X1_299 INVX8_29/A NAND2X1_299/B gnd OAI21X1_993/C vdd NAND2X1
XNAND2X1_288 BUFX4_291/Y NOR2X1_727/A gnd NAND2X1_288/Y vdd NAND2X1
XFILL_41_7_1 gnd vdd FILL
XFILL_40_2_0 gnd vdd FILL
XOAI21X1_750 OAI21X1_750/A AND2X2_29/Y OAI21X1_748/Y gnd NAND2X1_231/B vdd OAI21X1
XOAI21X1_772 INVX1_315/Y BUFX4_288/Y NAND2X1_237/Y gnd MUX2X1_211/B vdd OAI21X1
XOAI21X1_761 INVX1_312/Y BUFX4_281/Y NAND2X1_235/Y gnd MUX2X1_210/B vdd OAI21X1
XOAI21X1_794 BUFX4_146/Y NOR2X1_737/A BUFX4_236/Y gnd AOI21X1_348/C vdd OAI21X1
XOAI21X1_783 INVX1_320/Y BUFX4_226/Y OAI21X1_783/C gnd MUX2X1_214/B vdd OAI21X1
XMUX2X1_250 MUX2X1_250/A MUX2X1_250/B BUFX4_118/Y gnd MUX2X1_250/Y vdd MUX2X1
XMUX2X1_272 MUX2X1_1/B INVX1_224/Y NOR2X1_70/Y gnd MUX2X1_272/Y vdd MUX2X1
XMUX2X1_283 BUFX4_63/Y INVX1_347/Y NOR2X1_83/B gnd MUX2X1_283/Y vdd MUX2X1
XMUX2X1_261 MUX2X1_261/A MUX2X1_261/B BUFX4_86/Y gnd MUX2X1_261/Y vdd MUX2X1
XMUX2X1_294 BUFX4_443/Y INVX1_228/Y MUX2X1_55/S gnd MUX2X1_294/Y vdd MUX2X1
XFILL_49_8_1 gnd vdd FILL
XFILL_48_3_0 gnd vdd FILL
XFILL_32_7_1 gnd vdd FILL
XFILL_31_2_0 gnd vdd FILL
XCLKBUF1_14 BUFX4_2/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XCLKBUF1_25 BUFX4_1/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_47 BUFX4_2/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XCLKBUF1_36 BUFX4_5/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XCLKBUF1_69 BUFX4_1/Y gnd CLKBUF1_69/Y vdd CLKBUF1
XCLKBUF1_58 BUFX4_3/Y gnd CLKBUF1_58/Y vdd CLKBUF1
XFILL_39_3_0 gnd vdd FILL
XBUFX4_90 BUFX4_75/A gnd BUFX4_90/Y vdd BUFX4
XFILL_23_7_1 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XFILL_6_8_1 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XBUFX4_419 address[2] gnd BUFX4_419/Y vdd BUFX4
XBUFX4_408 INVX8_21/Y gnd BUFX4_408/Y vdd BUFX4
XFILL_14_7_1 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_1309 BUFX4_420/Y NAND2X1_39/Y OAI21X1_1308/Y gnd DFFPOSX1_183/D vdd OAI21X1
XOAI21X1_591 INVX1_250/Y BUFX4_259/Y OAI21X1_591/C gnd MUX2X1_179/B vdd OAI21X1
XOAI21X1_580 OAI21X1_580/A NOR2X1_371/Y BUFX4_415/Y gnd AOI21X1_265/A vdd OAI21X1
XAOI21X1_626 BUFX4_65/Y NOR2X1_737/B NOR2X1_738/Y gnd AOI21X1_626/Y vdd AOI21X1
XAOI21X1_615 BUFX4_73/Y NOR2X1_727/B NOR2X1_727/Y gnd AOI21X1_615/Y vdd AOI21X1
XAOI21X1_604 BUFX4_429/Y NOR2X1_716/B NOR2X1_716/Y gnd AOI21X1_604/Y vdd AOI21X1
XBUFX4_227 BUFX4_23/Y gnd BUFX4_227/Y vdd BUFX4
XBUFX4_205 address[3] gnd BUFX4_205/Y vdd BUFX4
XBUFX4_216 INVX8_11/Y gnd BUFX4_216/Y vdd BUFX4
XFILL_46_6_1 gnd vdd FILL
XBUFX4_249 BUFX4_24/Y gnd BUFX4_249/Y vdd BUFX4
XBUFX4_238 BUFX4_17/Y gnd AND2X2_51/B vdd BUFX4
XFILL_45_1_0 gnd vdd FILL
XNOR2X1_309 OR2X2_5/B OR2X2_5/A gnd NOR2X1_309/Y vdd NOR2X1
XOAI21X1_1128 OAI22X1_59/Y INVX8_28/A BUFX4_400/Y gnd OAI22X1_60/C vdd OAI21X1
XOAI21X1_1106 AOI21X1_470/Y AOI21X1_471/Y BUFX4_37/Y gnd NAND2X1_333/B vdd OAI21X1
XOAI21X1_1117 OAI22X1_54/Y BUFX4_40/Y BUFX4_168/Y gnd OAI22X1_55/B vdd OAI21X1
XDFFPOSX1_718 INVX1_48/A CLKBUF1_41/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XOAI21X1_1139 INVX1_26/A BUFX4_230/Y BUFX4_110/Y gnd OAI22X1_62/B vdd OAI21X1
XDFFPOSX1_707 OAI21X1_83/C CLKBUF1_28/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_729 NOR2X1_82/A CLKBUF1_12/Y AOI21X1_43/Y gnd vdd DFFPOSX1
XINVX1_452 INVX1_452/A gnd INVX1_452/Y vdd INVX1
XINVX1_441 INVX1_441/A gnd INVX1_441/Y vdd INVX1
XINVX1_430 INVX1_430/A gnd INVX1_430/Y vdd INVX1
XFILL_51_1 gnd vdd FILL
XFILL_37_6_1 gnd vdd FILL
XFILL_36_1_0 gnd vdd FILL
XAOI21X1_401 BUFX4_94/Y NOR2X1_695/A OAI21X1_926/Y gnd OAI22X1_38/B vdd AOI21X1
XFILL_20_5_1 gnd vdd FILL
XAOI21X1_412 BUFX4_153/Y AOI21X1_412/B AOI21X1_411/Y gnd MUX2X1_234/B vdd AOI21X1
XAOI21X1_423 BUFX4_412/Y MUX2X1_236/Y AOI21X1_423/C gnd AOI22X1_26/C vdd AOI21X1
XAOI21X1_434 BUFX4_366/Y AOI21X1_434/B AOI21X1_434/C gnd AOI21X1_434/Y vdd AOI21X1
XAOI21X1_467 BUFX4_92/Y AOI21X1_467/B AOI21X1_467/C gnd AOI21X1_467/Y vdd AOI21X1
XAOI21X1_445 BUFX4_417/Y MUX2X1_249/Y BUFX4_171/Y gnd AOI22X1_30/B vdd AOI21X1
XAOI21X1_456 NOR2X1_208/A BUFX4_246/Y AOI21X1_456/C gnd AOI21X1_456/Y vdd AOI21X1
XAOI21X1_478 INVX8_31/A INVX1_424/Y AND2X2_32/B gnd AOI21X1_478/Y vdd AOI21X1
XAOI21X1_489 AOI21X1_489/A AOI21X1_489/B BUFX4_413/Y gnd AOI21X1_489/Y vdd AOI21X1
XNAND3X1_27 INVX4_6/A INVX1_187/Y NAND3X1_7/C gnd NAND3X1_27/Y vdd NAND3X1
XNAND3X1_16 INVX4_6/Y INVX1_190/Y NAND3X1_16/C gnd NAND3X1_16/Y vdd NAND3X1
XNAND3X1_38 NOR2X1_309/Y NAND3X1_38/B NAND3X1_37/Y gnd BUFX4_306/A vdd NAND3X1
XNAND3X1_49 INVX1_200/A INVX1_203/A NOR3X1_7/Y gnd AOI22X1_6/C vdd NAND3X1
XNOR2X1_27 BUFX4_294/Y BUFX4_133/Y gnd NOR2X1_30/B vdd NOR2X1
XNOR2X1_16 NOR2X1_16/A BUFX4_57/Y gnd NOR2X1_16/Y vdd NOR2X1
XFILL_28_6_1 gnd vdd FILL
XFILL_3_6_1 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_38 INVX2_6/Y INVX2_8/Y gnd INVX8_10/A vdd NOR2X1
XNOR2X1_49 BUFX4_461/Y BUFX4_121/Y gnd MUX2X1_31/S vdd NOR2X1
XFILL_27_1_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XMUX2X1_34 MUX2X1_82/B INVX1_42/Y NOR2X1_54/Y gnd MUX2X1_34/Y vdd MUX2X1
XMUX2X1_12 INVX1_17/Y MUX2X1_8/B MUX2X1_9/S gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_23 INVX1_30/Y BUFX4_71/Y MUX2X1_21/S gnd MUX2X1_23/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_106 BUFX4_396/Y NOR2X1_96/B gnd NOR2X1_107/B vdd NOR2X1
XMUX2X1_45 BUFX4_465/Y INVX1_55/Y MUX2X1_45/S gnd MUX2X1_45/Y vdd MUX2X1
XNOR2X1_139 NOR2X1_596/A NOR2X1_137/B gnd AOI21X1_82/C vdd NOR2X1
XNOR2X1_128 NOR2X1_128/A AOI21X1_72/B gnd AOI21X1_74/C vdd NOR2X1
XNOR2X1_117 BUFX4_297/Y BUFX4_186/Y gnd NAND2X1_50/B vdd NOR2X1
XMUX2X1_78 INVX1_88/Y MUX2X1_61/B MUX2X1_76/S gnd MUX2X1_78/Y vdd MUX2X1
XMUX2X1_56 MUX2X1_64/B INVX1_66/Y MUX2X1_55/S gnd MUX2X1_56/Y vdd MUX2X1
XMUX2X1_67 INVX1_77/Y MUX2X1_71/B MUX2X1_70/S gnd MUX2X1_67/Y vdd MUX2X1
XMUX2X1_89 BUFX4_214/Y MUX2X1_89/B MUX2X1_89/S gnd MUX2X1_89/Y vdd MUX2X1
XDFFPOSX1_504 NOR2X1_434/A CLKBUF1_79/Y DFFPOSX1_504/D gnd vdd DFFPOSX1
XDFFPOSX1_515 NAND2X1_187/B CLKBUF1_62/Y DFFPOSX1_515/D gnd vdd DFFPOSX1
XDFFPOSX1_526 NOR2X1_726/A CLKBUF1_32/Y AOI21X1_614/Y gnd vdd DFFPOSX1
XDFFPOSX1_537 INVX1_386/A CLKBUF1_18/Y OAI21X1_1526/Y gnd vdd DFFPOSX1
XDFFPOSX1_559 INVX1_268/A CLKBUF1_53/Y MUX2X1_398/Y gnd vdd DFFPOSX1
XDFFPOSX1_548 NOR2X1_731/A CLKBUF1_57/Y AOI21X1_619/Y gnd vdd DFFPOSX1
XINVX1_271 INVX1_271/A gnd INVX1_271/Y vdd INVX1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 INVX8_21/A INVX8_7/A gnd NAND2X1_60/Y vdd NAND2X1
XNAND2X1_93 NAND2X1_93/A NAND2X1_6/B gnd NAND2X1_93/Y vdd NAND2X1
XNAND2X1_82 INVX8_27/A INVX4_3/Y gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_71 INVX8_23/A INVX8_9/A gnd MUX2X1_366/S vdd NAND2X1
XNOR2X1_640 NOR2X1_640/A NOR2X1_83/B gnd NOR2X1_640/Y vdd NOR2X1
XNOR2X1_662 NOR2X1_422/B NAND2X1_50/B gnd NOR2X1_662/Y vdd NOR2X1
XNOR2X1_651 NOR2X1_412/B NOR2X1_97/B gnd NOR2X1_651/Y vdd NOR2X1
XNOR2X1_673 NOR2X1_673/A NOR2X1_137/B gnd NOR2X1_673/Y vdd NOR2X1
XNOR2X1_695 NOR2X1_695/A MUX2X1_102/S gnd NOR2X1_695/Y vdd NOR2X1
XNOR2X1_684 NOR2X1_684/A NOR2X1_155/B gnd NOR2X1_684/Y vdd NOR2X1
XAOI21X1_231 NAND3X1_56/C AOI21X1_231/B OAI21X1_504/Y gnd OAI21X1_506/A vdd AOI21X1
XAOI21X1_242 INVX4_10/Y AOI21X1_242/B OAI21X1_497/A gnd AOI21X1_242/Y vdd AOI21X1
XAOI21X1_220 NAND3X1_30/Y OAI21X1_471/Y NAND3X1_31/Y gnd AOI21X1_221/B vdd AOI21X1
XAOI21X1_275 BUFX4_369/Y INVX1_257/Y AOI21X1_275/C gnd OAI21X1_601/A vdd AOI21X1
XAOI21X1_253 BUFX4_412/Y OAI21X1_562/Y BUFX4_167/Y gnd AOI22X1_11/B vdd AOI21X1
XAOI21X1_264 BUFX4_148/Y INVX1_242/Y AOI21X1_264/C gnd OAI21X1_583/B vdd AOI21X1
XAOI21X1_286 BUFX4_154/Y INVX1_270/Y AOI21X1_286/C gnd AOI21X1_286/Y vdd AOI21X1
XAOI21X1_297 OAI21X1_634/Y NOR2X1_377/Y AOI21X1_297/C gnd OAI22X1_8/A vdd AOI21X1
XOAI21X1_1492 NAND2X1_75/Y BUFX4_429/Y OAI21X1_1492/C gnd DFFPOSX1_496/D vdd OAI21X1
XOAI21X1_1481 BUFX4_192/Y BUFX4_160/Y AND2X2_23/B gnd OAI21X1_1481/Y vdd OAI21X1
XOAI21X1_1470 NAND2X1_72/Y BUFX4_72/Y OAI21X1_1470/C gnd OAI21X1_1470/Y vdd OAI21X1
XFILL_43_4_1 gnd vdd FILL
XDFFPOSX1_1011 OAI21X1_661/A CLKBUF1_36/Y OAI21X1_297/Y gnd vdd DFFPOSX1
XDFFPOSX1_1000 NOR2X1_470/A CLKBUF1_74/Y OAI21X1_283/Y gnd vdd DFFPOSX1
XDFFPOSX1_1022 INVX1_140/A CLKBUF1_62/Y MUX2X1_127/Y gnd vdd DFFPOSX1
XDFFPOSX1_1033 NOR2X1_237/A CLKBUF1_56/Y AOI21X1_150/Y gnd vdd DFFPOSX1
XDFFPOSX1_1044 OAI21X1_889/A CLKBUF1_36/Y OAI21X1_323/Y gnd vdd DFFPOSX1
XDFFPOSX1_1055 NOR2X1_251/A CLKBUF1_52/Y AOI21X1_160/Y gnd vdd DFFPOSX1
XFILL_34_4_1 gnd vdd FILL
XFILL_21_2 gnd vdd FILL
XOAI21X1_409 BUFX4_464/Y INVX4_2/A INVX1_402/A gnd OAI21X1_410/C vdd OAI21X1
XDFFPOSX1_301 INVX1_454/A CLKBUF1_48/Y MUX2X1_324/Y gnd vdd DFFPOSX1
XDFFPOSX1_312 INVX1_371/A CLKBUF1_16/Y MUX2X1_320/Y gnd vdd DFFPOSX1
XDFFPOSX1_323 OAI21X1_759/B CLKBUF1_75/Y DFFPOSX1_323/D gnd vdd DFFPOSX1
XDFFPOSX1_356 NAND2X1_274/B CLKBUF1_6/Y DFFPOSX1_356/D gnd vdd DFFPOSX1
XDFFPOSX1_334 INVX1_233/A CLKBUF1_55/Y OAI21X1_1333/Y gnd vdd DFFPOSX1
XDFFPOSX1_345 INVX1_453/A CLKBUF1_58/Y MUX2X1_318/Y gnd vdd DFFPOSX1
XDFFPOSX1_378 NOR2X1_640/A CLKBUF1_86/Y AOI21X1_528/Y gnd vdd DFFPOSX1
XDFFPOSX1_367 INVX1_450/A CLKBUF1_55/Y MUX2X1_298/Y gnd vdd DFFPOSX1
XDFFPOSX1_389 INVX1_410/A CLKBUF1_13/Y MUX2X1_282/Y gnd vdd DFFPOSX1
XFILL_0_4_1 gnd vdd FILL
XFILL_25_4_1 gnd vdd FILL
XNOR2X1_470 NOR2X1_470/A BUFX4_331/Y gnd OAI22X1_35/A vdd NOR2X1
XNOR2X1_481 BUFX4_362/Y INVX1_377/Y gnd NOR2X1_481/Y vdd NOR2X1
XNOR2X1_492 NOR2X1_492/A AND2X2_51/B gnd OAI22X1_40/D vdd NOR2X1
XOAI21X1_910 AOI21X1_392/Y NOR2X1_624/A OAI21X1_910/C gnd OAI21X1_910/Y vdd OAI21X1
XOAI21X1_921 INVX1_351/Y BUFX4_258/Y BUFX4_91/Y gnd AOI21X1_398/C vdd OAI21X1
XOAI21X1_932 BUFX4_102/Y NOR2X1_634/A OAI21X1_932/C gnd NAND2X1_280/A vdd OAI21X1
XOAI21X1_943 INVX1_369/Y BUFX4_418/Y NAND2X1_281/Y gnd AOI21X1_410/B vdd OAI21X1
XOAI21X1_954 BUFX4_370/Y INVX1_376/Y OAI21X1_954/C gnd OAI21X1_956/C vdd OAI21X1
XOAI21X1_976 INVX1_25/Y BUFX4_233/Y BUFX4_81/Y gnd AOI21X1_427/C vdd OAI21X1
XOAI21X1_965 NOR2X1_482/Y NOR2X1_483/Y BUFX4_290/Y gnd OAI21X1_965/Y vdd OAI21X1
XOAI21X1_987 OAI22X1_40/Y BUFX4_36/Y BUFX4_169/Y gnd OAI21X1_987/Y vdd OAI21X1
XOAI21X1_998 INVX1_120/Y BUFX4_93/Y BUFX4_247/Y gnd AOI21X1_432/C vdd OAI21X1
XMUX2X1_410 BUFX4_71/Y INVX1_391/Y MUX2X1_410/S gnd MUX2X1_410/Y vdd MUX2X1
XFILL_8_5_1 gnd vdd FILL
XDFFPOSX1_890 NOR2X1_586/A CLKBUF1_33/Y OAI21X1_207/Y gnd vdd DFFPOSX1
XFILL_7_0_0 gnd vdd FILL
XFILL_16_4_1 gnd vdd FILL
XOAI21X1_14 NOR2X1_16/A BUFX4_299/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_25 BUFX4_450/Y BUFX4_293/Y NOR2X1_560/A gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_47 BUFX4_62/Y BUFX4_460/Y OAI21X1_47/C gnd OAI21X1_48/C vdd OAI21X1
XOAI21X1_69 BUFX4_301/Y BUFX4_44/Y INVX1_332/A gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_58 OAI21X1_54/A BUFX4_316/Y OAI21X1_57/Y gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_36 OAI21X1_40/A BUFX4_443/Y OAI21X1_35/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_217 NAND2X1_62/Y AND2X2_2/B OAI21X1_217/C gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_206 BUFX4_143/Y BUFX4_404/Y NOR2X1_586/A gnd OAI21X1_207/C vdd OAI21X1
XOAI21X1_228 BUFX4_383/Y BUFX4_139/Y AND2X2_42/A gnd OAI21X1_228/Y vdd OAI21X1
XOAI21X1_239 NAND2X1_66/Y BUFX4_465/Y OAI21X1_239/C gnd OAI21X1_239/Y vdd OAI21X1
XAND2X2_17 AND2X2_17/A INVX4_9/Y gnd AND2X2_17/Y vdd AND2X2
XAND2X2_28 BUFX4_258/Y AND2X2_28/B gnd AND2X2_28/Y vdd AND2X2
XDFFPOSX1_120 NOR2X1_292/A CLKBUF1_63/Y AOI21X1_195/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 NOR2X1_696/A CLKBUF1_86/Y AOI21X1_584/Y gnd vdd DFFPOSX1
XDFFPOSX1_142 OAI21X1_557/B CLKBUF1_28/Y DFFPOSX1_142/D gnd vdd DFFPOSX1
XDFFPOSX1_164 INVX1_362/A CLKBUF1_35/Y MUX2X1_270/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 INVX1_185/A CLKBUF1_6/Y MUX2X1_171/Y gnd vdd DFFPOSX1
XAND2X2_39 BUFX4_95/Y AND2X2_39/B gnd AND2X2_39/Y vdd AND2X2
XNAND2X1_201 NOR2X1_282/A BUFX4_240/Y gnd NAND2X1_201/Y vdd NAND2X1
XDFFPOSX1_175 INVX1_309/A CLKBUF1_33/Y OAI21X1_1409/Y gnd vdd DFFPOSX1
XDFFPOSX1_197 OAI21X1_1396/C CLKBUF1_33/Y DFFPOSX1_197/D gnd vdd DFFPOSX1
XDFFPOSX1_186 OAI21X1_582/B CLKBUF1_8/Y OAI21X1_1399/Y gnd vdd DFFPOSX1
XNAND2X1_223 OAI21X1_101/C BUFX4_232/Y gnd OAI21X1_705/C vdd NAND2X1
XNAND2X1_212 INVX8_30/A OAI21X1_672/Y gnd AND2X2_26/B vdd NAND2X1
XNAND2X1_234 BUFX4_40/Y OAI21X1_757/Y gnd OAI21X1_758/C vdd NAND2X1
XNAND2X1_267 DFFPOSX1_7/Q BUFX4_226/Y gnd OAI21X1_887/C vdd NAND2X1
XNAND2X1_278 BUFX4_261/Y NOR2X1_680/A gnd NAND2X1_278/Y vdd NAND2X1
XNAND2X1_245 OAI21X1_795/Y OAI21X1_798/Y gnd NAND2X1_245/Y vdd NAND2X1
XNAND2X1_256 BUFX4_40/Y NAND2X1_256/B gnd AOI22X1_22/C vdd NAND2X1
XNAND2X1_289 BUFX4_220/Y NOR2X1_729/A gnd OAI21X1_968/C vdd NAND2X1
XFILL_40_2_1 gnd vdd FILL
XOAI21X1_740 BUFX4_110/Y NOR2X1_633/A AOI21X1_326/Y gnd AOI21X1_328/A vdd OAI21X1
XOAI21X1_751 INVX1_307/Y BUFX4_270/Y OAI21X1_751/C gnd AOI21X1_331/B vdd OAI21X1
XOAI21X1_773 BUFX4_348/Y INVX1_316/Y NAND2X1_238/Y gnd MUX2X1_211/A vdd OAI21X1
XOAI21X1_762 INVX1_313/Y BUFX4_283/Y OAI21X1_762/C gnd MUX2X1_210/A vdd OAI21X1
XOAI21X1_784 INVX1_321/Y AND2X2_37/B NAND2X1_243/Y gnd MUX2X1_214/A vdd OAI21X1
XOAI21X1_795 OAI21X1_795/A OAI21X1_795/B BUFX4_34/Y gnd OAI21X1_795/Y vdd OAI21X1
XMUX2X1_240 MUX2X1_240/A MUX2X1_240/B BUFX4_87/Y gnd MUX2X1_240/Y vdd MUX2X1
XMUX2X1_284 BUFX4_317/Y INVX1_411/Y NOR2X1_83/B gnd MUX2X1_284/Y vdd MUX2X1
XMUX2X1_273 BUFX4_421/Y INVX1_303/Y NOR2X1_70/Y gnd MUX2X1_273/Y vdd MUX2X1
XMUX2X1_262 OAI22X1_77/Y MUX2X1_262/B BUFX4_418/Y gnd OAI22X1_80/C vdd MUX2X1
XMUX2X1_251 MUX2X1_251/A MUX2X1_251/B BUFX4_74/Y gnd MUX2X1_251/Y vdd MUX2X1
XMUX2X1_295 BUFX4_430/Y INVX1_292/Y MUX2X1_55/S gnd MUX2X1_295/Y vdd MUX2X1
XFILL_48_3_1 gnd vdd FILL
XFILL_31_2_1 gnd vdd FILL
XCLKBUF1_15 BUFX4_9/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_37 BUFX4_8/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_26 BUFX4_6/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_48 BUFX4_5/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XCLKBUF1_59 BUFX4_8/Y gnd CLKBUF1_59/Y vdd CLKBUF1
XFILL_39_3_1 gnd vdd FILL
XBUFX4_80 BUFX4_75/A gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 BUFX4_75/A gnd BUFX4_91/Y vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 XNOR2X1_1/A XNOR2X1_1/B gnd INVX1_200/A vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XBUFX4_409 address[2] gnd INVX8_30/A vdd BUFX4
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XOAI21X1_581 BUFX4_148/Y OAI21X1_581/B BUFX4_342/Y gnd AOI21X1_263/C vdd OAI21X1
XOAI21X1_592 INVX1_251/Y BUFX4_261/Y NAND2X1_180/Y gnd MUX2X1_179/A vdd OAI21X1
XOAI21X1_570 INVX1_233/Y BUFX4_240/Y BUFX4_86/Y gnd OAI21X1_570/Y vdd OAI21X1
XAOI21X1_616 BUFX4_440/Y NOR2X1_729/B NOR2X1_728/Y gnd AOI21X1_616/Y vdd AOI21X1
XAOI21X1_605 BUFX4_72/Y NOR2X1_716/B NOR2X1_717/Y gnd AOI21X1_605/Y vdd AOI21X1
XAOI21X1_627 MUX2X1_4/B NOR2X1_737/B NOR2X1_739/Y gnd AOI21X1_627/Y vdd AOI21X1
XBUFX4_217 INVX8_11/Y gnd BUFX4_217/Y vdd BUFX4
XBUFX4_228 BUFX4_17/Y gnd AND2X2_37/B vdd BUFX4
XBUFX4_206 address[3] gnd BUFX4_206/Y vdd BUFX4
XBUFX4_239 BUFX4_19/Y gnd AND2X2_22/A vdd BUFX4
XFILL_45_1_1 gnd vdd FILL
XAND2X2_1 traffic_Street_1[0] traffic_Street_1[1] gnd AND2X2_1/Y vdd AND2X2
XOAI21X1_1129 BUFX4_222/Y NOR2X1_734/A AOI21X1_478/Y gnd OAI21X1_1131/C vdd OAI21X1
XOAI21X1_1118 BUFX4_327/Y OAI21X1_1348/C BUFX4_153/Y gnd OAI22X1_56/C vdd OAI21X1
XOAI21X1_1107 OAI22X1_52/Y BUFX4_391/Y INVX8_33/Y gnd OAI22X1_60/B vdd OAI21X1
XINVX1_420 INVX1_420/A gnd INVX1_420/Y vdd INVX1
XDFFPOSX1_708 OAI21X1_85/C CLKBUF1_35/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_719 INVX1_49/A CLKBUF1_38/Y MUX2X1_39/Y gnd vdd DFFPOSX1
XINVX1_431 INVX1_431/A gnd INVX1_431/Y vdd INVX1
XINVX1_453 INVX1_453/A gnd INVX1_453/Y vdd INVX1
XINVX1_442 INVX1_442/A gnd INVX1_442/Y vdd INVX1
XFILL_2_1 gnd vdd FILL
XFILL_51_2 gnd vdd FILL
XFILL_44_1 gnd vdd FILL
XFILL_36_1_1 gnd vdd FILL
XAOI21X1_424 BUFX4_413/Y MUX2X1_238/Y BUFX4_165/Y gnd AOI22X1_26/B vdd AOI21X1
XAOI21X1_413 BUFX4_393/Y MUX2X1_234/Y INVX8_33/Y gnd AOI22X1_25/B vdd AOI21X1
XAOI21X1_402 BUFX4_98/Y NOR2X1_700/A AOI21X1_402/C gnd OAI22X1_38/C vdd AOI21X1
XAOI21X1_446 BUFX4_51/Y AOI22X1_30/Y BUFX4_402/Y gnd AOI22X1_31/B vdd AOI21X1
XAOI21X1_435 BUFX4_265/Y INVX1_51/Y BUFX4_102/Y gnd AOI21X1_435/Y vdd AOI21X1
XAOI21X1_457 NOR2X1_216/A BUFX4_248/Y AOI21X1_457/C gnd AOI21X1_457/Y vdd AOI21X1
XAOI21X1_468 AND2X2_25/B INVX1_415/Y BUFX4_93/Y gnd AOI21X1_468/Y vdd AOI21X1
XAOI21X1_479 BUFX4_224/Y INVX1_425/Y AND2X2_33/B gnd AOI21X1_479/Y vdd AOI21X1
XNAND3X1_39 NAND3X1_39/A INVX1_198/A AOI22X1_4/Y gnd NAND3X1_39/Y vdd NAND3X1
XNAND3X1_28 INVX4_8/Y NAND3X1_6/C NAND3X1_28/C gnd NAND3X1_29/B vdd NAND3X1
XNAND3X1_17 INVX4_7/Y NAND3X1_17/B NAND3X1_17/C gnd NAND3X1_17/Y vdd NAND3X1
XNOR2X1_28 NOR2X1_28/A NOR2X1_30/B gnd AOI21X1_8/C vdd NOR2X1
XNOR2X1_17 NOR2X1_17/A NOR2X1_16/Y gnd NOR2X1_17/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_27_1_1 gnd vdd FILL
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B gnd NOR2X1_43/B vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XFILL_47_9_0 gnd vdd FILL
XMUX2X1_35 BUFX4_173/Y INVX1_43/Y NOR2X1_57/Y gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_24 INVX1_31/Y MUX2X1_8/B MUX2X1_21/S gnd MUX2X1_24/Y vdd MUX2X1
XMUX2X1_13 INVX1_18/Y MUX2X1_1/B MUX2X1_14/S gnd MUX2X1_13/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XNOR2X1_129 NOR2X1_129/A AOI21X1_72/B gnd AOI21X1_75/C vdd NOR2X1
XMUX2X1_46 BUFX4_217/Y INVX1_56/Y NOR2X1_85/B gnd MUX2X1_46/Y vdd MUX2X1
XNOR2X1_118 NOR2X1_118/A NAND2X1_50/B gnd NOR2X1_118/Y vdd NOR2X1
XMUX2X1_57 MUX2X1_57/A INVX1_67/Y MUX2X1_55/S gnd MUX2X1_57/Y vdd MUX2X1
XMUX2X1_68 INVX1_78/Y MUX2X1_77/B MUX2X1_70/S gnd MUX2X1_68/Y vdd MUX2X1
XMUX2X1_79 INVX1_89/Y MUX2X1_58/A MUX2X1_76/S gnd MUX2X1_79/Y vdd MUX2X1
XNOR2X1_107 NOR2X1_107/A NOR2X1_107/B gnd AOI21X1_59/C vdd NOR2X1
XFILL_30_8_0 gnd vdd FILL
XDFFPOSX1_505 NOR2X1_484/A CLKBUF1_18/Y DFFPOSX1_505/D gnd vdd DFFPOSX1
XDFFPOSX1_516 NAND2X1_242/B CLKBUF1_17/Y DFFPOSX1_516/D gnd vdd DFFPOSX1
XDFFPOSX1_538 OAI21X1_1527/C CLKBUF1_64/Y DFFPOSX1_538/D gnd vdd DFFPOSX1
XDFFPOSX1_527 MUX2X1_182/B CLKBUF1_67/Y DFFPOSX1_527/D gnd vdd DFFPOSX1
XINVX1_250 INVX1_250/A gnd INVX1_250/Y vdd INVX1
XDFFPOSX1_549 NOR2X1_732/A CLKBUF1_57/Y AOI21X1_620/Y gnd vdd DFFPOSX1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XINVX1_294 INVX1_294/A gnd INVX1_294/Y vdd INVX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XNAND2X1_50 traffic_Street_1[2] NAND2X1_50/B gnd NAND2X1_50/Y vdd NAND2X1
XNAND2X1_61 INVX8_21/A INVX4_4/Y gnd NAND2X1_61/Y vdd NAND2X1
XFILL_38_9_0 gnd vdd FILL
XNAND2X1_94 NAND2X1_94/A OAI21X1_7/B gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_83 INVX8_27/A INVX4_4/Y gnd MUX2X1_406/S vdd NAND2X1
XNAND2X1_72 INVX8_24/A INVX4_4/Y gnd NAND2X1_72/Y vdd NAND2X1
XNOR2X1_652 NOR2X1_652/A NOR2X1_97/B gnd NOR2X1_652/Y vdd NOR2X1
XNOR2X1_630 NOR2X1_630/A NOR2X1_60/Y gnd NOR2X1_630/Y vdd NOR2X1
XNOR2X1_641 NOR2X1_641/A NOR2X1_83/B gnd NOR2X1_641/Y vdd NOR2X1
XNOR2X1_696 NOR2X1_696/A MUX2X1_102/S gnd NOR2X1_696/Y vdd NOR2X1
XNOR2X1_674 NOR2X1_674/A NOR2X1_137/B gnd NOR2X1_674/Y vdd NOR2X1
XNOR2X1_663 NOR2X1_539/B NAND2X1_50/B gnd NOR2X1_663/Y vdd NOR2X1
XNOR2X1_685 NOR2X1_685/A NOR2X1_155/B gnd NOR2X1_685/Y vdd NOR2X1
XFILL_21_8_0 gnd vdd FILL
XAOI21X1_232 INVX2_24/Y NOR2X1_319/Y NOR3X1_11/Y gnd AND2X2_11/A vdd AOI21X1
XAOI21X1_243 NOR2X1_339/Y NOR3X1_13/Y AOI21X1_242/Y gnd AOI22X1_8/C vdd AOI21X1
XAOI21X1_210 NAND3X1_15/C OAI21X1_473/B INVX4_8/Y gnd NOR3X1_5/A vdd AOI21X1
XAOI21X1_221 NOR2X1_311/Y AOI21X1_221/B OR2X2_5/B gnd NAND3X1_43/C vdd AOI21X1
XAOI21X1_254 BUFX4_82/Y INVX1_229/Y NOR2X1_365/Y gnd OAI21X1_566/B vdd AOI21X1
XAOI21X1_265 AOI21X1_265/A AOI21X1_265/B AND2X2_48/B gnd AOI21X1_265/Y vdd AOI21X1
XAOI21X1_276 BUFX4_268/Y INVX1_258/Y AOI21X1_276/C gnd OAI21X1_601/B vdd AOI21X1
XAOI21X1_287 BUFX4_146/Y INVX1_271/Y OAI21X1_617/Y gnd AOI21X1_287/Y vdd AOI21X1
XAOI21X1_298 BUFX4_417/Y MUX2X1_197/Y AOI21X1_298/C gnd AOI21X1_299/C vdd AOI21X1
XOAI21X1_1460 NAND2X1_70/Y BUFX4_420/Y OAI21X1_1460/C gnd OAI21X1_1460/Y vdd OAI21X1
XOAI21X1_1493 BUFX4_457/Y BUFX4_298/Y NOR2X1_485/B gnd OAI21X1_1493/Y vdd OAI21X1
XOAI21X1_1482 BUFX4_445/Y NAND2X1_74/Y OAI21X1_1481/Y gnd OAI21X1_1482/Y vdd OAI21X1
XOAI21X1_1471 BUFX4_451/Y BUFX4_164/Y INVX1_431/A gnd OAI21X1_1471/Y vdd OAI21X1
XFILL_29_9_0 gnd vdd FILL
XFILL_4_9_0 gnd vdd FILL
XFILL_12_8_0 gnd vdd FILL
XDFFPOSX1_1001 AND2X2_47/A CLKBUF1_7/Y OAI21X1_285/Y gnd vdd DFFPOSX1
XDFFPOSX1_1034 NOR2X1_238/A CLKBUF1_34/Y AOI21X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_1023 INVX1_283/A CLKBUF1_16/Y OAI21X1_305/Y gnd vdd DFFPOSX1
XDFFPOSX1_1012 OAI21X1_895/A CLKBUF1_67/Y OAI21X1_299/Y gnd vdd DFFPOSX1
XDFFPOSX1_1045 INVX1_408/A CLKBUF1_64/Y OAI21X1_325/Y gnd vdd DFFPOSX1
XDFFPOSX1_1056 NOR2X1_252/A CLKBUF1_52/Y AOI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_302 NOR2X1_666/A CLKBUF1_90/Y AOI21X1_554/Y gnd vdd DFFPOSX1
XDFFPOSX1_313 NOR2X1_665/A CLKBUF1_17/Y AOI21X1_553/Y gnd vdd DFFPOSX1
XDFFPOSX1_346 INVX1_231/A CLKBUF1_96/Y MUX2X1_313/Y gnd vdd DFFPOSX1
XDFFPOSX1_324 NAND2X1_282/B CLKBUF1_16/Y OAI21X1_1347/Y gnd vdd DFFPOSX1
XDFFPOSX1_335 INVX1_298/A CLKBUF1_6/Y OAI21X1_1335/Y gnd vdd DFFPOSX1
XDFFPOSX1_368 INVX1_368/A CLKBUF1_50/Y MUX2X1_299/Y gnd vdd DFFPOSX1
XDFFPOSX1_379 NOR2X1_641/A CLKBUF1_13/Y AOI21X1_529/Y gnd vdd DFFPOSX1
XDFFPOSX1_357 AOI21X1_470/B CLKBUF1_55/Y OAI21X1_1330/Y gnd vdd DFFPOSX1
XNOR2X1_460 NOR2X1_460/A BUFX4_331/Y gnd NOR2X1_460/Y vdd NOR2X1
XNOR2X1_493 NOR2X1_35/A BUFX4_332/Y gnd NOR2X1_493/Y vdd NOR2X1
XNOR2X1_482 NOR2X1_721/A BUFX4_153/Y gnd NOR2X1_482/Y vdd NOR2X1
XNOR2X1_471 BUFX4_365/Y INVX1_347/Y gnd NOR2X1_471/Y vdd NOR2X1
XOAI21X1_900 OAI21X1_900/A BUFX4_240/Y BUFX4_82/Y gnd OAI22X1_33/B vdd OAI21X1
XOAI21X1_933 BUFX4_157/Y OAI21X1_933/B BUFX4_363/Y gnd NOR2X1_475/B vdd OAI21X1
XOAI21X1_922 INVX1_353/Y BUFX4_260/Y BUFX4_150/Y gnd OAI21X1_922/Y vdd OAI21X1
XOAI21X1_911 INVX1_342/Y BUFX4_246/Y OAI21X1_911/C gnd MUX2X1_228/B vdd OAI21X1
XOAI21X1_966 NOR2X1_484/Y NOR2X1_485/Y BUFX4_357/Y gnd AOI21X1_422/B vdd OAI21X1
XOAI21X1_944 MUX2X1_232/Y BUFX4_335/Y BUFX4_152/Y gnd AOI21X1_410/C vdd OAI21X1
XOAI21X1_955 INVX1_378/Y BUFX4_281/Y BUFX4_115/Y gnd OAI21X1_956/B vdd OAI21X1
XOAI21X1_977 INVX1_20/Y BUFX4_350/Y BUFX4_146/Y gnd OAI21X1_977/Y vdd OAI21X1
XOAI21X1_988 INVX1_392/Y BUFX4_241/Y OAI21X1_988/C gnd MUX2X1_240/B vdd OAI21X1
XOAI21X1_999 INVX1_118/Y BUFX4_96/Y BUFX4_345/Y gnd OAI21X1_999/Y vdd OAI21X1
XMUX2X1_411 MUX2X1_4/B INVX1_425/Y MUX2X1_410/S gnd MUX2X1_411/Y vdd MUX2X1
XMUX2X1_400 BUFX4_71/Y INVX1_389/Y MUX2X1_400/S gnd MUX2X1_400/Y vdd MUX2X1
XOAI21X1_1290 BUFX4_120/Y BUFX4_476/Y INVX1_225/A gnd OAI21X1_1291/C vdd OAI21X1
XDFFPOSX1_880 NOR2X1_155/A CLKBUF1_101/Y AOI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_891 INVX1_285/A CLKBUF1_45/Y OAI21X1_209/Y gnd vdd DFFPOSX1
XFILL_7_0_1 gnd vdd FILL
XFILL_44_7_0 gnd vdd FILL
XOAI21X1_15 OAI21X1_11/A BUFX4_64/Y OAI21X1_14/Y gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_26 OAI21X1_24/A MUX2X1_8/B OAI21X1_25/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_59 BUFX4_191/Y BUFX4_461/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_37 NOR2X1_39/A BUFX4_303/Y NOR2X1_438/A gnd OAI21X1_38/C vdd OAI21X1
XOAI21X1_48 BUFX4_70/Y OAI21X1_48/B OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XFILL_35_7_0 gnd vdd FILL
XOAI21X1_218 BUFX4_119/Y BUFX4_404/Y OAI21X1_846/A gnd OAI21X1_219/C vdd OAI21X1
XOAI21X1_207 BUFX4_465/Y NAND2X1_60/Y OAI21X1_207/C gnd OAI21X1_207/Y vdd OAI21X1
XOAI21X1_229 NAND2X1_64/Y BUFX4_377/Y OAI21X1_228/Y gnd OAI21X1_229/Y vdd OAI21X1
XAND2X2_18 AND2X2_18/A AND2X2_18/B gnd AND2X2_18/Y vdd AND2X2
XDFFPOSX1_121 NOR2X1_293/A CLKBUF1_4/Y AOI21X1_196/Y gnd vdd DFFPOSX1
XAND2X2_29 AND2X2_29/A AND2X2_29/B gnd AND2X2_29/Y vdd AND2X2
XDFFPOSX1_110 OAI21X1_413/C CLKBUF1_63/Y OAI21X1_414/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 INVX1_240/A CLKBUF1_86/Y MUX2X1_340/Y gnd vdd DFFPOSX1
XDFFPOSX1_143 OAI21X1_741/B CLKBUF1_24/Y DFFPOSX1_143/D gnd vdd DFFPOSX1
XDFFPOSX1_132 INVX1_186/A CLKBUF1_51/Y MUX2X1_172/Y gnd vdd DFFPOSX1
XDFFPOSX1_198 INVX1_242/A CLKBUF1_101/Y MUX2X1_339/Y gnd vdd DFFPOSX1
XDFFPOSX1_165 NOR2X1_628/A CLKBUF1_19/Y AOI21X1_516/Y gnd vdd DFFPOSX1
XNAND2X1_202 NOR2X1_286/A BUFX4_242/Y gnd NAND2X1_202/Y vdd NAND2X1
XDFFPOSX1_176 NAND2X1_281/B CLKBUF1_7/Y DFFPOSX1_176/D gnd vdd DFFPOSX1
XDFFPOSX1_187 OAI21X1_756/B CLKBUF1_45/Y OAI21X1_1401/Y gnd vdd DFFPOSX1
XNAND2X1_235 BUFX4_280/Y NOR2X1_667/A gnd NAND2X1_235/Y vdd NAND2X1
XNAND2X1_213 address[6] MUX2X1_199/Y gnd AOI22X1_18/D vdd NAND2X1
XNAND2X1_224 NAND2X1_224/A BUFX4_236/Y gnd NAND2X1_224/Y vdd NAND2X1
XNAND2X1_268 OAI21X1_306/C BUFX4_231/Y gnd NAND2X1_268/Y vdd NAND2X1
XNAND2X1_257 NAND2X1_257/A BUFX4_275/Y gnd OAI21X1_860/C vdd NAND2X1
XNAND2X1_246 BUFX4_171/Y NAND2X1_245/Y gnd NAND2X1_246/Y vdd NAND2X1
XNAND2X1_279 BUFX4_391/Y OAI22X1_37/Y gnd AOI22X1_24/C vdd NAND2X1
XFILL_26_7_0 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XNOR2X1_290 NOR2X1_290/A NOR2X1_43/B gnd NOR2X1_290/Y vdd NOR2X1
XOAI21X1_741 BUFX4_157/Y OAI21X1_741/B BUFX4_334/Y gnd NOR2X1_418/B vdd OAI21X1
XOAI21X1_730 OAI21X1_730/A NOR2X1_416/Y BUFX4_31/Y gnd AOI22X1_19/A vdd OAI21X1
XOAI21X1_763 BUFX4_413/Y OAI22X1_20/Y AOI21X1_336/Y gnd OAI21X1_770/C vdd OAI21X1
XOAI21X1_785 NOR2X1_432/Y NOR2X1_433/Y BUFX4_229/Y gnd AOI21X1_341/A vdd OAI21X1
XOAI21X1_752 BUFX4_271/Y OAI21X1_752/B BUFX4_115/Y gnd AOI21X1_330/C vdd OAI21X1
XOAI21X1_774 INVX1_317/Y BUFX4_290/Y OAI21X1_774/C gnd MUX2X1_212/B vdd OAI21X1
XOAI21X1_796 BUFX4_154/Y OAI21X1_796/B BUFX4_351/Y gnd AOI21X1_349/C vdd OAI21X1
XMUX2X1_241 MUX2X1_241/A MUX2X1_241/B BUFX4_98/Y gnd MUX2X1_241/Y vdd MUX2X1
XMUX2X1_230 MUX2X1_230/A MUX2X1_230/B BUFX4_415/Y gnd NOR2X1_479/B vdd MUX2X1
XMUX2X1_274 BUFX4_64/Y INVX1_360/Y NOR2X1_70/Y gnd MUX2X1_274/Y vdd MUX2X1
XMUX2X1_263 MUX2X1_263/A OAI22X1_83/Y BUFX4_411/Y gnd MUX2X1_263/Y vdd MUX2X1
XMUX2X1_252 MUX2X1_251/Y MUX2X1_250/Y INVX8_30/A gnd MUX2X1_252/Y vdd MUX2X1
XMUX2X1_296 BUFX4_70/Y INVX1_367/Y MUX2X1_55/S gnd MUX2X1_296/Y vdd MUX2X1
XMUX2X1_285 BUFX4_424/Y INVX1_299/Y NOR2X1_85/B gnd MUX2X1_285/Y vdd MUX2X1
XFILL_9_8_0 gnd vdd FILL
XFILL_17_7_0 gnd vdd FILL
XCLKBUF1_27 BUFX4_8/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_38 BUFX4_2/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XCLKBUF1_16 BUFX4_2/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_49 BUFX4_10/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XBUFX4_70 INVX8_4/Y gnd BUFX4_70/Y vdd BUFX4
XBUFX4_92 BUFX4_11/Y gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 BUFX4_11/Y gnd BUFX4_81/Y vdd BUFX4
XFILL_50_5_0 gnd vdd FILL
XXNOR2X1_2 AOI22X1_6/A INVX2_23/Y gnd AND2X2_9/A vdd XNOR2X1
XFILL_41_5_0 gnd vdd FILL
XINVX1_2 read_Write gnd INVX1_2/Y vdd INVX1
XOAI21X1_560 BUFX4_153/Y INVX1_225/Y AOI21X1_252/Y gnd OAI21X1_560/Y vdd OAI21X1
XOAI21X1_571 OAI21X1_570/Y AND2X2_22/Y OAI21X1_571/C gnd MUX2X1_178/B vdd OAI21X1
XOAI21X1_593 BUFX4_263/Y INVX1_252/Y AOI21X1_273/Y gnd OAI21X1_593/Y vdd OAI21X1
XOAI21X1_582 BUFX4_148/Y OAI21X1_582/B BUFX4_248/Y gnd AOI21X1_264/C vdd OAI21X1
XFILL_49_6_0 gnd vdd FILL
XFILL_32_5_0 gnd vdd FILL
XAOI21X1_606 BUFX4_318/Y NOR2X1_716/B NOR2X1_718/Y gnd AOI21X1_606/Y vdd AOI21X1
XAOI21X1_617 BUFX4_72/Y NOR2X1_729/B NOR2X1_729/Y gnd AOI21X1_617/Y vdd AOI21X1
XFILL_23_5_0 gnd vdd FILL
XFILL_6_6_0 gnd vdd FILL
XBUFX4_218 INVX8_11/Y gnd BUFX4_218/Y vdd BUFX4
XBUFX4_207 address[3] gnd BUFX4_207/Y vdd BUFX4
XBUFX4_229 BUFX4_18/Y gnd BUFX4_229/Y vdd BUFX4
XFILL_14_5_0 gnd vdd FILL
XOAI21X1_1119 BUFX4_289/Y OAI21X1_1119/B BUFX4_101/Y gnd OAI22X1_56/B vdd OAI21X1
XOAI21X1_1108 INVX1_420/Y BUFX4_280/Y BUFX4_151/Y gnd OAI21X1_1108/Y vdd OAI21X1
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XDFFPOSX1_709 OAI21X1_87/C CLKBUF1_94/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XOAI21X1_390 OAI21X1_24/A BUFX4_213/Y OAI21X1_389/Y gnd DFFPOSX1_90/D vdd OAI21X1
XINVX1_410 INVX1_410/A gnd INVX1_410/Y vdd INVX1
XINVX1_443 INVX1_443/A gnd INVX1_443/Y vdd INVX1
XINVX1_432 INVX1_432/A gnd INVX1_432/Y vdd INVX1
XINVX1_421 INVX1_421/A gnd INVX1_421/Y vdd INVX1
XINVX1_454 INVX1_454/A gnd INVX1_454/Y vdd INVX1
XFILL_2_2 gnd vdd FILL
XFILL_51_3 gnd vdd FILL
XFILL_37_1 gnd vdd FILL
XAOI21X1_425 INVX8_28/A AOI22X1_26/Y BUFX4_400/Y gnd AOI22X1_28/B vdd AOI21X1
XAOI21X1_403 BUFX4_50/Y OAI22X1_38/Y INVX8_33/Y gnd AOI22X1_24/D vdd AOI21X1
XAOI21X1_414 BUFX4_277/Y AOI21X1_414/B BUFX4_112/Y gnd OAI21X1_951/C vdd AOI21X1
XAOI21X1_447 BUFX4_111/Y AOI21X1_447/B NOR2X1_504/Y gnd AOI21X1_447/Y vdd AOI21X1
XAOI21X1_458 NOR2X1_253/A AND2X2_27/A BUFX4_83/Y gnd AOI21X1_458/Y vdd AOI21X1
XAOI21X1_436 INVX1_54/Y BUFX4_345/Y BUFX4_152/Y gnd AOI21X1_436/Y vdd AOI21X1
XAOI21X1_469 BUFX4_370/Y INVX1_416/Y BUFX4_156/Y gnd AOI21X1_469/Y vdd AOI21X1
XNAND3X1_29 NAND3X1_29/A NAND3X1_29/B NAND3X1_29/C gnd NOR3X1_8/C vdd NAND3X1
XNAND3X1_18 NOR2X1_351/B AND2X2_6/A NAND3X1_18/C gnd NAND3X1_19/C vdd NAND3X1
XNOR2X1_18 NOR2X1_18/A NOR2X1_16/Y gnd AOI21X1_2/C vdd NOR2X1
XNOR2X1_29 NOR2X1_29/A NOR2X1_30/B gnd NOR2X1_29/Y vdd NOR2X1
XFILL_47_9_1 gnd vdd FILL
XFILL_46_4_0 gnd vdd FILL
XMUX2X1_25 BUFX4_421/Y INVX1_33/Y NOR2X1_33/Y gnd MUX2X1_25/Y vdd MUX2X1
XMUX2X1_36 MUX2X1_82/B INVX1_44/Y NOR2X1_57/Y gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_14 INVX1_19/Y MUX2X1_6/B MUX2X1_14/S gnd MUX2X1_14/Y vdd MUX2X1
XMUX2X1_47 MUX2X1_49/A INVX1_57/Y NOR2X1_85/B gnd MUX2X1_47/Y vdd MUX2X1
XNOR2X1_119 NOR2X1_591/A NAND2X1_50/B gnd NOR2X1_119/Y vdd NOR2X1
XNOR2X1_108 NOR2X1_108/A NOR2X1_107/B gnd NOR2X1_108/Y vdd NOR2X1
XMUX2X1_69 INVX1_79/Y MUX2X1_61/B MUX2X1_70/S gnd MUX2X1_69/Y vdd MUX2X1
XMUX2X1_58 MUX2X1_58/A INVX1_68/Y MUX2X1_55/S gnd MUX2X1_58/Y vdd MUX2X1
XFILL_30_8_1 gnd vdd FILL
XDFFPOSX1_517 NAND2X1_286/B CLKBUF1_16/Y OAI21X1_1510/Y gnd vdd DFFPOSX1
XDFFPOSX1_506 NOR2X1_566/A CLKBUF1_79/Y OAI21X1_1504/Y gnd vdd DFFPOSX1
XDFFPOSX1_528 NAND2X1_244/A CLKBUF1_64/Y DFFPOSX1_528/D gnd vdd DFFPOSX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XINVX1_262 INVX1_262/A gnd INVX1_262/Y vdd INVX1
XDFFPOSX1_539 NOR2X1_728/A CLKBUF1_36/Y AOI21X1_616/Y gnd vdd DFFPOSX1
XINVX1_273 INVX1_273/A gnd INVX1_273/Y vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XINVX1_284 INVX1_284/A gnd INVX1_284/Y vdd INVX1
XNAND2X1_51 INVX8_19/A INVX8_6/A gnd NAND2X1_51/Y vdd NAND2X1
XNAND2X1_40 INVX8_17/A INVX4_4/Y gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_95 NAND2X1_95/A OAI21X1_7/B gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_84 INVX8_27/A INVX4_5/Y gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_73 INVX8_24/A INVX8_8/A gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_62 INVX8_21/A INVX4_5/Y gnd NAND2X1_62/Y vdd NAND2X1
XFILL_37_4_0 gnd vdd FILL
XFILL_38_9_1 gnd vdd FILL
XNOR2X1_620 INVX1_130/A BUFX4_359/Y gnd NOR2X1_620/Y vdd NOR2X1
XNOR2X1_642 NOR2X1_642/A NOR2X1_85/B gnd NOR2X1_642/Y vdd NOR2X1
XNOR2X1_631 NOR2X1_521/A NOR2X1_60/Y gnd NOR2X1_631/Y vdd NOR2X1
XNOR2X1_653 NOR2X1_653/A MUX2X1_75/S gnd NOR2X1_653/Y vdd NOR2X1
XNOR2X1_686 NOR2X1_686/A NOR2X1_155/B gnd NOR2X1_686/Y vdd NOR2X1
XNOR2X1_675 NOR2X1_427/B MUX2X1_89/S gnd NOR2X1_675/Y vdd NOR2X1
XNOR2X1_664 NOR2X1_423/A MUX2X1_320/S gnd NOR2X1_664/Y vdd NOR2X1
XAOI21X1_200 BUFX4_470/Y NOR2X1_47/B NOR2X1_297/Y gnd AOI21X1_200/Y vdd AOI21X1
XNOR2X1_697 NOR2X1_697/A MUX2X1_108/S gnd NOR2X1_697/Y vdd NOR2X1
XAOI21X1_233 AND2X2_11/Y NOR2X1_334/Y INVX1_208/A gnd NAND3X1_58/A vdd AOI21X1
XAOI21X1_222 NAND3X1_34/Y OAI21X1_475/Y BUFX2_3/A gnd NAND3X1_35/B vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XFILL_21_8_1 gnd vdd FILL
XAOI21X1_211 traffic_Street_0[0] traffic_Street_0[1] traffic_Street_0[2] gnd NOR2X1_308/B
+ vdd AOI21X1
XAOI21X1_244 INVX2_26/Y INVX4_12/Y OAI21X1_536/Y gnd AOI21X1_244/Y vdd AOI21X1
XAOI21X1_255 BUFX4_413/Y AOI21X1_255/B BUFX4_201/Y gnd AOI22X1_12/C vdd AOI21X1
XAOI21X1_266 BUFX4_204/Y OAI22X1_4/Y AOI21X1_265/Y gnd MUX2X1_180/B vdd AOI21X1
XAOI21X1_277 BUFX4_369/Y INVX1_259/Y OAI21X1_602/Y gnd OAI21X1_604/A vdd AOI21X1
XAOI21X1_288 OAI21X1_615/Y OAI21X1_618/Y BUFX4_201/Y gnd AOI21X1_288/Y vdd AOI21X1
XAOI21X1_299 BUFX4_171/Y MUX2X1_196/Y AOI21X1_299/C gnd OAI22X1_8/C vdd AOI21X1
XOAI21X1_1450 BUFX4_384/Y BUFX4_431/Y OAI21X1_958/B gnd OAI21X1_1451/C vdd OAI21X1
XOAI21X1_1472 NAND2X1_72/Y BUFX4_320/Y OAI21X1_1471/Y gnd DFFPOSX1_482/D vdd OAI21X1
XOAI21X1_1483 BUFX4_192/Y BUFX4_164/Y NOR2X1_431/A gnd OAI21X1_1484/C vdd OAI21X1
XOAI21X1_1461 BUFX4_126/Y BUFX4_431/Y OAI21X1_961/B gnd OAI21X1_1461/Y vdd OAI21X1
XOAI21X1_1494 NAND2X1_75/Y BUFX4_72/Y OAI21X1_1493/Y gnd OAI21X1_1494/Y vdd OAI21X1
XFILL_4_9_1 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XFILL_28_4_0 gnd vdd FILL
XFILL_29_9_1 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_12_8_1 gnd vdd FILL
XDFFPOSX1_1002 NOR2X1_616/A CLKBUF1_7/Y OAI21X1_287/Y gnd vdd DFFPOSX1
XDFFPOSX1_1024 OAI21X1_306/C CLKBUF1_56/Y OAI21X1_307/Y gnd vdd DFFPOSX1
XDFFPOSX1_1035 NOR2X1_381/A CLKBUF1_36/Y OAI21X1_313/Y gnd vdd DFFPOSX1
XDFFPOSX1_1013 NOR2X1_517/A CLKBUF1_36/Y OAI21X1_301/Y gnd vdd DFFPOSX1
XDFFPOSX1_1057 NOR2X1_253/A CLKBUF1_57/Y AOI21X1_162/Y gnd vdd DFFPOSX1
XDFFPOSX1_1046 AOI21X1_510/A CLKBUF1_60/Y OAI21X1_327/Y gnd vdd DFFPOSX1
XFILL_19_4_0 gnd vdd FILL
XDFFPOSX1_303 NOR2X1_667/A CLKBUF1_56/Y AOI21X1_555/Y gnd vdd DFFPOSX1
XDFFPOSX1_314 NOR2X1_642/A CLKBUF1_97/Y AOI21X1_530/Y gnd vdd DFFPOSX1
XDFFPOSX1_325 OAI21X1_1348/C CLKBUF1_16/Y DFFPOSX1_325/D gnd vdd DFFPOSX1
XDFFPOSX1_347 INVX1_295/A CLKBUF1_87/Y MUX2X1_314/Y gnd vdd DFFPOSX1
XDFFPOSX1_336 INVX1_343/A CLKBUF1_99/Y OAI21X1_1337/Y gnd vdd DFFPOSX1
XDFFPOSX1_369 INVX1_416/A CLKBUF1_95/Y MUX2X1_300/Y gnd vdd DFFPOSX1
XDFFPOSX1_358 INVX1_230/A CLKBUF1_87/Y MUX2X1_305/Y gnd vdd DFFPOSX1
XBUFX4_390 INVX8_28/Y gnd BUFX4_390/Y vdd BUFX4
XNOR2X1_461 INVX1_124/A BUFX4_237/Y gnd NOR2X1_461/Y vdd NOR2X1
XNOR2X1_450 BUFX4_413/Y NOR2X1_450/B gnd OAI22X1_28/A vdd NOR2X1
XNOR2X1_472 BUFX4_354/Y INVX1_352/Y gnd NOR2X1_472/Y vdd NOR2X1
XNOR2X1_494 NOR2X1_494/A BUFX4_244/Y gnd NOR2X1_494/Y vdd NOR2X1
XNOR2X1_483 BUFX4_74/Y NOR2X1_483/B gnd NOR2X1_483/Y vdd NOR2X1
XOAI21X1_934 AND2X2_32/B NOR2X1_626/A AOI21X1_405/Y gnd NAND3X1_76/B vdd OAI21X1
XOAI21X1_923 OAI21X1_922/Y NOR2X1_472/Y BUFX4_39/Y gnd OAI22X1_37/A vdd OAI21X1
XOAI21X1_912 INVX1_343/Y BUFX4_248/Y NAND2X1_272/Y gnd MUX2X1_228/A vdd OAI21X1
XOAI21X1_901 OAI22X1_33/Y BUFX4_33/Y BUFX4_166/Y gnd OAI22X1_36/A vdd OAI21X1
XOAI21X1_956 NOR2X1_481/Y OAI21X1_956/B OAI21X1_956/C gnd MUX2X1_235/A vdd OAI21X1
XOAI21X1_967 INVX1_385/Y AND2X2_46/B NAND2X1_288/Y gnd MUX2X1_237/B vdd OAI21X1
XOAI21X1_945 NOR2X1_479/Y OAI21X1_942/Y NOR2X1_480/Y gnd AOI22X1_25/A vdd OAI21X1
XOAI21X1_978 OAI21X1_977/Y NOR2X1_489/Y BUFX4_414/Y gnd OAI21X1_981/B vdd OAI21X1
XOAI21X1_989 INVX1_39/Y AND2X2_47/B OAI21X1_989/C gnd MUX2X1_240/A vdd OAI21X1
XMUX2X1_401 BUFX4_441/Y INVX1_269/Y NOR2X1_261/B gnd MUX2X1_401/Y vdd MUX2X1
XOAI21X1_1280 NAND2X1_31/Y MUX2X1_4/B OAI21X1_1279/Y gnd DFFPOSX1_149/D vdd OAI21X1
XOAI21X1_1291 NAND2X1_36/Y BUFX4_440/Y OAI21X1_1291/C gnd DFFPOSX1_230/D vdd OAI21X1
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XDFFPOSX1_870 NOR2X1_144/A CLKBUF1_93/Y AOI21X1_85/Y gnd vdd DFFPOSX1
XDFFPOSX1_881 MUX2X1_247/B CLKBUF1_44/Y AOI21X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_892 NOR2X1_447/A CLKBUF1_33/Y OAI21X1_211/Y gnd vdd DFFPOSX1
XFILL_44_7_1 gnd vdd FILL
XFILL_43_2_0 gnd vdd FILL
XOAI21X1_16 BUFX4_295/Y BUFX4_299/Y OAI21X1_16/C gnd OAI21X1_17/C vdd OAI21X1
XOAI21X1_27 BUFX4_125/Y BUFX4_293/Y INVX1_274/A gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_38 OAI21X1_40/A MUX2X1_27/B OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_49 BUFX4_62/Y NOR2X1_39/A AND2X2_51/A gnd OAI21X1_50/C vdd OAI21X1
XFILL_35_7_1 gnd vdd FILL
XFILL_34_2_0 gnd vdd FILL
XOAI21X1_219 NAND2X1_62/Y BUFX4_174/Y OAI21X1_219/C gnd OAI21X1_219/Y vdd OAI21X1
XOAI21X1_208 BUFX4_452/Y BUFX4_403/Y INVX1_285/A gnd OAI21X1_209/C vdd OAI21X1
XAND2X2_19 AND2X2_18/Y INVX4_9/A gnd AND2X2_19/Y vdd AND2X2
XDFFPOSX1_100 OAI21X1_401/C CLKBUF1_84/Y OAI21X1_402/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 AND2X2_36/A CLKBUF1_88/Y OAI21X1_416/Y gnd vdd DFFPOSX1
XDFFPOSX1_144 OAI21X1_933/B CLKBUF1_76/Y OAI21X1_1286/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 INVX1_281/A CLKBUF1_99/Y OAI21X1_422/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 NOR2X1_298/A CLKBUF1_99/Y AOI21X1_201/Y gnd vdd DFFPOSX1
XDFFPOSX1_155 NOR2X1_687/A CLKBUF1_71/Y AOI21X1_575/Y gnd vdd DFFPOSX1
XDFFPOSX1_166 NOR2X1_678/A CLKBUF1_69/Y AOI21X1_566/Y gnd vdd DFFPOSX1
XDFFPOSX1_188 MUX2X1_231/B CLKBUF1_74/Y OAI21X1_1403/Y gnd vdd DFFPOSX1
XDFFPOSX1_177 NOR2X1_536/B CLKBUF1_45/Y OAI21X1_1413/Y gnd vdd DFFPOSX1
XNAND2X1_214 OAI21X1_184/C AND2X2_41/A gnd NAND2X1_214/Y vdd NAND2X1
XNAND2X1_203 NOR2X1_275/A BUFX4_244/Y gnd OAI21X1_648/C vdd NAND2X1
XDFFPOSX1_199 NOR2X1_684/A CLKBUF1_45/Y AOI21X1_572/Y gnd vdd DFFPOSX1
XNAND2X1_225 NOR2X1_92/A AND2X2_51/B gnd OAI21X1_711/C vdd NAND2X1
XNAND2X1_258 NOR2X1_137/A BUFX4_111/Y gnd NAND2X1_258/Y vdd NAND2X1
XNAND2X1_269 NOR2X1_236/A BUFX4_233/Y gnd OAI21X1_893/C vdd NAND2X1
XNAND2X1_236 BUFX4_282/Y INVX1_456/A gnd OAI21X1_762/C vdd NAND2X1
XNAND2X1_247 NOR2X1_62/A BUFX4_248/Y gnd NAND2X1_247/Y vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_26_7_1 gnd vdd FILL
XNOR2X1_280 NOR2X1_280/A AOI21X1_7/B gnd NOR2X1_280/Y vdd NOR2X1
XNOR2X1_291 NOR2X1_291/A NOR2X1_43/B gnd NOR2X1_291/Y vdd NOR2X1
XOAI21X1_742 BUFX4_157/Y NOR2X1_630/A AND2X2_23/A gnd OAI21X1_742/Y vdd OAI21X1
XOAI21X1_731 BUFX4_253/Y INVX1_297/Y OAI21X1_731/C gnd OAI21X1_733/C vdd OAI21X1
XOAI21X1_720 INVX1_81/A BUFX4_244/Y BUFX4_98/Y gnd OAI22X1_19/B vdd OAI21X1
XOAI21X1_764 BUFX4_361/Y NOR2X1_670/A BUFX4_154/Y gnd OAI22X1_21/C vdd OAI21X1
XOAI21X1_753 INVX1_309/Y BUFX4_274/Y NAND2X1_233/Y gnd OAI21X1_753/Y vdd OAI21X1
XOAI21X1_775 INVX1_318/Y AND2X2_46/B NAND2X1_240/Y gnd MUX2X1_212/A vdd OAI21X1
XOAI21X1_797 BUFX4_146/Y OAI21X1_797/B BUFX4_237/Y gnd OAI21X1_797/Y vdd OAI21X1
XOAI21X1_786 NOR2X1_434/Y NOR2X1_435/Y BUFX4_357/Y gnd AOI21X1_341/B vdd OAI21X1
XMUX2X1_220 MUX2X1_220/A MUX2X1_220/B BUFX4_325/Y gnd MUX2X1_221/B vdd MUX2X1
XMUX2X1_231 NOR2X1_691/A MUX2X1_231/B BUFX4_416/Y gnd MUX2X1_231/Y vdd MUX2X1
XMUX2X1_253 MUX2X1_253/A MUX2X1_252/Y BUFX4_202/Y gnd MUX2X1_253/Y vdd MUX2X1
XMUX2X1_242 OAI22X1_44/Y MUX2X1_242/B BUFX4_394/Y gnd MUX2X1_242/Y vdd MUX2X1
XMUX2X1_264 MUX2X1_264/A MUX2X1_264/B BUFX4_414/Y gnd OAI22X1_91/C vdd MUX2X1
XMUX2X1_297 INVX1_449/Y BUFX4_437/Y MUX2X1_59/S gnd MUX2X1_297/Y vdd MUX2X1
XMUX2X1_275 INVX1_220/Y AND2X2_5/B MUX2X1_42/S gnd MUX2X1_275/Y vdd MUX2X1
XFILL_9_8_1 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XMUX2X1_286 BUFX4_63/Y INVX1_349/Y NOR2X1_85/B gnd MUX2X1_286/Y vdd MUX2X1
XFILL_16_2_0 gnd vdd FILL
XFILL_17_7_1 gnd vdd FILL
XCLKBUF1_28 BUFX4_7/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_17 BUFX4_5/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XCLKBUF1_39 BUFX4_9/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XBUFX4_71 INVX8_4/Y gnd BUFX4_71/Y vdd BUFX4
XBUFX4_60 INVX8_6/Y gnd BUFX4_60/Y vdd BUFX4
XBUFX4_93 BUFX4_82/A gnd BUFX4_93/Y vdd BUFX4
XBUFX4_82 BUFX4_82/A gnd BUFX4_82/Y vdd BUFX4
XFILL_50_5_1 gnd vdd FILL
XOR2X2_1 traffic_Street_1[1] traffic_Street_1[2] gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 INVX4_12/A INVX2_23/A gnd AND2X2_9/B vdd XNOR2X1
XFILL_41_5_1 gnd vdd FILL
XINVX8_30 INVX8_30/A gnd BUFX4_33/A vdd INVX8
XFILL_40_0_0 gnd vdd FILL
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_550 INVX2_1/Y BUFX4_189/Y OAI21X1_550/C gnd OAI21X1_550/Y vdd OAI21X1
XOAI21X1_561 INVX1_226/Y BUFX4_79/Y AND2X2_37/B gnd OAI21X1_562/B vdd OAI21X1
XOAI21X1_583 OAI21X1_583/A OAI21X1_583/B BUFX4_40/Y gnd AOI21X1_265/B vdd OAI21X1
XOAI21X1_572 INVX1_234/Y BUFX4_241/Y BUFX4_87/Y gnd AOI21X1_260/C vdd OAI21X1
XOAI21X1_594 INVX1_253/Y BUFX4_265/Y BUFX4_95/Y gnd OAI21X1_595/A vdd OAI21X1
XFILL_49_6_1 gnd vdd FILL
XFILL_48_1_0 gnd vdd FILL
XFILL_32_5_1 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XAOI21X1_607 BUFX4_445/Y NOR2X1_231/B NOR2X1_719/Y gnd AOI21X1_607/Y vdd AOI21X1
XAOI21X1_618 BUFX4_439/Y NOR2X1_733/B NOR2X1_730/Y gnd AOI21X1_618/Y vdd AOI21X1
XFILL_39_1_0 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XBUFX4_208 INVX8_11/Y gnd AND2X2_2/B vdd BUFX4
XFILL_6_6_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XBUFX4_219 BUFX4_23/Y gnd AND2X2_46/B vdd BUFX4
XFILL_13_0_0 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XOAI21X1_1109 OAI21X1_1108/Y NOR2X1_531/Y BUFX4_40/Y gnd AOI21X1_473/C vdd OAI21X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XINVX1_411 INVX1_411/A gnd INVX1_411/Y vdd INVX1
XOAI21X1_391 BUFX4_450/Y NOR2X1_16/A NOR2X1_451/A gnd OAI21X1_392/C vdd OAI21X1
XOAI21X1_380 BUFX4_292/Y BUFX4_303/Y INVX1_280/A gnd OAI21X1_380/Y vdd OAI21X1
XINVX1_400 INVX1_400/A gnd INVX1_400/Y vdd INVX1
XINVX1_444 INVX1_444/A gnd INVX1_444/Y vdd INVX1
XINVX1_422 INVX1_422/A gnd INVX1_422/Y vdd INVX1
XINVX1_433 INVX1_433/A gnd INVX1_433/Y vdd INVX1
XINVX1_455 INVX1_455/A gnd INVX1_455/Y vdd INVX1
XAOI21X1_415 NOR2X1_709/A BUFX4_355/Y BUFX4_114/Y gnd OAI21X1_954/C vdd AOI21X1
XAOI21X1_404 BUFX4_101/Y INVX1_360/Y BUFX4_333/Y gnd OAI21X1_932/C vdd AOI21X1
XAOI21X1_437 INVX1_398/Y BUFX4_351/Y AOI21X1_437/C gnd AOI21X1_437/Y vdd AOI21X1
XAOI21X1_426 BUFX4_230/Y INVX1_391/Y BUFX4_79/Y gnd OAI21X1_973/C vdd AOI21X1
XAOI21X1_459 NOR2X1_243/A BUFX4_259/Y AOI21X1_459/C gnd NOR2X1_520/A vdd AOI21X1
XAOI21X1_448 NOR2X1_296/A BUFX4_290/Y BUFX4_113/Y gnd AOI21X1_448/Y vdd AOI21X1
XNAND3X1_19 INVX2_14/A NAND3X1_19/B NAND3X1_19/C gnd AND2X2_7/B vdd NAND3X1
XNOR2X1_19 NOR2X1_19/A NOR2X1_16/Y gnd AOI21X1_3/C vdd NOR2X1
XFILL_46_4_1 gnd vdd FILL
XMUX2X1_15 INVX1_20/Y BUFX4_71/Y MUX2X1_14/S gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_26 INVX1_34/Y BUFX4_443/Y MUX2X1_29/S gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_59 INVX1_69/Y MUX2X1_59/B MUX2X1_59/S gnd MUX2X1_59/Y vdd MUX2X1
XMUX2X1_37 MUX2X1_40/B INVX1_45/Y NOR2X1_70/Y gnd MUX2X1_37/Y vdd MUX2X1
XNOR2X1_109 NOR2X1_109/A NOR2X1_107/B gnd NOR2X1_109/Y vdd NOR2X1
XMUX2X1_48 BUFX4_381/Y INVX1_58/Y NOR2X1_85/B gnd MUX2X1_48/Y vdd MUX2X1
XDFFPOSX1_518 NAND2X1_338/B CLKBUF1_62/Y OAI21X1_1512/Y gnd vdd DFFPOSX1
XDFFPOSX1_529 INVX1_385/A CLKBUF1_60/Y OAI21X1_1518/Y gnd vdd DFFPOSX1
XDFFPOSX1_507 NOR2X1_719/A CLKBUF1_67/Y AOI21X1_607/Y gnd vdd DFFPOSX1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XINVX1_252 INVX1_252/A gnd INVX1_252/Y vdd INVX1
XINVX1_274 INVX1_274/A gnd INVX1_274/Y vdd INVX1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XINVX1_285 INVX1_285/A gnd INVX1_285/Y vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XNAND2X1_30 INVX8_12/A INVX4_2/Y gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_52 INVX8_19/A INVX4_3/Y gnd NAND2X1_52/Y vdd NAND2X1
XNAND2X1_41 INVX8_17/A INVX4_5/Y gnd MUX2X1_59/S vdd NAND2X1
XNAND2X1_85 INVX8_27/A INVX8_9/A gnd NAND2X1_85/Y vdd NAND2X1
XNAND2X1_74 INVX8_24/A INVX8_9/A gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_63 INVX8_22/A INVX4_2/Y gnd MUX2X1_97/S vdd NAND2X1
XFILL_37_4_1 gnd vdd FILL
XNAND2X1_96 NAND2X1_96/A OAI21X1_7/B gnd NAND2X1_96/Y vdd NAND2X1
XNOR2X1_610 NOR2X1_610/A BUFX4_237/Y gnd OAI22X1_85/D vdd NOR2X1
XNOR2X1_632 NOR2X1_632/A NOR2X1_65/Y gnd NOR2X1_632/Y vdd NOR2X1
XNOR2X1_643 NOR2X1_643/A MUX2X1_50/S gnd NOR2X1_643/Y vdd NOR2X1
XNOR2X1_621 NOR2X1_621/A BUFX4_247/Y gnd NOR2X1_621/Y vdd NOR2X1
XNOR2X1_676 NOR2X1_676/A MUX2X1_89/S gnd NOR2X1_676/Y vdd NOR2X1
XNOR2X1_665 NOR2X1_665/A MUX2X1_320/S gnd NOR2X1_665/Y vdd NOR2X1
XNOR2X1_654 NOR2X1_654/A MUX2X1_75/S gnd NOR2X1_654/Y vdd NOR2X1
XNOR2X1_687 NOR2X1_687/A MUX2X1_340/S gnd NOR2X1_687/Y vdd NOR2X1
XNOR2X1_698 NOR2X1_698/A INVX1_219/A gnd NOR2X1_698/Y vdd NOR2X1
XAOI21X1_212 INVX2_17/Y AOI21X1_212/B OAI21X1_461/Y gnd OAI21X1_462/C vdd AOI21X1
XAOI21X1_234 OAI21X1_507/Y AOI21X1_234/B NOR3X1_11/Y gnd NOR3X1_12/A vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_201 BUFX4_470/Y MUX2X1_31/S NOR2X1_298/Y gnd AOI21X1_201/Y vdd AOI21X1
XAOI21X1_223 INVX1_189/A NOR3X1_4/B OAI21X1_476/Y gnd NAND3X1_36/B vdd AOI21X1
XAOI21X1_245 NAND3X1_66/Y AOI21X1_244/Y AOI21X1_245/C gnd AND2X2_18/A vdd AOI21X1
XAOI21X1_267 BUFX4_250/Y NOR2X1_671/A AOI21X1_267/C gnd OAI22X1_5/B vdd AOI21X1
XAOI21X1_256 BUFX4_236/Y INVX1_231/Y OAI21X1_568/Y gnd AOI21X1_257/C vdd AOI21X1
XAOI21X1_289 NAND2X1_11/A BUFX4_288/Y OAI21X1_619/Y gnd AOI21X1_289/Y vdd AOI21X1
XAOI21X1_278 BUFX4_270/Y INVX1_260/Y AOI21X1_278/C gnd OAI21X1_604/B vdd AOI21X1
XOAI21X1_1440 BUFX4_60/Y BUFX4_435/Y NAND2X1_239/B gnd OAI21X1_1440/Y vdd OAI21X1
XOAI21X1_1473 BUFX4_135/Y BUFX4_160/Y AOI21X1_273/B gnd OAI21X1_1473/Y vdd OAI21X1
XOAI21X1_1484 BUFX4_422/Y NAND2X1_74/Y OAI21X1_1484/C gnd DFFPOSX1_492/D vdd OAI21X1
XOAI21X1_1451 NAND2X1_69/Y BUFX4_68/Y OAI21X1_1451/C gnd DFFPOSX1_292/D vdd OAI21X1
XOAI21X1_1462 NAND2X1_70/Y BUFX4_68/Y OAI21X1_1461/Y gnd DFFPOSX1_457/D vdd OAI21X1
XOAI21X1_1495 BUFX4_456/Y BUFX4_298/Y NOR2X1_567/B gnd OAI21X1_1496/C vdd OAI21X1
XFILL_28_4_1 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XFILL_11_3_1 gnd vdd FILL
XDFFPOSX1_1025 NAND2X1_329/A CLKBUF1_16/Y OAI21X1_309/Y gnd vdd DFFPOSX1
XDFFPOSX1_1036 INVX1_341/A CLKBUF1_60/Y OAI21X1_315/Y gnd vdd DFFPOSX1
XDFFPOSX1_1003 NOR2X1_383/A CLKBUF1_60/Y OAI21X1_289/Y gnd vdd DFFPOSX1
XDFFPOSX1_1014 OAI21X1_302/C CLKBUF1_18/Y OAI21X1_303/Y gnd vdd DFFPOSX1
XDFFPOSX1_1047 NOR2X1_246/A CLKBUF1_36/Y AOI21X1_156/Y gnd vdd DFFPOSX1
XOAI22X1_1 XOR2X1_3/A INVX2_22/A XNOR2X1_4/A INVX2_21/A gnd OAI22X1_1/Y vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XDFFPOSX1_304 NOR2X1_668/A CLKBUF1_97/Y AOI21X1_556/Y gnd vdd DFFPOSX1
XDFFPOSX1_315 INVX1_299/A CLKBUF1_92/Y MUX2X1_285/Y gnd vdd DFFPOSX1
XDFFPOSX1_326 INVX1_248/A CLKBUF1_42/Y OAI21X1_1340/Y gnd vdd DFFPOSX1
XDFFPOSX1_337 OAI21X1_1096/B CLKBUF1_58/Y OAI21X1_1339/Y gnd vdd DFFPOSX1
XDFFPOSX1_359 INVX1_294/A CLKBUF1_47/Y MUX2X1_306/Y gnd vdd DFFPOSX1
XDFFPOSX1_348 NOR2X1_653/A CLKBUF1_78/Y AOI21X1_541/Y gnd vdd DFFPOSX1
XBUFX4_391 INVX8_28/Y gnd BUFX4_391/Y vdd BUFX4
XBUFX4_380 INVX8_14/Y gnd BUFX4_380/Y vdd BUFX4
XNOR2X1_451 NOR2X1_451/A BUFX4_280/Y gnd NOR2X1_451/Y vdd NOR2X1
XNOR2X1_440 NOR2X1_440/A BUFX4_244/Y gnd OAI22X1_23/D vdd NOR2X1
XNOR2X1_462 NOR2X1_188/A BUFX4_359/Y gnd OAI22X1_32/A vdd NOR2X1
XNOR2X1_473 BUFX4_170/Y NOR2X1_473/B gnd OAI22X1_42/A vdd NOR2X1
XNOR2X1_484 NOR2X1_484/A BUFX4_155/Y gnd NOR2X1_484/Y vdd NOR2X1
XNOR2X1_495 NOR2X1_42/A BUFX4_355/Y gnd OAI22X1_41/A vdd NOR2X1
XOAI21X1_902 BUFX4_341/Y NOR2X1_207/A BUFX4_147/Y gnd OAI22X1_34/C vdd OAI21X1
XOAI21X1_924 BUFX4_356/Y OAI21X1_924/B BUFX4_150/Y gnd AOI21X1_399/C vdd OAI21X1
XOAI21X1_913 INVX1_344/Y BUFX4_250/Y NAND2X1_274/Y gnd MUX2X1_229/B vdd OAI21X1
XOAI21X1_957 BUFX4_348/Y OAI21X1_957/B BUFX4_147/Y gnd OAI21X1_957/Y vdd OAI21X1
XOAI21X1_935 AND2X2_33/B OAI21X1_935/B AOI21X1_406/Y gnd NAND3X1_76/C vdd OAI21X1
XOAI21X1_946 INVX1_370/Y BUFX4_270/Y OAI21X1_946/C gnd AOI21X1_412/B vdd OAI21X1
XOAI21X1_979 INVX1_10/Y BUFX4_347/Y OAI21X1_979/C gnd NAND3X1_78/B vdd OAI21X1
XOAI21X1_968 INVX1_386/Y INVX8_31/A OAI21X1_968/C gnd MUX2X1_237/A vdd OAI21X1
XMUX2X1_402 MUX2X1_18/B INVX1_327/Y NOR2X1_261/B gnd MUX2X1_402/Y vdd MUX2X1
XOAI21X1_1270 NAND2X1_30/Y BUFX4_64/Y OAI21X1_1270/C gnd DFFPOSX1_240/D vdd OAI21X1
XOAI21X1_1281 BUFX4_125/Y BUFX4_43/Y OAI21X1_557/B gnd OAI21X1_1282/C vdd OAI21X1
XDFFPOSX1_860 INVX1_103/A CLKBUF1_34/Y MUX2X1_90/Y gnd vdd DFFPOSX1
XOAI21X1_1292 BUFX4_120/Y BUFX4_476/Y INVX1_300/A gnd OAI21X1_1293/C vdd OAI21X1
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XDFFPOSX1_871 NOR2X1_146/A CLKBUF1_2/Y AOI21X1_86/Y gnd vdd DFFPOSX1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XDFFPOSX1_893 MUX2X1_246/A CLKBUF1_7/Y OAI21X1_213/Y gnd vdd DFFPOSX1
XDFFPOSX1_882 NOR2X1_157/A CLKBUF1_33/Y AOI21X1_94/Y gnd vdd DFFPOSX1
XFILL_43_2_1 gnd vdd FILL
XOAI21X1_17 OAI21X1_11/A MUX2X1_8/B OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 NAND2X1_24/Y MUX2X1_1/B OAI21X1_27/Y gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_39 BUFX4_460/Y BUFX4_303/Y NOR2X1_494/A gnd OAI21X1_40/C vdd OAI21X1
XFILL_34_2_1 gnd vdd FILL
XOAI21X1_209 NAND2X1_61/Y AND2X2_2/B OAI21X1_209/C gnd OAI21X1_209/Y vdd OAI21X1
XDFFPOSX1_101 OAI21X1_403/C CLKBUF1_91/Y OAI21X1_404/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 AOI21X1_449/A CLKBUF1_51/Y OAI21X1_418/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 OAI21X1_1091/B CLKBUF1_35/Y DFFPOSX1_145/D gnd vdd DFFPOSX1
XDFFPOSX1_134 OAI21X1_429/C CLKBUF1_47/Y OAI21X1_430/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 INVX1_338/A CLKBUF1_99/Y OAI21X1_424/Y gnd vdd DFFPOSX1
XDFFPOSX1_178 INVX1_220/A CLKBUF1_101/Y MUX2X1_275/Y gnd vdd DFFPOSX1
XDFFPOSX1_167 NOR2X1_679/A CLKBUF1_93/Y AOI21X1_567/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 MUX2X1_232/A CLKBUF1_71/Y AOI21X1_576/Y gnd vdd DFFPOSX1
XDFFPOSX1_189 NOR2X1_534/A CLKBUF1_71/Y DFFPOSX1_189/D gnd vdd DFFPOSX1
XNAND2X1_215 NOR2X1_146/A BUFX4_281/Y gnd OAI21X1_684/C vdd NAND2X1
XNAND2X1_204 NOR2X1_279/A BUFX4_246/Y gnd NAND2X1_204/Y vdd NAND2X1
XNAND2X1_226 BUFX4_37/Y OAI22X1_19/Y gnd AOI21X1_316/A vdd NAND2X1
XNAND2X1_259 NAND2X1_259/A BUFX4_113/Y gnd OAI21X1_863/C vdd NAND2X1
XNAND2X1_248 BUFX4_393/Y MUX2X1_218/Y gnd AOI22X1_23/D vdd NAND2X1
XNAND2X1_237 BUFX4_287/Y NOR2X1_704/A gnd NAND2X1_237/Y vdd NAND2X1
XFILL_25_2_1 gnd vdd FILL
XNOR2X1_270 BUFX4_196/Y BUFX4_133/Y gnd MUX2X1_410/S vdd NOR2X1
XFILL_0_2_1 gnd vdd FILL
XNOR2X1_281 NOR2X1_281/A AOI21X1_7/B gnd NOR2X1_281/Y vdd NOR2X1
XNOR2X1_292 NOR2X1_292/A NOR2X1_43/B gnd NOR2X1_292/Y vdd NOR2X1
XOAI21X1_721 NOR2X1_411/Y BUFX4_392/Y OAI21X1_709/Y gnd MUX2X1_207/A vdd OAI21X1
XOAI21X1_732 INVX1_298/Y BUFX4_255/Y AND2X2_32/B gnd OAI21X1_733/A vdd OAI21X1
XOAI21X1_710 INVX1_61/Y BUFX4_237/Y NAND2X1_224/Y gnd MUX2X1_206/B vdd OAI21X1
XOAI21X1_743 BUFX4_157/Y NOR2X1_627/A BUFX4_352/Y gnd OAI21X1_743/Y vdd OAI21X1
XOAI21X1_765 BUFX4_285/Y OAI21X1_765/B BUFX4_74/Y gnd OAI22X1_21/B vdd OAI21X1
XOAI21X1_754 BUFX4_275/Y OAI21X1_754/B BUFX4_116/Y gnd AOI21X1_333/C vdd OAI21X1
XOAI21X1_776 BUFX4_341/Y NOR2X1_711/A BUFX4_147/Y gnd OAI22X1_22/C vdd OAI21X1
XOAI21X1_798 AOI21X1_349/Y AOI21X1_350/Y BUFX4_419/Y gnd OAI21X1_798/Y vdd OAI21X1
XOAI21X1_787 BUFX4_231/Y INVX1_322/Y AOI21X1_343/Y gnd OAI21X1_787/Y vdd OAI21X1
XMUX2X1_210 MUX2X1_210/A MUX2X1_210/B BUFX4_118/Y gnd MUX2X1_210/Y vdd MUX2X1
XMUX2X1_221 MUX2X1_221/A MUX2X1_221/B BUFX4_412/Y gnd MUX2X1_221/Y vdd MUX2X1
XMUX2X1_232 MUX2X1_232/A NOR2X1_685/A BUFX4_419/Y gnd MUX2X1_232/Y vdd MUX2X1
XMUX2X1_265 MUX2X1_265/A MUX2X1_265/B BUFX4_110/Y gnd MUX2X1_265/Y vdd MUX2X1
XMUX2X1_243 MUX2X1_243/A MUX2X1_243/B BUFX4_99/Y gnd NOR2X1_496/B vdd MUX2X1
XMUX2X1_254 MUX2X1_254/A MUX2X1_254/B BUFX4_80/Y gnd MUX2X1_254/Y vdd MUX2X1
XDFFPOSX1_690 NOR2X1_56/A CLKBUF1_31/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XMUX2X1_287 BUFX4_322/Y INVX1_413/Y NOR2X1_85/B gnd MUX2X1_287/Y vdd MUX2X1
XMUX2X1_276 INVX1_446/Y BUFX4_429/Y MUX2X1_42/S gnd MUX2X1_276/Y vdd MUX2X1
XMUX2X1_298 INVX1_450/Y MUX2X1_27/B MUX2X1_59/S gnd MUX2X1_298/Y vdd MUX2X1
XFILL_8_3_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XCLKBUF1_29 BUFX4_8/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XCLKBUF1_18 BUFX4_4/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XBUFX4_50 address[4] gnd BUFX4_50/Y vdd BUFX4
XBUFX4_61 INVX8_6/Y gnd BUFX4_61/Y vdd BUFX4
XBUFX4_94 BUFX4_87/A gnd BUFX4_94/Y vdd BUFX4
XBUFX4_83 BUFX4_85/A gnd BUFX4_83/Y vdd BUFX4
XBUFX4_72 INVX8_4/Y gnd BUFX4_72/Y vdd BUFX4
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 XNOR2X1_4/A XNOR2X1_4/B gnd XNOR2X1_4/Y vdd XNOR2X1
XINVX8_20 INVX8_20/A gnd INVX8_20/Y vdd INVX8
XINVX8_31 INVX8_31/A gnd BUFX4_28/A vdd INVX8
XFILL_40_0_1 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_10_9_0 gnd vdd FILL
XOAI21X1_540 AOI22X1_10/D AOI22X1_9/C NOR2X1_353/Y gnd AOI21X1_246/B vdd OAI21X1
XOAI21X1_573 INVX1_236/Y AND2X2_47/B BUFX4_151/Y gnd OAI21X1_573/Y vdd OAI21X1
XOAI21X1_584 INVX1_243/Y BUFX4_249/Y BUFX4_90/Y gnd AOI21X1_267/C vdd OAI21X1
XOAI21X1_562 AND2X2_21/Y OAI21X1_562/B OAI21X1_560/Y gnd OAI21X1_562/Y vdd OAI21X1
XOAI21X1_551 AND2X2_20/Y INVX2_3/Y INVX1_219/Y gnd OAI21X1_551/Y vdd OAI21X1
XOAI21X1_595 OAI21X1_595/A AND2X2_23/Y OAI21X1_593/Y gnd MUX2X1_181/B vdd OAI21X1
XFILL_48_1_1 gnd vdd FILL
XAOI21X1_608 BUFX4_429/Y NOR2X1_231/B NOR2X1_720/Y gnd AOI21X1_608/Y vdd AOI21X1
XFILL_31_0_1 gnd vdd FILL
XAOI21X1_619 BUFX4_424/Y NOR2X1_733/B NOR2X1_731/Y gnd AOI21X1_619/Y vdd AOI21X1
XFILL_39_1_1 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XBUFX4_209 INVX8_11/Y gnd BUFX4_209/Y vdd BUFX4
XFILL_5_1_1 gnd vdd FILL
XFILL_42_8_0 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_392 OAI21X1_24/A BUFX4_178/Y OAI21X1_392/C gnd DFFPOSX1_91/D vdd OAI21X1
XOAI21X1_370 BUFX4_375/Y NAND2X1_2/Y NAND2X1_88/Y gnd OAI21X1_370/Y vdd OAI21X1
XOAI21X1_381 OAI21X1_11/A BUFX4_209/Y OAI21X1_380/Y gnd OAI21X1_381/Y vdd OAI21X1
XINVX1_401 INVX1_401/A gnd INVX1_401/Y vdd INVX1
XAND2X2_4 traffic_Street_0[0] traffic_Street_0[1] gnd AND2X2_4/Y vdd AND2X2
XINVX1_434 INVX1_434/A gnd INVX1_434/Y vdd INVX1
XINVX1_423 INVX1_423/A gnd INVX1_423/Y vdd INVX1
XINVX1_412 INVX1_412/A gnd INVX1_412/Y vdd INVX1
XINVX1_456 INVX1_456/A gnd INVX1_456/Y vdd INVX1
XINVX1_445 INVX1_445/A gnd INVX1_445/Y vdd INVX1
XFILL_33_8_0 gnd vdd FILL
XAOI21X1_416 BUFX4_348/Y INVX1_379/Y OAI21X1_957/Y gnd OAI21X1_959/A vdd AOI21X1
XAOI21X1_405 BUFX4_104/Y INVX1_361/Y BUFX4_361/Y gnd AOI21X1_405/Y vdd AOI21X1
XAOI21X1_438 BUFX4_103/Y AOI21X1_438/B AOI21X1_437/Y gnd AOI21X1_438/Y vdd AOI21X1
XAOI21X1_427 NAND2X1_13/A BUFX4_234/Y AOI21X1_427/C gnd AOI21X1_427/Y vdd AOI21X1
XAOI21X1_449 AOI21X1_449/A BUFX4_222/Y AOI21X1_449/C gnd NOR2X1_508/A vdd AOI21X1
XFILL_24_8_0 gnd vdd FILL
XFILL_7_9_0 gnd vdd FILL
XMUX2X1_27 INVX1_35/Y MUX2X1_27/B MUX2X1_29/S gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_16 INVX1_21/Y MUX2X1_4/B MUX2X1_14/S gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_38 BUFX4_372/Y INVX1_46/Y NOR2X1_70/Y gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A INVX1_59/Y MUX2X1_50/S gnd MUX2X1_49/Y vdd MUX2X1
XFILL_15_8_0 gnd vdd FILL
XDFFPOSX1_519 INVX1_267/A CLKBUF1_97/Y MUX2X1_385/Y gnd vdd DFFPOSX1
XDFFPOSX1_508 NOR2X1_720/A CLKBUF1_60/Y AOI21X1_608/Y gnd vdd DFFPOSX1
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_275 INVX1_275/A gnd INVX1_275/Y vdd INVX1
XINVX1_264 INVX1_264/A gnd INVX1_264/Y vdd INVX1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XNAND2X1_20 traffic_Street_0[3] AOI21X1_7/B gnd OAI21X1_18/C vdd NAND2X1
XNAND2X1_31 INVX8_12/A INVX4_4/Y gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_42 INVX8_17/A INVX8_9/A gnd MUX2X1_66/S vdd NAND2X1
XNAND2X1_53 INVX8_19/A INVX4_4/Y gnd NAND2X1_53/Y vdd NAND2X1
XNAND2X1_86 AND2X2_24/B NAND2X1_2/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_75 INVX8_25/A INVX4_2/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_64 INVX8_22/A INVX4_3/Y gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_97 NAND2X1_97/A OAI21X1_7/B gnd NAND2X1_97/Y vdd NAND2X1
XNOR2X1_600 address[6] OAI22X1_81/Y gnd OAI22X1_94/A vdd NOR2X1
XFILL_42_1 gnd vdd FILL
XNOR2X1_633 NOR2X1_633/A NOR2X1_65/Y gnd NOR2X1_633/Y vdd NOR2X1
XNOR2X1_644 NOR2X1_644/A MUX2X1_50/S gnd NOR2X1_644/Y vdd NOR2X1
XNOR2X1_611 NOR2X1_611/A BUFX4_364/Y gnd OAI22X1_85/A vdd NOR2X1
XNOR2X1_622 NOR2X1_231/A BUFX4_366/Y gnd OAI22X1_92/A vdd NOR2X1
XNOR2X1_666 NOR2X1_666/A AOI21X1_72/B gnd NOR2X1_666/Y vdd NOR2X1
XNOR2X1_677 NOR2X1_677/A MUX2X1_92/S gnd NOR2X1_677/Y vdd NOR2X1
XNOR2X1_655 NOR2X1_655/A NOR2X1_107/B gnd NOR2X1_655/Y vdd NOR2X1
XNOR2X1_699 AND2X2_29/B INVX1_219/A gnd NOR2X1_699/Y vdd NOR2X1
XNOR2X1_688 MUX2X1_232/A MUX2X1_340/S gnd NOR2X1_688/Y vdd NOR2X1
XAOI21X1_213 INVX2_16/Y AND2X2_2/A AOI21X1_213/C gnd OR2X2_5/A vdd AOI21X1
XAOI21X1_202 BUFX4_174/Y MUX2X1_57/A AND2X2_3/B gnd AOI21X1_212/B vdd AOI21X1
XAOI21X1_224 AOI21X1_224/A OAI21X1_477/Y AND2X2_8/Y gnd AOI21X1_224/Y vdd AOI21X1
XAOI21X1_235 XOR2X1_3/A NAND3X1_46/B NAND3X1_47/Y gnd AOI21X1_235/Y vdd AOI21X1
XAOI21X1_257 BUFX4_149/Y OAI21X1_567/Y AOI21X1_257/C gnd MUX2X1_178/A vdd AOI21X1
XAOI21X1_246 AOI22X1_10/Y AOI21X1_246/B AOI21X1_246/C gnd OAI22X1_3/C vdd AOI21X1
XAOI21X1_268 BUFX4_356/Y INVX1_246/Y AOI21X1_268/C gnd AOI21X1_268/Y vdd AOI21X1
XAOI21X1_279 AOI21X1_279/A OAI21X1_604/Y BUFX4_207/Y gnd AOI21X1_280/C vdd AOI21X1
XOAI21X1_1441 BUFX4_420/Y NAND2X1_68/Y OAI21X1_1440/Y gnd OAI21X1_1441/Y vdd OAI21X1
XOAI21X1_1430 BUFX4_123/Y BUFX4_141/Y INVX1_237/A gnd OAI21X1_1431/C vdd OAI21X1
XOAI21X1_1463 BUFX4_126/Y BUFX4_433/Y OAI21X1_1157/B gnd OAI21X1_1463/Y vdd OAI21X1
XOAI21X1_1452 BUFX4_384/Y BUFX4_433/Y OAI21X1_1452/C gnd OAI21X1_1453/C vdd OAI21X1
XOAI21X1_1474 BUFX4_445/Y NAND2X1_73/Y OAI21X1_1473/Y gnd OAI21X1_1474/Y vdd OAI21X1
XOAI21X1_1496 NAND2X1_75/Y BUFX4_318/Y OAI21X1_1496/C gnd DFFPOSX1_498/D vdd OAI21X1
XOAI21X1_1485 BUFX4_188/Y BUFX4_161/Y AND2X2_41/B gnd OAI21X1_1486/C vdd OAI21X1
XDFFPOSX1_1026 OAI21X1_310/C CLKBUF1_2/Y OAI21X1_311/Y gnd vdd DFFPOSX1
XDFFPOSX1_1004 NOR2X1_459/A CLKBUF1_60/Y OAI21X1_291/Y gnd vdd DFFPOSX1
XDFFPOSX1_1015 NOR2X1_384/A CLKBUF1_67/Y AOI21X1_144/Y gnd vdd DFFPOSX1
XDFFPOSX1_1037 INVX1_407/A CLKBUF1_64/Y OAI21X1_317/Y gnd vdd DFFPOSX1
XDFFPOSX1_1048 NOR2X1_247/A CLKBUF1_67/Y AOI21X1_157/Y gnd vdd DFFPOSX1
XOAI22X1_2 OAI22X1_2/A OAI22X1_2/B OAI22X1_2/C OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XFILL_47_7_0 gnd vdd FILL
XFILL_30_6_0 gnd vdd FILL
XDFFPOSX1_305 NOR2X1_669/A CLKBUF1_2/Y AOI21X1_557/Y gnd vdd DFFPOSX1
XDFFPOSX1_338 NOR2X1_655/A CLKBUF1_88/Y AOI21X1_543/Y gnd vdd DFFPOSX1
XDFFPOSX1_316 INVX1_349/A CLKBUF1_48/Y MUX2X1_286/Y gnd vdd DFFPOSX1
XDFFPOSX1_327 NOR2X1_422/B CLKBUF1_75/Y AOI21X1_550/Y gnd vdd DFFPOSX1
XDFFPOSX1_349 NOR2X1_654/A CLKBUF1_58/Y AOI21X1_542/Y gnd vdd DFFPOSX1
XFILL_38_7_0 gnd vdd FILL
XBUFX4_370 BUFX4_25/Y gnd BUFX4_370/Y vdd BUFX4
XBUFX4_381 INVX8_14/Y gnd BUFX4_381/Y vdd BUFX4
XNOR2X1_452 NOR2X1_452/A BUFX4_346/Y gnd NOR2X1_452/Y vdd NOR2X1
XBUFX4_392 INVX8_28/Y gnd BUFX4_392/Y vdd BUFX4
XNOR2X1_441 OAI21X1_61/C BUFX4_364/Y gnd OAI22X1_23/A vdd NOR2X1
XNOR2X1_430 BUFX4_416/Y NOR2X1_430/B gnd NOR2X1_430/Y vdd NOR2X1
XNOR2X1_474 BUFX4_103/Y NOR2X1_474/B gnd NOR2X1_475/A vdd NOR2X1
XNOR2X1_485 INVX8_32/A NOR2X1_485/B gnd NOR2X1_485/Y vdd NOR2X1
XNOR2X1_463 BUFX4_419/Y NOR2X1_463/B gnd OAI22X1_36/B vdd NOR2X1
XNOR2X1_496 BUFX4_417/Y NOR2X1_496/B gnd NOR2X1_496/Y vdd NOR2X1
XOAI21X1_925 INVX1_355/Y BUFX4_262/Y NAND2X1_278/Y gnd OAI21X1_925/Y vdd OAI21X1
XFILL_21_6_0 gnd vdd FILL
XOAI21X1_914 INVX1_345/Y BUFX4_252/Y OAI21X1_914/C gnd MUX2X1_229/A vdd OAI21X1
XOAI21X1_903 NOR2X1_211/A BUFX4_242/Y BUFX4_83/Y gnd OAI22X1_34/B vdd OAI21X1
XOAI21X1_947 BUFX4_271/Y OAI21X1_947/B BUFX4_110/Y gnd AOI21X1_411/C vdd OAI21X1
XOAI21X1_936 BUFX4_35/Y INVX1_363/Y BUFX4_266/Y gnd OAI21X1_936/Y vdd OAI21X1
XOAI21X1_958 BUFX4_282/Y OAI21X1_958/B BUFX4_116/Y gnd AOI21X1_417/C vdd OAI21X1
XOAI21X1_969 INVX1_387/Y BUFX4_223/Y NAND2X1_291/Y gnd MUX2X1_238/B vdd OAI21X1
XMUX2X1_403 BUFX4_324/Y INVX1_424/Y NOR2X1_261/B gnd MUX2X1_403/Y vdd MUX2X1
XDFFPOSX1_850 NOR2X1_134/A CLKBUF1_62/Y AOI21X1_78/Y gnd vdd DFFPOSX1
XOAI21X1_1282 NAND2X1_32/Y BUFX4_442/Y OAI21X1_1282/C gnd DFFPOSX1_142/D vdd OAI21X1
XOAI21X1_1271 BUFX4_301/Y BUFX4_44/Y OAI21X1_1087/B gnd OAI21X1_1272/C vdd OAI21X1
XOAI21X1_1260 INVX1_445/Y BUFX4_259/Y BUFX4_155/Y gnd OAI21X1_1260/Y vdd OAI21X1
XDFFPOSX1_872 INVX1_107/A CLKBUF1_5/Y MUX2X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_861 INVX1_104/A CLKBUF1_93/Y MUX2X1_91/Y gnd vdd DFFPOSX1
XOAI21X1_1293 NAND2X1_36/Y BUFX4_424/Y OAI21X1_1293/C gnd DFFPOSX1_231/D vdd OAI21X1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XDFFPOSX1_883 INVX1_287/A CLKBUF1_86/Y OAI21X1_193/Y gnd vdd DFFPOSX1
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XDFFPOSX1_894 NOR2X1_588/A CLKBUF1_8/Y OAI21X1_215/Y gnd vdd DFFPOSX1
XFILL_4_7_0 gnd vdd FILL
XFILL_29_7_0 gnd vdd FILL
XOAI21X1_18 INVX1_32/Y AOI21X1_7/B OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 BUFX4_125/Y BUFX4_295/Y INVX1_331/A gnd OAI21X1_30/C vdd OAI21X1
XFILL_12_6_0 gnd vdd FILL
XDFFPOSX1_102 NOR2X1_286/A CLKBUF1_103/Y AOI21X1_189/Y gnd vdd DFFPOSX1
XDFFPOSX1_146 INVX1_223/A CLKBUF1_80/Y OAI21X1_1274/Y gnd vdd DFFPOSX1
XDFFPOSX1_135 NAND2X1_261/A CLKBUF1_6/Y OAI21X1_432/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 INVX1_401/A CLKBUF1_100/Y OAI21X1_426/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 OAI21X1_419/C CLKBUF1_88/Y OAI21X1_420/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 NOR2X1_689/A CLKBUF1_45/Y AOI21X1_577/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 NOR2X1_680/A CLKBUF1_26/Y AOI21X1_568/Y gnd vdd DFFPOSX1
XDFFPOSX1_179 INVX1_446/A CLKBUF1_89/Y MUX2X1_276/Y gnd vdd DFFPOSX1
XNAND2X1_205 NOR2X1_294/A BUFX4_248/Y gnd OAI21X1_650/C vdd NAND2X1
XNAND2X1_216 NOR2X1_159/A BUFX4_285/Y gnd NAND2X1_216/Y vdd NAND2X1
XNAND2X1_238 NAND2X1_238/A BUFX4_348/Y gnd NAND2X1_238/Y vdd NAND2X1
XNAND2X1_227 enable INVX1_2/Y gnd NOR2X1_624/A vdd NAND2X1
XNAND2X1_249 OAI21X1_111/C BUFX4_255/Y gnd NAND2X1_249/Y vdd NAND2X1
XNOR2X1_260 BUFX4_198/Y BUFX4_57/Y gnd NOR2X1_261/B vdd NOR2X1
XNOR2X1_293 NOR2X1_293/A NOR2X1_43/B gnd NOR2X1_293/Y vdd NOR2X1
XNOR2X1_282 NOR2X1_282/A NOR2X1_30/B gnd NOR2X1_282/Y vdd NOR2X1
XNOR2X1_271 NOR2X1_271/A MUX2X1_410/S gnd NOR2X1_271/Y vdd NOR2X1
XOAI21X1_722 INVX2_2/Y read_Write BUFX2_5/A gnd OAI21X1_723/C vdd OAI21X1
XOAI21X1_700 NOR2X1_58/A BUFX4_227/Y BUFX4_92/Y gnd OAI22X1_16/B vdd OAI21X1
XOAI21X1_733 OAI21X1_733/A AND2X2_27/Y OAI21X1_733/C gnd OAI21X1_733/Y vdd OAI21X1
XOAI21X1_711 INVX1_65/Y AND2X2_22/A OAI21X1_711/C gnd MUX2X1_206/A vdd OAI21X1
XOAI21X1_766 BUFX4_354/Y OAI21X1_766/B BUFX4_150/Y gnd OAI21X1_768/B vdd OAI21X1
XOAI21X1_744 OAI21X1_743/Y NOR2X1_420/Y BUFX4_41/Y gnd OAI21X1_744/Y vdd OAI21X1
XOAI21X1_755 BUFX4_367/Y NOR2X1_684/A BUFX4_148/Y gnd OAI21X1_757/B vdd OAI21X1
XOAI21X1_788 INVX1_323/Y BUFX4_233/Y BUFX4_84/Y gnd OAI21X1_788/Y vdd OAI21X1
XOAI21X1_799 BUFX4_360/Y INVX1_19/A BUFX4_149/Y gnd AOI21X1_351/C vdd OAI21X1
XOAI21X1_777 INVX8_31/A NOR2X1_712/A BUFX4_77/Y gnd OAI22X1_22/B vdd OAI21X1
XMUX2X1_211 MUX2X1_211/A MUX2X1_211/B INVX8_32/A gnd MUX2X1_213/A vdd MUX2X1
XMUX2X1_200 MUX2X1_200/A MUX2X1_200/B BUFX4_86/Y gnd MUX2X1_200/Y vdd MUX2X1
XMUX2X1_222 MUX2X1_222/A MUX2X1_221/Y BUFX4_165/Y gnd MUX2X1_222/Y vdd MUX2X1
XOAI21X1_1090 BUFX4_334/Y NOR2X1_635/A BUFX4_157/Y gnd OAI22X1_49/C vdd OAI21X1
XMUX2X1_233 MUX2X1_233/A MUX2X1_233/B BUFX4_111/Y gnd MUX2X1_233/Y vdd MUX2X1
XMUX2X1_244 MUX2X1_244/A MUX2X1_244/B BUFX4_100/Y gnd MUX2X1_244/Y vdd MUX2X1
XMUX2X1_255 MUX2X1_255/A OAI22X1_46/Y INVX8_33/Y gnd MUX2X1_255/Y vdd MUX2X1
XMUX2X1_299 INVX1_368/Y BUFX4_68/Y MUX2X1_59/S gnd MUX2X1_299/Y vdd MUX2X1
XMUX2X1_266 MUX2X1_266/A MUX2X1_266/B BUFX4_111/Y gnd MUX2X1_266/Y vdd MUX2X1
XDFFPOSX1_691 NOR2X1_58/A CLKBUF1_94/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XMUX2X1_288 BUFX4_440/Y INVX1_226/Y MUX2X1_50/S gnd MUX2X1_288/Y vdd MUX2X1
XDFFPOSX1_680 NOR2X1_50/A CLKBUF1_87/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XMUX2X1_277 INVX1_346/Y BUFX4_63/Y MUX2X1_42/S gnd MUX2X1_277/Y vdd MUX2X1
XFILL_44_5_0 gnd vdd FILL
XCLKBUF1_19 BUFX4_1/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_51 address[4] gnd BUFX4_51/Y vdd BUFX4
XBUFX4_40 BUFX4_33/A gnd BUFX4_40/Y vdd BUFX4
XBUFX4_62 INVX8_6/Y gnd BUFX4_62/Y vdd BUFX4
XBUFX4_95 BUFX4_14/Y gnd BUFX4_95/Y vdd BUFX4
XBUFX4_84 BUFX4_87/A gnd BUFX4_84/Y vdd BUFX4
XBUFX4_73 INVX8_4/Y gnd BUFX4_73/Y vdd BUFX4
XFILL_35_5_0 gnd vdd FILL
XOR2X2_3 traffic_Street_0[1] traffic_Street_0[2] gnd OR2X2_3/Y vdd OR2X2
XXNOR2X1_5 AOI22X1_7/C XNOR2X1_5/B gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XINVX8_10 INVX8_10/A gnd INVX8_10/Y vdd INVX8
XINVX8_21 INVX8_21/A gnd INVX8_21/Y vdd INVX8
XINVX8_32 INVX8_32/A gnd INVX8_32/Y vdd INVX8
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOAI21X1_530 OAI21X1_515/Y INVX4_9/A INVX1_211/A gnd AND2X2_14/A vdd OAI21X1
XOAI21X1_541 BUFX4_307/Y INVX4_11/Y NOR2X1_352/A gnd OAI21X1_541/Y vdd OAI21X1
XFILL_10_9_1 gnd vdd FILL
XOAI21X1_574 OAI21X1_573/Y NOR2X1_368/Y BUFX4_35/Y gnd OAI22X1_4/A vdd OAI21X1
XOAI21X1_563 INVX1_227/Y BUFX4_230/Y OAI21X1_563/C gnd MUX2X1_177/B vdd OAI21X1
XOAI21X1_552 BUFX4_220/Y NOR2X1_637/A AOI21X1_247/Y gnd NAND3X1_71/B vdd OAI21X1
XOAI21X1_596 BUFX4_341/Y INVX1_254/Y OAI21X1_596/C gnd OAI21X1_598/C vdd OAI21X1
XOAI21X1_585 INVX1_245/Y BUFX4_251/Y BUFX4_150/Y gnd OAI21X1_585/Y vdd OAI21X1
.ends

