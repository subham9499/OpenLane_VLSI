magic
tech scmos
timestamp 1607101874
<< metal1 >>
rect 848 5103 850 5107
rect 854 5103 857 5107
rect 861 5103 864 5107
rect 1872 5103 1874 5107
rect 1878 5103 1881 5107
rect 1885 5103 1888 5107
rect 2888 5103 2890 5107
rect 2894 5103 2897 5107
rect 2901 5103 2904 5107
rect 3920 5103 3922 5107
rect 3926 5103 3929 5107
rect 3933 5103 3936 5107
rect 4936 5103 4938 5107
rect 4942 5103 4945 5107
rect 4949 5103 4952 5107
rect 3398 5088 3409 5091
rect 634 5078 641 5081
rect 1086 5078 1102 5081
rect 2462 5078 2470 5081
rect 2502 5078 2521 5081
rect 3406 5081 3409 5088
rect 2718 5078 2729 5081
rect 2734 5078 2753 5081
rect 2870 5078 2881 5081
rect 3406 5078 3425 5081
rect 3526 5078 3537 5081
rect 3570 5078 3571 5082
rect 3830 5078 3841 5081
rect 4342 5078 4353 5081
rect 1726 5076 1730 5078
rect 2718 5077 2722 5078
rect 2870 5077 2874 5078
rect 3526 5077 3530 5078
rect 3830 5077 3834 5078
rect 4342 5077 4346 5078
rect 94 5071 98 5074
rect 94 5068 105 5071
rect 270 5071 274 5074
rect 270 5068 281 5071
rect 318 5068 326 5071
rect 858 5068 865 5071
rect 886 5068 894 5071
rect 1110 5068 1121 5071
rect 1234 5068 1241 5071
rect 1250 5068 1257 5071
rect 1326 5068 1342 5071
rect 1586 5068 1601 5071
rect 2418 5068 2433 5071
rect 2470 5068 2486 5071
rect 2494 5068 2502 5071
rect 2754 5068 2761 5071
rect 2898 5068 2921 5071
rect 3118 5068 3129 5071
rect 3302 5068 3314 5071
rect 3958 5068 3966 5071
rect 38 5058 46 5061
rect 118 5061 121 5068
rect 118 5058 129 5061
rect 166 5058 174 5061
rect 286 5058 305 5061
rect 354 5058 369 5061
rect 414 5058 425 5061
rect 718 5058 726 5061
rect 754 5058 761 5061
rect 786 5058 793 5061
rect 882 5058 905 5061
rect 966 5058 978 5061
rect 1118 5062 1121 5068
rect 1246 5058 1254 5061
rect 1282 5058 1297 5061
rect 1438 5058 1449 5061
rect 1958 5058 1966 5061
rect 2470 5058 2473 5068
rect 2886 5058 2918 5061
rect 3118 5061 3121 5068
rect 3078 5058 3097 5061
rect 3102 5058 3121 5061
rect 3266 5058 3273 5061
rect 3538 5058 3545 5061
rect 5114 5058 5121 5061
rect 5254 5058 5265 5061
rect 302 5048 305 5058
rect 974 5057 978 5058
rect 1438 5057 1442 5058
rect 334 5048 361 5051
rect 762 5048 766 5052
rect 774 5048 782 5051
rect 842 5048 862 5051
rect 3078 5048 3081 5058
rect 3174 5048 3177 5058
rect 3838 5051 3841 5058
rect 3838 5048 3849 5051
rect 5254 5048 5257 5058
rect 106 5038 113 5041
rect 606 5041 610 5044
rect 594 5038 610 5041
rect 2187 5038 2190 5042
rect 3426 5038 3433 5041
rect 5278 5038 5302 5041
rect 4454 5028 4470 5031
rect 4474 5018 4481 5021
rect 4994 5018 4995 5022
rect 5045 5018 5046 5022
rect 5242 5018 5243 5022
rect 328 5003 330 5007
rect 334 5003 337 5007
rect 341 5003 344 5007
rect 1352 5003 1354 5007
rect 1358 5003 1361 5007
rect 1365 5003 1368 5007
rect 2384 5003 2386 5007
rect 2390 5003 2393 5007
rect 2397 5003 2400 5007
rect 3400 5003 3402 5007
rect 3406 5003 3409 5007
rect 3413 5003 3416 5007
rect 4424 5003 4426 5007
rect 4430 5003 4433 5007
rect 4437 5003 4440 5007
rect 501 4988 502 4992
rect 666 4988 668 4992
rect 1941 4988 1942 4992
rect 3634 4988 3635 4992
rect 533 4968 534 4972
rect 834 4968 835 4972
rect 882 4968 883 4972
rect 2043 4968 2046 4972
rect 3227 4968 3230 4972
rect 3450 4968 3453 4972
rect 3541 4968 3542 4972
rect 3850 4968 3853 4972
rect 258 4958 265 4961
rect 626 4958 630 4962
rect 986 4958 993 4961
rect 138 4948 145 4951
rect 698 4948 713 4951
rect 782 4948 790 4951
rect 806 4948 825 4951
rect 850 4948 881 4951
rect 990 4948 1001 4951
rect 1030 4948 1046 4951
rect 1062 4951 1065 4958
rect 1054 4948 1065 4951
rect 822 4942 825 4948
rect 990 4942 993 4948
rect 1206 4948 1217 4951
rect 1238 4951 1242 4954
rect 1334 4952 1338 4954
rect 1238 4948 1257 4951
rect 1262 4948 1278 4951
rect 1398 4948 1410 4951
rect 1514 4948 1521 4951
rect 1678 4951 1682 4953
rect 1670 4948 1682 4951
rect 1926 4951 1929 4961
rect 2074 4958 2081 4961
rect 2214 4958 2222 4961
rect 1910 4948 1929 4951
rect 1406 4946 1410 4948
rect 2394 4948 2401 4951
rect 2490 4948 2497 4951
rect 2950 4948 2958 4951
rect 3006 4951 3009 4958
rect 2998 4948 3009 4951
rect 3142 4948 3150 4951
rect 3278 4951 3281 4961
rect 3666 4958 3670 4962
rect 3278 4948 3297 4951
rect 3562 4948 3569 4951
rect 4166 4951 4169 4961
rect 4498 4958 4502 4962
rect 5038 4952 5041 4961
rect 4150 4948 4169 4951
rect 4482 4948 4497 4951
rect 4594 4948 4601 4951
rect 4630 4948 4649 4951
rect 326 4938 350 4941
rect 390 4938 398 4941
rect 554 4938 561 4941
rect 762 4938 769 4941
rect 786 4938 793 4941
rect 1010 4938 1017 4941
rect 1062 4938 1074 4941
rect 1170 4938 1177 4941
rect 1220 4938 1222 4942
rect 1294 4938 1305 4941
rect 1390 4938 1401 4941
rect 1766 4938 1778 4941
rect 1954 4938 1969 4941
rect 2598 4938 2609 4941
rect 2886 4938 2921 4941
rect 2982 4938 3001 4941
rect 3606 4938 3614 4941
rect 3869 4938 3870 4942
rect 3918 4938 3946 4941
rect 4482 4938 4489 4941
rect 4630 4938 4638 4941
rect 4646 4938 4654 4941
rect 1070 4936 1074 4938
rect 1398 4932 1401 4938
rect 346 4928 353 4931
rect 390 4928 401 4931
rect 2189 4928 2190 4932
rect 2350 4928 2369 4931
rect 2374 4928 2390 4931
rect 2438 4928 2457 4931
rect 2486 4928 2489 4938
rect 2598 4932 2601 4938
rect 2886 4928 2889 4938
rect 2898 4928 2910 4931
rect 3014 4931 3018 4933
rect 3230 4932 3234 4936
rect 3006 4928 3018 4931
rect 3130 4928 3131 4932
rect 4662 4931 4666 4933
rect 4654 4928 4666 4931
rect 4766 4928 4785 4931
rect 5062 4931 5066 4936
rect 5062 4928 5078 4931
rect 470 4921 473 4928
rect 470 4918 481 4921
rect 1882 4918 1889 4921
rect 3418 4918 3433 4921
rect 848 4903 850 4907
rect 854 4903 857 4907
rect 861 4903 864 4907
rect 1872 4903 1874 4907
rect 1878 4903 1881 4907
rect 1885 4903 1888 4907
rect 2888 4903 2890 4907
rect 2894 4903 2897 4907
rect 2901 4903 2904 4907
rect 3920 4903 3922 4907
rect 3926 4903 3929 4907
rect 3933 4903 3936 4907
rect 4936 4903 4938 4907
rect 4942 4903 4945 4907
rect 4949 4903 4952 4907
rect 533 4888 534 4892
rect 1866 4888 1867 4892
rect 2382 4888 2393 4891
rect 4205 4888 4206 4892
rect 4934 4888 4945 4891
rect 106 4878 113 4881
rect 682 4878 689 4881
rect 902 4878 913 4881
rect 198 4868 217 4871
rect 238 4868 246 4871
rect 382 4868 390 4871
rect 578 4868 585 4871
rect 642 4868 649 4871
rect 670 4868 689 4871
rect 738 4868 753 4871
rect 838 4868 854 4871
rect 878 4868 897 4871
rect 966 4871 969 4881
rect 1518 4878 1530 4881
rect 1822 4878 1833 4881
rect 2006 4878 2025 4881
rect 2126 4878 2137 4881
rect 2170 4878 2171 4882
rect 2390 4881 2393 4888
rect 2390 4878 2409 4881
rect 2646 4878 2654 4881
rect 2838 4878 2849 4881
rect 3294 4878 3313 4881
rect 4014 4878 4033 4881
rect 4118 4878 4126 4881
rect 4238 4878 4246 4881
rect 966 4868 974 4871
rect 1286 4871 1290 4874
rect 1278 4868 1290 4871
rect 1394 4868 1401 4871
rect 234 4858 257 4861
rect 346 4858 369 4861
rect 378 4858 401 4861
rect 586 4858 593 4861
rect 598 4858 617 4861
rect 666 4858 678 4861
rect 686 4861 689 4868
rect 878 4862 881 4868
rect 686 4858 702 4861
rect 830 4858 862 4861
rect 950 4861 953 4868
rect 1478 4871 1481 4878
rect 1526 4877 1530 4878
rect 1822 4877 1826 4878
rect 2126 4877 2130 4878
rect 2838 4877 2842 4878
rect 4286 4872 4289 4881
rect 4438 4878 4446 4881
rect 4550 4878 4561 4881
rect 4742 4878 4754 4881
rect 4942 4881 4945 4888
rect 4942 4878 4961 4881
rect 4550 4877 4554 4878
rect 4750 4877 4754 4878
rect 1478 4868 1489 4871
rect 1494 4868 1502 4871
rect 2586 4868 2593 4871
rect 2866 4868 2873 4871
rect 2942 4868 2958 4871
rect 3110 4868 3118 4871
rect 3382 4868 3398 4871
rect 3558 4868 3566 4871
rect 4578 4868 4585 4871
rect 4838 4868 4850 4871
rect 4978 4868 4985 4871
rect 950 4858 961 4861
rect 1038 4858 1057 4861
rect 1070 4858 1078 4861
rect 1262 4858 1273 4861
rect 1330 4858 1345 4861
rect 2574 4858 2593 4861
rect 2650 4858 2657 4861
rect 2854 4858 2873 4861
rect 2958 4858 2961 4868
rect 3046 4858 3065 4861
rect 3110 4858 3129 4861
rect 3342 4858 3361 4861
rect 3374 4858 3382 4861
rect 3518 4858 3537 4861
rect 3634 4858 3641 4861
rect 3702 4858 3721 4861
rect 3766 4858 3785 4861
rect 3942 4858 3961 4861
rect 4242 4858 4249 4861
rect 4566 4858 4585 4861
rect 4618 4858 4625 4861
rect 4654 4858 4673 4861
rect 4718 4858 4737 4861
rect 4794 4858 4809 4861
rect 4966 4858 4985 4861
rect 158 4848 166 4851
rect 302 4848 310 4851
rect 1054 4848 1057 4858
rect 1186 4848 1190 4852
rect 3046 4848 3049 4858
rect 3358 4848 3361 4858
rect 3534 4848 3537 4858
rect 3610 4848 3614 4852
rect 3674 4848 3678 4852
rect 3686 4848 3694 4851
rect 3718 4848 3721 4858
rect 3782 4848 3785 4858
rect 3958 4848 3961 4858
rect 258 4838 259 4842
rect 402 4838 403 4842
rect 138 4818 139 4822
rect 466 4818 467 4822
rect 874 4818 875 4822
rect 2637 4818 2638 4822
rect 3034 4818 3035 4822
rect 3373 4818 3374 4822
rect 3733 4818 3734 4822
rect 4058 4818 4059 4822
rect 4253 4818 4254 4822
rect 4429 4818 4430 4822
rect 5266 4818 5267 4822
rect 328 4803 330 4807
rect 334 4803 337 4807
rect 341 4803 344 4807
rect 1352 4803 1354 4807
rect 1358 4803 1361 4807
rect 1365 4803 1368 4807
rect 2384 4803 2386 4807
rect 2390 4803 2393 4807
rect 2397 4803 2400 4807
rect 3400 4803 3402 4807
rect 3406 4803 3409 4807
rect 3413 4803 3416 4807
rect 4424 4803 4426 4807
rect 4430 4803 4433 4807
rect 4437 4803 4440 4807
rect 114 4788 115 4792
rect 522 4788 523 4792
rect 773 4788 774 4792
rect 1501 4788 1502 4792
rect 802 4778 803 4782
rect 914 4768 915 4772
rect 2827 4768 2830 4772
rect 182 4758 190 4761
rect 678 4758 689 4761
rect 1338 4758 1345 4761
rect 3050 4758 3057 4761
rect 678 4752 682 4754
rect 174 4748 190 4751
rect 70 4738 78 4741
rect 230 4741 233 4748
rect 582 4748 590 4751
rect 726 4748 734 4751
rect 774 4748 798 4751
rect 818 4748 830 4751
rect 858 4748 873 4751
rect 986 4748 993 4751
rect 1062 4748 1078 4751
rect 1230 4748 1238 4751
rect 1310 4748 1329 4751
rect 222 4738 233 4741
rect 346 4738 353 4741
rect 486 4738 494 4741
rect 570 4738 577 4741
rect 582 4738 585 4748
rect 706 4738 713 4741
rect 782 4738 790 4741
rect 1358 4738 1366 4741
rect 1662 4741 1665 4751
rect 1718 4748 1737 4751
rect 2038 4748 2046 4751
rect 2270 4748 2278 4751
rect 2354 4748 2361 4751
rect 2574 4748 2593 4751
rect 2630 4742 2633 4751
rect 2854 4742 2857 4751
rect 2982 4748 2990 4751
rect 3710 4751 3713 4761
rect 3814 4753 3818 4758
rect 5190 4756 5194 4758
rect 3694 4748 3713 4751
rect 3918 4748 3942 4751
rect 4006 4742 4009 4751
rect 4106 4748 4113 4751
rect 4186 4748 4201 4751
rect 4526 4748 4545 4751
rect 4810 4748 4825 4751
rect 4894 4748 4910 4751
rect 5158 4742 5161 4751
rect 1650 4738 1665 4741
rect 1670 4738 1678 4741
rect 1718 4738 1726 4741
rect 1906 4738 1914 4741
rect 2174 4738 2193 4741
rect 2238 4738 2257 4741
rect 2750 4738 2762 4741
rect 3066 4738 3073 4741
rect 3926 4738 3950 4741
rect 4010 4738 4025 4741
rect 4054 4738 4073 4741
rect 4182 4738 4190 4741
rect 4718 4738 4737 4741
rect 4854 4738 4866 4741
rect 4990 4738 4998 4741
rect 5138 4738 5145 4741
rect 94 4728 105 4731
rect 486 4728 489 4738
rect 1342 4732 1345 4738
rect 566 4728 577 4731
rect 1342 4728 1350 4732
rect 1614 4728 1633 4731
rect 1750 4731 1754 4733
rect 1742 4728 1754 4731
rect 1766 4731 1770 4736
rect 1766 4728 1782 4731
rect 2190 4728 2193 4738
rect 2238 4728 2241 4738
rect 3470 4736 3474 4738
rect 2562 4728 2563 4732
rect 2662 4731 2666 4733
rect 2630 4728 2649 4731
rect 2654 4728 2666 4731
rect 2894 4728 2902 4731
rect 3038 4731 3042 4733
rect 3598 4732 3602 4736
rect 3038 4728 3049 4731
rect 3894 4728 3905 4731
rect 3974 4728 3985 4731
rect 4070 4728 4073 4738
rect 4206 4728 4214 4731
rect 4518 4728 4521 4738
rect 4734 4728 4737 4738
rect 5190 4731 5194 4733
rect 5158 4728 5177 4731
rect 5182 4728 5194 4731
rect 36 4718 38 4722
rect 846 4718 854 4721
rect 1018 4718 1020 4722
rect 1549 4718 1550 4722
rect 4950 4718 4966 4721
rect 848 4703 850 4707
rect 854 4703 857 4707
rect 861 4703 864 4707
rect 1872 4703 1874 4707
rect 1878 4703 1881 4707
rect 1885 4703 1888 4707
rect 2888 4703 2890 4707
rect 2894 4703 2897 4707
rect 2901 4703 2904 4707
rect 3920 4703 3922 4707
rect 3926 4703 3929 4707
rect 3933 4703 3936 4707
rect 4936 4703 4938 4707
rect 4942 4703 4945 4707
rect 4949 4703 4952 4707
rect 226 4688 227 4692
rect 668 4688 670 4692
rect 690 4688 697 4691
rect 1350 4688 1358 4691
rect 2026 4688 2027 4692
rect 3918 4688 3929 4691
rect 4914 4688 4929 4691
rect 102 4662 105 4671
rect 198 4671 201 4681
rect 190 4668 201 4671
rect 254 4668 265 4671
rect 366 4668 369 4678
rect 430 4671 433 4681
rect 462 4678 478 4681
rect 414 4668 433 4671
rect 726 4668 742 4671
rect 898 4668 913 4671
rect 970 4668 977 4671
rect 1150 4668 1169 4671
rect 1250 4668 1257 4671
rect 1318 4671 1321 4678
rect 1334 4671 1337 4681
rect 1370 4678 1377 4681
rect 1630 4678 1641 4681
rect 1774 4678 1793 4681
rect 1630 4677 1634 4678
rect 1318 4668 1329 4671
rect 1334 4668 1353 4671
rect 1390 4668 1398 4671
rect 1994 4668 2001 4671
rect 2302 4671 2305 4681
rect 2442 4678 2449 4681
rect 2466 4678 2473 4681
rect 2510 4678 2529 4681
rect 2534 4678 2542 4681
rect 2302 4668 2321 4671
rect 2566 4671 2569 4681
rect 2658 4678 2674 4681
rect 2670 4674 2674 4678
rect 2782 4678 2793 4681
rect 3046 4678 3057 4681
rect 3158 4678 3177 4681
rect 3762 4678 3763 4682
rect 3802 4678 3809 4681
rect 3926 4681 3929 4688
rect 3926 4678 3945 4681
rect 4030 4678 4049 4681
rect 4058 4678 4066 4681
rect 2782 4677 2786 4678
rect 3046 4677 3050 4678
rect 4062 4677 4066 4678
rect 2550 4668 2569 4671
rect 2878 4668 2913 4671
rect 3074 4668 3081 4671
rect 3134 4668 3142 4671
rect 3426 4668 3433 4671
rect 3542 4668 3561 4671
rect 3962 4668 3969 4671
rect 4374 4671 4377 4681
rect 4246 4668 4258 4671
rect 4358 4668 4377 4671
rect 4518 4671 4521 4678
rect 4510 4668 4521 4671
rect 4694 4671 4697 4681
rect 4862 4678 4881 4681
rect 4678 4668 4697 4671
rect 5078 4671 5081 4681
rect 5078 4668 5097 4671
rect 5106 4668 5121 4671
rect 198 4662 201 4668
rect 38 4658 46 4661
rect 118 4658 145 4661
rect 222 4658 241 4661
rect 446 4658 457 4661
rect 726 4658 729 4668
rect 782 4658 809 4661
rect 834 4658 841 4661
rect 902 4658 918 4661
rect 1094 4658 1102 4661
rect 1114 4658 1121 4661
rect 1774 4658 1777 4668
rect 2126 4658 2145 4661
rect 2538 4658 2545 4661
rect 2798 4658 2806 4661
rect 2810 4658 2817 4661
rect 3062 4658 3081 4661
rect 3294 4658 3313 4661
rect 3526 4658 3545 4661
rect 3582 4658 3601 4661
rect 3774 4658 3793 4661
rect 3950 4658 3969 4661
rect 4114 4658 4121 4661
rect 4398 4658 4406 4661
rect 4642 4658 4649 4661
rect 4758 4658 4766 4661
rect 5154 4658 5161 4661
rect 5250 4658 5265 4661
rect 214 4651 217 4658
rect 166 4648 177 4651
rect 206 4648 217 4651
rect 238 4648 241 4658
rect 1102 4648 1113 4651
rect 1210 4648 1217 4651
rect 3582 4648 3585 4658
rect 4614 4652 4618 4657
rect 1102 4642 1105 4648
rect 618 4638 633 4641
rect 842 4638 843 4642
rect 1875 4638 1878 4642
rect 1414 4628 1417 4638
rect 1229 4618 1230 4622
rect 1301 4618 1302 4622
rect 3221 4618 3222 4622
rect 3442 4618 3443 4622
rect 3474 4618 3475 4622
rect 3570 4618 3571 4622
rect 3918 4618 3934 4621
rect 4650 4618 4651 4622
rect 5037 4618 5038 4622
rect 328 4603 330 4607
rect 334 4603 337 4607
rect 341 4603 344 4607
rect 1352 4603 1354 4607
rect 1358 4603 1361 4607
rect 1365 4603 1368 4607
rect 2384 4603 2386 4607
rect 2390 4603 2393 4607
rect 2397 4603 2400 4607
rect 3400 4603 3402 4607
rect 3406 4603 3409 4607
rect 3413 4603 3416 4607
rect 4424 4603 4426 4607
rect 4430 4603 4433 4607
rect 4437 4603 4440 4607
rect 906 4588 907 4592
rect 1282 4588 1283 4592
rect 2522 4588 2523 4592
rect 4221 4588 4222 4592
rect 5141 4588 5142 4592
rect 1118 4572 1121 4581
rect 125 4568 126 4572
rect 154 4568 155 4572
rect 250 4568 251 4572
rect 594 4568 614 4571
rect 1230 4568 1241 4571
rect 3611 4568 3614 4572
rect 1238 4562 1241 4568
rect 202 4558 209 4561
rect 130 4548 153 4551
rect 286 4548 294 4551
rect 630 4551 633 4561
rect 740 4558 742 4562
rect 1434 4558 1441 4561
rect 2382 4558 2390 4561
rect 2870 4558 2878 4561
rect 630 4548 638 4551
rect 818 4548 841 4551
rect 1014 4548 1030 4551
rect 1186 4548 1201 4551
rect 1378 4548 1385 4551
rect 1442 4548 1449 4551
rect 1614 4551 1617 4558
rect 1614 4548 1625 4551
rect 1814 4551 1818 4553
rect 1798 4548 1818 4551
rect 1866 4548 1873 4551
rect 2458 4548 2465 4551
rect 2690 4548 2705 4551
rect 3262 4548 3270 4551
rect 3302 4551 3305 4561
rect 3314 4558 3318 4562
rect 3826 4558 3830 4562
rect 4066 4558 4070 4562
rect 3286 4548 3305 4551
rect 3450 4548 3457 4551
rect 3494 4548 3521 4551
rect 3646 4548 3657 4551
rect 3862 4548 3870 4551
rect 3654 4542 3657 4548
rect 4058 4548 4065 4551
rect 4254 4548 4262 4551
rect 4278 4548 4286 4551
rect 4554 4548 4569 4551
rect 4710 4548 4718 4551
rect 4846 4548 4854 4551
rect 5058 4548 5065 4551
rect 5258 4548 5273 4551
rect 34 4538 41 4541
rect 134 4538 142 4541
rect 442 4538 457 4541
rect 474 4538 481 4541
rect 486 4538 497 4541
rect 654 4538 673 4541
rect 774 4538 793 4541
rect 810 4538 830 4541
rect 866 4538 897 4541
rect 946 4538 958 4541
rect 1238 4538 1246 4541
rect 1254 4538 1273 4541
rect 1398 4538 1425 4541
rect 1902 4538 1910 4541
rect 2070 4538 2082 4541
rect 2214 4538 2222 4541
rect 2330 4538 2337 4541
rect 2810 4538 2825 4541
rect 3238 4538 3257 4541
rect 3266 4538 3273 4541
rect 3930 4538 3945 4541
rect 4462 4538 4481 4541
rect 4662 4538 4681 4541
rect 4750 4538 4758 4541
rect 5034 4538 5041 4541
rect 5150 4538 5158 4541
rect 654 4528 657 4538
rect 790 4528 793 4538
rect 1030 4528 1054 4531
rect 1606 4531 1610 4533
rect 1606 4528 1617 4531
rect 1950 4528 1969 4531
rect 1982 4531 1986 4533
rect 1978 4528 1986 4531
rect 2166 4531 2170 4533
rect 2166 4528 2174 4531
rect 2182 4528 2201 4531
rect 2838 4528 2857 4531
rect 2878 4528 2897 4531
rect 3238 4528 3241 4538
rect 3630 4531 3634 4533
rect 3630 4528 3641 4531
rect 3738 4528 3745 4531
rect 3754 4528 3761 4531
rect 4190 4528 4198 4531
rect 4246 4528 4254 4531
rect 4310 4531 4314 4533
rect 4302 4528 4314 4531
rect 4478 4528 4481 4538
rect 4766 4528 4785 4531
rect 5190 4528 5193 4538
rect 61 4518 62 4522
rect 590 4518 598 4521
rect 990 4521 993 4528
rect 990 4518 1007 4521
rect 1229 4518 1230 4522
rect 1770 4518 1771 4522
rect 2894 4521 2897 4528
rect 2894 4518 2905 4521
rect 4994 4518 5001 4521
rect 848 4503 850 4507
rect 854 4503 857 4507
rect 861 4503 864 4507
rect 1872 4503 1874 4507
rect 1878 4503 1881 4507
rect 1885 4503 1888 4507
rect 2888 4503 2890 4507
rect 2894 4503 2897 4507
rect 2901 4503 2904 4507
rect 3920 4503 3922 4507
rect 3926 4503 3929 4507
rect 3933 4503 3936 4507
rect 4936 4503 4938 4507
rect 4942 4503 4945 4507
rect 4949 4503 4952 4507
rect 98 4488 105 4491
rect 302 4488 310 4491
rect 862 4488 870 4491
rect 1381 4488 1382 4492
rect 2910 4488 2921 4491
rect 3037 4488 3038 4492
rect 54 4468 65 4471
rect 150 4471 153 4481
rect 454 4478 465 4481
rect 134 4468 153 4471
rect 190 4468 214 4471
rect 446 4468 454 4471
rect 486 4468 505 4471
rect 586 4468 601 4471
rect 694 4468 705 4471
rect 1054 4471 1057 4481
rect 1266 4478 1273 4481
rect 1462 4478 1481 4481
rect 1646 4478 1665 4481
rect 1670 4472 1673 4481
rect 1814 4478 1833 4481
rect 1966 4478 1977 4481
rect 2134 4478 2146 4481
rect 2438 4478 2449 4481
rect 2486 4478 2498 4481
rect 2910 4481 2913 4488
rect 2894 4478 2913 4481
rect 1966 4477 1970 4478
rect 2142 4477 2146 4478
rect 2494 4477 2498 4478
rect 1054 4468 1081 4471
rect 1154 4468 1166 4471
rect 1342 4468 1385 4471
rect 1394 4468 1401 4471
rect 1982 4468 1993 4471
rect 2638 4468 2657 4471
rect 2738 4468 2745 4471
rect 62 4462 65 4468
rect 3078 4471 3081 4478
rect 3094 4472 3097 4481
rect 3558 4478 3577 4481
rect 3678 4478 3689 4481
rect 4006 4478 4017 4481
rect 4214 4478 4226 4481
rect 3678 4477 3682 4478
rect 2870 4468 2881 4471
rect 3078 4468 3089 4471
rect 3142 4468 3153 4471
rect 3254 4471 3258 4474
rect 3246 4468 3258 4471
rect 3426 4468 3433 4471
rect 3518 4468 3534 4471
rect 3550 4468 3558 4471
rect 3910 4471 3913 4478
rect 4006 4477 4010 4478
rect 4222 4477 4226 4478
rect 4486 4478 4505 4481
rect 4710 4478 4726 4481
rect 3910 4468 3922 4471
rect 4046 4468 4054 4471
rect 4254 4468 4257 4478
rect 4710 4474 4714 4478
rect 4506 4468 4513 4471
rect 5182 4468 5190 4471
rect 338 4458 345 4461
rect 606 4458 625 4461
rect 650 4458 657 4461
rect 662 4458 694 4461
rect 794 4458 801 4461
rect 890 4458 897 4461
rect 1002 4458 1028 4461
rect 1186 4458 1201 4461
rect 2878 4462 2881 4468
rect 3150 4462 3153 4468
rect 1858 4458 1870 4461
rect 2030 4458 2049 4461
rect 2110 4458 2118 4461
rect 2126 4458 2134 4461
rect 2194 4458 2201 4461
rect 2318 4458 2334 4461
rect 2410 4458 2417 4461
rect 2622 4458 2641 4461
rect 2678 4458 2686 4461
rect 2706 4458 2713 4461
rect 2950 4458 2958 4461
rect 3226 4458 3233 4461
rect 3530 4458 3537 4461
rect 4154 4458 4169 4461
rect 4394 4458 4409 4461
rect 4470 4458 4478 4461
rect 4578 4458 4593 4461
rect 4658 4458 4673 4461
rect 4678 4458 4698 4461
rect 4746 4458 4753 4461
rect 4946 4458 4961 4461
rect 898 4448 902 4452
rect 1786 4448 1793 4451
rect 2046 4448 2049 4458
rect 2678 4448 2681 4458
rect 3194 4448 3198 4452
rect 3350 4448 3353 4458
rect 4694 4457 4698 4458
rect 4330 4448 4334 4452
rect 4422 4448 4449 4451
rect 910 4438 921 4441
rect 1114 4438 1121 4441
rect 2162 4438 2165 4442
rect 3086 4438 3094 4441
rect 2002 4418 2003 4422
rect 2666 4418 2667 4422
rect 2754 4418 2755 4422
rect 3698 4418 3699 4422
rect 4085 4418 4086 4422
rect 4410 4418 4411 4422
rect 4802 4418 4803 4422
rect 328 4403 330 4407
rect 334 4403 337 4407
rect 341 4403 344 4407
rect 1352 4403 1354 4407
rect 1358 4403 1361 4407
rect 1365 4403 1368 4407
rect 2384 4403 2386 4407
rect 2390 4403 2393 4407
rect 2397 4403 2400 4407
rect 3400 4403 3402 4407
rect 3406 4403 3409 4407
rect 3413 4403 3416 4407
rect 4424 4403 4426 4407
rect 4430 4403 4433 4407
rect 4437 4403 4440 4407
rect 434 4388 436 4392
rect 554 4388 555 4392
rect 830 4388 838 4391
rect 1914 4388 1915 4392
rect 2549 4388 2550 4392
rect 3954 4388 3955 4392
rect 14 4368 22 4371
rect 76 4368 78 4372
rect 230 4368 254 4371
rect 805 4368 806 4372
rect 1142 4371 1145 4381
rect 1126 4368 1145 4371
rect 1182 4371 1185 4381
rect 1182 4368 1202 4371
rect 2955 4368 2958 4372
rect 3381 4368 3382 4372
rect 3574 4368 3585 4371
rect 570 4358 577 4361
rect 1126 4358 1129 4368
rect 1198 4366 1202 4368
rect 4198 4366 4202 4368
rect 1718 4358 1729 4361
rect 1946 4358 1950 4362
rect 2682 4358 2686 4362
rect 3562 4358 3566 4362
rect 3786 4358 3790 4362
rect 1718 4356 1722 4358
rect 150 4348 161 4351
rect 310 4348 337 4351
rect 510 4348 518 4351
rect 606 4348 614 4351
rect 1238 4348 1257 4351
rect 1302 4348 1310 4351
rect 38 4338 49 4341
rect 94 4338 97 4348
rect 158 4342 161 4348
rect 334 4342 337 4348
rect 1406 4342 1409 4351
rect 1614 4348 1622 4351
rect 1730 4348 1737 4351
rect 1898 4348 1913 4351
rect 1930 4348 1945 4351
rect 2114 4348 2121 4351
rect 2238 4351 2241 4358
rect 2238 4348 2249 4351
rect 2358 4348 2390 4351
rect 2686 4348 2702 4351
rect 2918 4348 2934 4351
rect 2990 4348 3009 4351
rect 3410 4348 3425 4351
rect 4118 4348 4126 4351
rect 4166 4348 4174 4351
rect 166 4338 185 4341
rect 830 4338 838 4341
rect 958 4338 972 4341
rect 998 4338 1014 4341
rect 1214 4338 1225 4341
rect 1882 4338 1905 4341
rect 2194 4338 2201 4341
rect 2378 4338 2393 4341
rect 3213 4338 3214 4342
rect 3542 4338 3545 4348
rect 4230 4342 4233 4351
rect 4406 4348 4414 4351
rect 4818 4348 4833 4351
rect 4918 4348 4926 4351
rect 5122 4348 5137 4351
rect 3670 4338 3682 4341
rect 3854 4338 3862 4341
rect 470 4331 473 4338
rect 958 4332 961 4338
rect 470 4328 481 4331
rect 878 4328 886 4331
rect 1018 4328 1025 4331
rect 1042 4328 1049 4331
rect 1438 4331 1442 4333
rect 1406 4328 1425 4331
rect 1430 4328 1442 4331
rect 2342 4331 2346 4333
rect 2342 4328 2353 4331
rect 4054 4328 4062 4331
rect 4126 4328 4129 4338
rect 4558 4332 4561 4342
rect 4738 4338 4745 4341
rect 4910 4341 4913 4348
rect 4902 4338 4913 4341
rect 5278 4332 5282 4336
rect 4230 4328 4249 4331
rect 4366 4328 4385 4331
rect 4662 4328 4681 4331
rect 4926 4328 4945 4331
rect 1085 4318 1086 4322
rect 3882 4318 3883 4322
rect 4194 4318 4195 4322
rect 4942 4321 4945 4328
rect 4942 4318 4953 4321
rect 848 4303 850 4307
rect 854 4303 857 4307
rect 861 4303 864 4307
rect 1872 4303 1874 4307
rect 1878 4303 1881 4307
rect 1885 4303 1888 4307
rect 2888 4303 2890 4307
rect 2894 4303 2897 4307
rect 2901 4303 2904 4307
rect 3920 4303 3922 4307
rect 3926 4303 3929 4307
rect 3933 4303 3936 4307
rect 4936 4303 4938 4307
rect 4942 4303 4945 4307
rect 4949 4303 4952 4307
rect 170 4288 172 4292
rect 334 4288 350 4291
rect 789 4288 790 4292
rect 882 4288 889 4291
rect 1133 4288 1134 4292
rect 410 4278 417 4281
rect 45 4268 46 4272
rect 126 4268 137 4271
rect 226 4268 233 4271
rect 478 4262 481 4271
rect 638 4268 657 4271
rect 838 4268 854 4271
rect 934 4271 937 4281
rect 1318 4278 1337 4281
rect 1398 4272 1401 4281
rect 1406 4278 1414 4281
rect 2222 4272 2225 4281
rect 2382 4278 2409 4281
rect 3134 4278 3145 4281
rect 3182 4278 3193 4281
rect 3230 4278 3249 4281
rect 3366 4278 3377 4281
rect 3134 4277 3138 4278
rect 3366 4277 3370 4278
rect 922 4268 937 4271
rect 1102 4268 1113 4271
rect 1426 4268 1433 4271
rect 1470 4268 1481 4271
rect 2062 4268 2081 4271
rect 2166 4268 2177 4271
rect 2350 4268 2361 4271
rect 2430 4268 2449 4271
rect 2582 4271 2586 4274
rect 2574 4268 2586 4271
rect 2670 4268 2682 4271
rect 2778 4268 2785 4271
rect 2802 4268 2809 4271
rect 2862 4268 2870 4271
rect 2878 4268 2905 4271
rect 2958 4268 2969 4271
rect 398 4258 409 4261
rect 446 4258 462 4261
rect 542 4258 561 4261
rect 582 4258 590 4261
rect 798 4261 801 4268
rect 1102 4262 1105 4268
rect 754 4258 761 4261
rect 798 4258 809 4261
rect 1230 4258 1246 4261
rect 2174 4262 2177 4268
rect 1694 4258 1710 4261
rect 1910 4258 1918 4261
rect 2430 4258 2433 4268
rect 3006 4262 3009 4271
rect 3150 4268 3161 4271
rect 3394 4268 3417 4271
rect 3506 4268 3513 4271
rect 3586 4268 3593 4271
rect 3654 4268 3662 4271
rect 4082 4268 4089 4271
rect 4326 4268 4345 4271
rect 4374 4268 4385 4271
rect 4534 4268 4553 4271
rect 4614 4271 4617 4281
rect 4854 4278 4866 4281
rect 4962 4278 4977 4281
rect 4982 4278 5001 4281
rect 5082 4278 5089 4281
rect 5094 4278 5113 4281
rect 4862 4277 4866 4278
rect 4614 4268 4633 4271
rect 4950 4268 4974 4271
rect 2502 4258 2521 4261
rect 2830 4258 2849 4261
rect 2854 4258 2862 4261
rect 3186 4258 3193 4261
rect 3214 4258 3222 4261
rect 3382 4258 3417 4261
rect 3606 4258 3614 4261
rect 3646 4258 3654 4261
rect 3710 4258 3718 4261
rect 3730 4258 3737 4261
rect 3794 4258 3801 4261
rect 4070 4258 4089 4261
rect 4238 4258 4246 4261
rect 4430 4258 4446 4261
rect 4554 4258 4561 4261
rect 4690 4258 4705 4261
rect 4774 4258 4782 4261
rect 4790 4261 4793 4268
rect 4790 4258 4801 4261
rect 4834 4258 4841 4261
rect 4846 4258 4854 4261
rect 5238 4258 5246 4261
rect 1070 4256 1074 4258
rect 1062 4248 1073 4251
rect 1778 4248 1782 4252
rect 2438 4248 2441 4258
rect 2518 4248 2521 4258
rect 2818 4248 2822 4252
rect 2830 4248 2833 4258
rect 4562 4248 4566 4252
rect 629 4238 630 4242
rect 882 4238 889 4241
rect 946 4238 947 4242
rect 1693 4238 1694 4242
rect 1854 4238 1862 4241
rect 1947 4238 1950 4242
rect 2747 4238 2750 4242
rect 3634 4238 3635 4242
rect 3802 4238 3803 4242
rect 4666 4238 4669 4242
rect 218 4218 219 4222
rect 1501 4218 1502 4222
rect 1626 4218 1627 4222
rect 1813 4218 1814 4222
rect 1989 4218 1990 4222
rect 2474 4218 2475 4222
rect 3738 4218 3739 4222
rect 4170 4218 4171 4222
rect 4205 4218 4206 4222
rect 4266 4218 4267 4222
rect 4354 4218 4355 4222
rect 5045 4218 5046 4222
rect 5069 4218 5070 4222
rect 5154 4218 5155 4222
rect 328 4203 330 4207
rect 334 4203 337 4207
rect 341 4203 344 4207
rect 1352 4203 1354 4207
rect 1358 4203 1361 4207
rect 1365 4203 1368 4207
rect 2384 4203 2386 4207
rect 2390 4203 2393 4207
rect 2397 4203 2400 4207
rect 3400 4203 3402 4207
rect 3406 4203 3409 4207
rect 3413 4203 3416 4207
rect 4424 4203 4426 4207
rect 4430 4203 4433 4207
rect 4437 4203 4440 4207
rect 101 4188 102 4192
rect 362 4188 363 4192
rect 493 4188 494 4192
rect 549 4188 550 4192
rect 846 4188 854 4191
rect 1250 4188 1251 4192
rect 1509 4188 1510 4192
rect 1685 4188 1686 4192
rect 2642 4188 2643 4192
rect 2946 4188 2947 4192
rect 3797 4188 3798 4192
rect 4357 4188 4358 4192
rect 5202 4188 5203 4192
rect 5274 4188 5275 4192
rect 3026 4178 3027 4182
rect 4733 4178 4734 4182
rect 206 4168 222 4171
rect 618 4168 633 4171
rect 1890 4168 1891 4172
rect 4394 4168 4397 4172
rect 4922 4168 4945 4171
rect 134 4151 137 4161
rect 190 4158 209 4161
rect 310 4158 321 4161
rect 670 4158 678 4161
rect 1186 4158 1190 4162
rect 102 4148 121 4151
rect 118 4142 121 4148
rect 134 4148 153 4151
rect 278 4148 286 4151
rect 346 4148 361 4151
rect 698 4148 721 4151
rect 134 4142 137 4148
rect 1130 4148 1137 4151
rect 1198 4151 1201 4161
rect 1198 4148 1217 4151
rect 1262 4151 1265 4161
rect 1262 4148 1281 4151
rect 1446 4148 1462 4151
rect 1494 4151 1497 4161
rect 1478 4148 1497 4151
rect 1702 4151 1706 4153
rect 1902 4152 1905 4161
rect 2526 4158 2537 4161
rect 1690 4148 1706 4151
rect 1882 4148 1889 4151
rect 1926 4148 1934 4151
rect 2058 4148 2065 4151
rect 2090 4148 2097 4151
rect 2154 4148 2161 4151
rect 2358 4148 2377 4151
rect 2654 4151 2657 4161
rect 2654 4148 2673 4151
rect 2758 4151 2761 4161
rect 2802 4158 2806 4162
rect 2754 4148 2761 4151
rect 2958 4151 2961 4161
rect 5110 4153 5114 4158
rect 2938 4148 2945 4151
rect 2958 4148 2977 4151
rect 3154 4148 3169 4151
rect 3282 4148 3289 4151
rect 14 4138 33 4141
rect 702 4138 710 4141
rect 734 4138 745 4141
rect 762 4138 785 4141
rect 878 4138 902 4141
rect 1422 4138 1433 4141
rect 1542 4138 1561 4141
rect 2110 4138 2118 4141
rect 2358 4138 2366 4141
rect 2494 4138 2505 4141
rect 2922 4138 2937 4141
rect 3006 4138 3017 4141
rect 3086 4138 3089 4148
rect 3478 4142 3481 4151
rect 3150 4138 3158 4141
rect 3314 4138 3321 4141
rect 3326 4138 3346 4141
rect 3430 4138 3446 4141
rect 3510 4141 3513 4151
rect 3734 4148 3753 4151
rect 4030 4148 4038 4151
rect 4106 4148 4113 4151
rect 4358 4148 4366 4151
rect 4606 4142 4609 4151
rect 4754 4148 4761 4151
rect 4870 4142 4873 4151
rect 5158 4142 5161 4151
rect 3506 4138 3513 4141
rect 3730 4138 3737 4141
rect 3746 4138 3753 4141
rect 3902 4138 3930 4141
rect 4218 4138 4233 4141
rect 4462 4138 4490 4141
rect 4658 4138 4665 4141
rect 4810 4138 4817 4141
rect 5030 4138 5042 4141
rect 278 4131 281 4138
rect 270 4128 281 4131
rect 454 4131 458 4136
rect 442 4128 458 4131
rect 754 4128 777 4131
rect 818 4128 833 4131
rect 1566 4128 1569 4138
rect 2494 4136 2498 4138
rect 3342 4136 3346 4138
rect 2382 4128 2398 4131
rect 3182 4131 3186 4133
rect 3358 4132 3362 4136
rect 3174 4128 3186 4131
rect 3302 4128 3313 4131
rect 3462 4128 3481 4131
rect 3718 4131 3722 4133
rect 3718 4128 3729 4131
rect 4014 4131 4018 4133
rect 4014 4128 4025 4131
rect 4062 4128 4073 4131
rect 4246 4131 4250 4133
rect 4238 4128 4250 4131
rect 4574 4131 4578 4133
rect 4574 4128 4585 4131
rect 4590 4128 4609 4131
rect 4662 4128 4665 4138
rect 4902 4132 4905 4138
rect 4670 4128 4689 4131
rect 4870 4128 4889 4131
rect 4902 4128 4910 4132
rect 5126 4131 5130 4133
rect 5126 4128 5137 4131
rect 5142 4128 5161 4131
rect 60 4118 62 4122
rect 602 4118 604 4122
rect 946 4118 948 4122
rect 2173 4118 2174 4122
rect 4786 4118 4787 4122
rect 848 4103 850 4107
rect 854 4103 857 4107
rect 861 4103 864 4107
rect 1872 4103 1874 4107
rect 1878 4103 1881 4107
rect 1885 4103 1888 4107
rect 2888 4103 2890 4107
rect 2894 4103 2897 4107
rect 2901 4103 2904 4107
rect 3920 4103 3922 4107
rect 3926 4103 3929 4107
rect 3933 4103 3936 4107
rect 4936 4103 4938 4107
rect 4942 4103 4945 4107
rect 4949 4103 4952 4107
rect 132 4088 134 4092
rect 165 4088 166 4092
rect 454 4088 465 4091
rect 626 4088 627 4092
rect 462 4082 465 4088
rect 414 4078 430 4081
rect 750 4078 766 4081
rect 846 4078 873 4081
rect 1166 4078 1185 4081
rect 1318 4078 1337 4081
rect 1342 4078 1358 4081
rect 1542 4078 1561 4081
rect 1870 4078 1886 4081
rect 2014 4078 2026 4081
rect 414 4072 417 4078
rect 750 4074 754 4078
rect 2022 4077 2026 4078
rect 2286 4078 2297 4081
rect 2330 4078 2331 4082
rect 3198 4078 3209 4081
rect 3742 4078 3753 4081
rect 3870 4078 3881 4081
rect 4202 4078 4203 4082
rect 4330 4078 4337 4081
rect 4830 4078 4842 4081
rect 2286 4077 2290 4078
rect 3198 4077 3202 4078
rect 3870 4077 3874 4078
rect 4838 4077 4842 4078
rect 4734 4072 4738 4074
rect 174 4068 182 4071
rect 234 4068 249 4071
rect 554 4068 569 4071
rect 414 4058 433 4061
rect 582 4058 593 4061
rect 942 4062 945 4071
rect 1846 4068 1854 4071
rect 2354 4068 2361 4071
rect 2630 4068 2641 4071
rect 2678 4068 2686 4071
rect 3994 4068 4009 4071
rect 4146 4068 4153 4071
rect 922 4058 929 4061
rect 982 4058 990 4061
rect 1002 4058 1009 4061
rect 1346 4058 1377 4061
rect 1394 4058 1409 4061
rect 1470 4058 1489 4061
rect 1506 4058 1521 4061
rect 1826 4058 1833 4061
rect 1838 4058 1846 4061
rect 2230 4058 2238 4061
rect 2442 4058 2449 4061
rect 2630 4061 2633 4068
rect 2590 4058 2609 4061
rect 2614 4058 2633 4061
rect 2654 4058 2662 4061
rect 2698 4058 2705 4061
rect 2758 4058 2766 4061
rect 2790 4058 2809 4061
rect 2822 4058 2830 4061
rect 2946 4058 2953 4061
rect 3062 4058 3081 4061
rect 3214 4058 3222 4061
rect 3342 4058 3350 4061
rect 3390 4061 3393 4068
rect 3366 4058 3393 4061
rect 4262 4062 4265 4071
rect 4374 4068 4382 4071
rect 5102 4068 5110 4071
rect 3646 4058 3665 4061
rect 3682 4058 3697 4061
rect 3902 4058 3937 4061
rect 4038 4058 4046 4061
rect 4166 4058 4174 4061
rect 4226 4058 4241 4061
rect 5070 4058 5089 4061
rect 5098 4058 5121 4061
rect 5126 4058 5145 4061
rect 5234 4058 5249 4061
rect 590 4052 593 4058
rect 898 4048 902 4052
rect 1486 4048 1489 4058
rect 1498 4048 1502 4052
rect 2298 4048 2305 4051
rect 2590 4048 2593 4058
rect 2806 4048 2809 4058
rect 2818 4048 2822 4052
rect 3078 4048 3081 4058
rect 3542 4052 3546 4057
rect 3374 4048 3390 4051
rect 3634 4048 3638 4052
rect 3646 4048 3649 4058
rect 3934 4048 3937 4058
rect 5058 4048 5062 4052
rect 5070 4048 5073 4058
rect 5142 4048 5145 4058
rect 1626 4038 1629 4042
rect 1861 4038 1862 4042
rect 1981 4038 1982 4042
rect 3093 4038 3094 4042
rect 858 4018 873 4021
rect 1410 4018 1411 4022
rect 1805 4018 1806 4022
rect 2173 4018 2174 4022
rect 2370 4018 2371 4022
rect 2418 4018 2419 4022
rect 4242 4018 4243 4022
rect 328 4003 330 4007
rect 334 4003 337 4007
rect 341 4003 344 4007
rect 1352 4003 1354 4007
rect 1358 4003 1361 4007
rect 1365 4003 1368 4007
rect 2384 4003 2386 4007
rect 2390 4003 2393 4007
rect 2397 4003 2400 4007
rect 3400 4003 3402 4007
rect 3406 4003 3409 4007
rect 3413 4003 3416 4007
rect 4424 4003 4426 4007
rect 4430 4003 4433 4007
rect 4437 4003 4440 4007
rect 101 3988 102 3992
rect 541 3988 542 3992
rect 1034 3988 1035 3992
rect 1522 3988 1523 3992
rect 2106 3988 2107 3992
rect 3205 3988 3206 3992
rect 3394 3988 3395 3992
rect 4061 3988 4062 3992
rect 4362 3988 4363 3992
rect 5194 3988 5195 3992
rect 3093 3978 3094 3982
rect 3437 3978 3438 3982
rect 226 3968 265 3971
rect 458 3968 459 3972
rect 931 3968 934 3972
rect 1066 3968 1067 3972
rect 1290 3968 1291 3972
rect 2338 3968 2339 3972
rect 3330 3968 3331 3972
rect 4763 3968 4766 3972
rect 198 3961 201 3968
rect 30 3938 62 3941
rect 94 3941 97 3951
rect 150 3951 153 3961
rect 190 3958 201 3961
rect 242 3958 249 3961
rect 614 3958 622 3961
rect 134 3948 153 3951
rect 530 3948 537 3951
rect 642 3948 665 3951
rect 670 3948 686 3951
rect 90 3938 97 3941
rect 110 3938 121 3941
rect 406 3938 409 3948
rect 650 3938 657 3941
rect 706 3938 713 3941
rect 782 3941 785 3951
rect 982 3951 985 3961
rect 982 3948 1001 3951
rect 1138 3948 1145 3951
rect 1214 3948 1222 3951
rect 1234 3948 1241 3951
rect 1302 3951 1305 3961
rect 1302 3948 1321 3951
rect 1366 3948 1374 3951
rect 1422 3951 1425 3961
rect 1386 3948 1401 3951
rect 1406 3948 1425 3951
rect 1686 3951 1689 3961
rect 1686 3948 1705 3951
rect 1710 3948 1729 3951
rect 1782 3951 1785 3961
rect 1982 3958 1993 3961
rect 2002 3958 2006 3962
rect 2034 3958 2038 3962
rect 1782 3948 1801 3951
rect 2130 3948 2137 3951
rect 2158 3948 2177 3951
rect 2182 3948 2190 3951
rect 758 3938 777 3941
rect 782 3938 798 3941
rect 814 3938 833 3941
rect 1438 3938 1446 3941
rect 1542 3941 1545 3948
rect 1542 3938 1553 3941
rect 1562 3938 1570 3941
rect 1726 3941 1729 3948
rect 2158 3942 2161 3948
rect 2350 3951 2353 3961
rect 2350 3948 2369 3951
rect 1726 3938 1737 3941
rect 2534 3938 2537 3948
rect 2990 3948 3006 3951
rect 3078 3951 3081 3961
rect 3062 3948 3081 3951
rect 3342 3951 3345 3961
rect 3406 3958 3422 3961
rect 3626 3958 3630 3962
rect 3342 3948 3361 3951
rect 3370 3948 3393 3951
rect 3502 3948 3510 3951
rect 3702 3951 3705 3961
rect 3714 3958 3718 3962
rect 4802 3958 4806 3962
rect 3674 3948 3681 3951
rect 3686 3948 3705 3951
rect 3786 3948 3793 3951
rect 4222 3951 4225 3958
rect 2894 3938 2918 3941
rect 3102 3938 3121 3941
rect 3261 3938 3262 3942
rect 3822 3938 3834 3941
rect 4118 3941 4121 3948
rect 4222 3948 4233 3951
rect 4110 3938 4121 3941
rect 4270 3941 4273 3948
rect 4814 3951 4817 3961
rect 5002 3958 5006 3962
rect 4814 3948 4833 3951
rect 4974 3948 4982 3951
rect 5074 3948 5081 3951
rect 4230 3938 4241 3941
rect 4262 3938 4273 3941
rect 4690 3938 4698 3941
rect 4862 3938 4881 3941
rect 110 3932 113 3938
rect 758 3928 761 3938
rect 814 3928 817 3938
rect 2246 3932 2250 3936
rect 2402 3928 2409 3931
rect 2678 3931 2682 3933
rect 2678 3928 2689 3931
rect 2806 3928 2825 3931
rect 3470 3931 3473 3938
rect 3450 3928 3457 3931
rect 3462 3928 3473 3931
rect 3502 3928 3513 3931
rect 3966 3928 3985 3931
rect 4214 3931 4218 3933
rect 4598 3932 4602 3936
rect 4214 3928 4225 3931
rect 1429 3918 1430 3922
rect 4322 3918 4323 3922
rect 848 3903 850 3907
rect 854 3903 857 3907
rect 861 3903 864 3907
rect 1872 3903 1874 3907
rect 1878 3903 1881 3907
rect 1885 3903 1888 3907
rect 2888 3903 2890 3907
rect 2894 3903 2897 3907
rect 2901 3903 2904 3907
rect 3920 3903 3922 3907
rect 3926 3903 3929 3907
rect 3933 3903 3936 3907
rect 4936 3903 4938 3907
rect 4942 3903 4945 3907
rect 4949 3903 4952 3907
rect 814 3888 822 3891
rect 3290 3888 3291 3892
rect 3422 3888 3433 3891
rect 357 3878 358 3882
rect 614 3878 630 3881
rect 614 3874 618 3878
rect 46 3868 62 3871
rect 310 3868 318 3871
rect 558 3868 566 3871
rect 890 3868 891 3872
rect 958 3871 961 3881
rect 1126 3878 1145 3881
rect 958 3868 977 3871
rect 1070 3868 1078 3871
rect 1098 3868 1105 3871
rect 1630 3871 1633 3881
rect 1662 3872 1665 3881
rect 2062 3878 2073 3881
rect 1614 3868 1633 3871
rect 1878 3868 1886 3871
rect 2022 3868 2030 3871
rect 2246 3868 2254 3871
rect 2278 3871 2281 3881
rect 2838 3872 2841 3881
rect 3022 3878 3033 3881
rect 3422 3881 3425 3888
rect 3174 3878 3186 3881
rect 3358 3878 3369 3881
rect 3406 3878 3425 3881
rect 3670 3878 3689 3881
rect 3990 3878 4002 3881
rect 4158 3878 4170 3881
rect 4434 3878 4449 3881
rect 4454 3878 4473 3881
rect 5198 3878 5210 3881
rect 3022 3877 3026 3878
rect 3182 3877 3186 3878
rect 3998 3877 4002 3878
rect 4166 3877 4170 3878
rect 5206 3877 5210 3878
rect 4638 3872 4642 3874
rect 2278 3868 2297 3871
rect 2706 3868 2721 3871
rect 3050 3868 3057 3871
rect 3390 3868 3401 3871
rect 3734 3868 3742 3871
rect 3902 3868 3910 3871
rect 3954 3868 3961 3871
rect 38 3858 46 3861
rect 94 3858 113 3861
rect 150 3858 158 3861
rect 302 3858 310 3861
rect 322 3858 345 3861
rect 398 3858 417 3861
rect 446 3858 458 3861
rect 538 3858 545 3861
rect 550 3858 569 3861
rect 1102 3862 1105 3868
rect 1154 3858 1161 3861
rect 1166 3858 1174 3861
rect 1390 3858 1409 3861
rect 1626 3858 1633 3861
rect 1742 3858 1750 3861
rect 1806 3858 1814 3861
rect 1950 3858 1977 3861
rect 2358 3858 2374 3861
rect 2630 3858 2638 3861
rect 2874 3858 2902 3861
rect 3038 3858 3057 3861
rect 3150 3858 3169 3861
rect 3234 3858 3241 3861
rect 3882 3858 3889 3861
rect 3894 3858 3902 3861
rect 3922 3858 3929 3861
rect 4118 3858 4137 3861
rect 4366 3858 4385 3861
rect 4574 3858 4606 3861
rect 4934 3858 4969 3861
rect 94 3848 97 3858
rect 454 3856 458 3858
rect 146 3848 150 3852
rect 254 3848 262 3851
rect 298 3848 302 3852
rect 542 3848 545 3858
rect 998 3848 1009 3851
rect 1390 3848 1393 3858
rect 2626 3848 2630 3852
rect 3858 3848 3862 3852
rect 4118 3848 4121 3858
rect 4366 3848 4369 3858
rect 4846 3852 4850 3854
rect 1006 3842 1009 3848
rect 117 3838 118 3842
rect 2606 3838 2618 3841
rect 3546 3838 3547 3842
rect 5074 3838 5077 3842
rect 5226 3838 5229 3842
rect 4866 3828 4867 3832
rect 1445 3818 1446 3822
rect 1730 3818 1731 3822
rect 1765 3818 1766 3822
rect 1914 3818 1915 3822
rect 1989 3818 1990 3822
rect 2114 3818 2115 3822
rect 2146 3818 2147 3822
rect 3101 3818 3102 3822
rect 4354 3818 4355 3822
rect 4514 3818 4515 3822
rect 4618 3818 4619 3822
rect 4970 3818 4971 3822
rect 5002 3818 5003 3822
rect 5189 3818 5190 3822
rect 328 3803 330 3807
rect 334 3803 337 3807
rect 341 3803 344 3807
rect 1352 3803 1354 3807
rect 1358 3803 1361 3807
rect 1365 3803 1368 3807
rect 2384 3803 2386 3807
rect 2390 3803 2393 3807
rect 2397 3803 2400 3807
rect 3400 3803 3402 3807
rect 3406 3803 3409 3807
rect 3413 3803 3416 3807
rect 4424 3803 4426 3807
rect 4430 3803 4433 3807
rect 4437 3803 4440 3807
rect 18 3788 19 3792
rect 282 3788 283 3792
rect 362 3788 363 3792
rect 3162 3788 3163 3792
rect 5109 3788 5110 3792
rect 114 3768 115 3772
rect 627 3768 630 3772
rect 1477 3768 1478 3772
rect 1858 3768 1859 3772
rect 2802 3768 2803 3772
rect 3930 3768 3946 3771
rect 4410 3768 4417 3771
rect 3030 3766 3034 3768
rect 70 3758 78 3761
rect 258 3758 265 3761
rect 398 3751 401 3758
rect 382 3748 401 3751
rect 782 3748 790 3751
rect 858 3748 865 3751
rect 922 3748 929 3751
rect 1222 3751 1225 3761
rect 1210 3748 1225 3751
rect 1390 3751 1393 3761
rect 1390 3748 1409 3751
rect 1462 3751 1465 3761
rect 1418 3748 1441 3751
rect 1446 3748 1465 3751
rect 1722 3748 1729 3751
rect 1870 3751 1873 3761
rect 1882 3758 1897 3761
rect 1870 3748 1905 3751
rect 1910 3748 1934 3751
rect 1942 3748 1958 3751
rect 2022 3748 2030 3751
rect 2042 3748 2049 3751
rect 2634 3748 2641 3751
rect 2742 3751 2745 3758
rect 2742 3748 2753 3751
rect 2774 3748 2782 3751
rect 2826 3748 2833 3751
rect 2990 3748 2998 3751
rect 406 3738 433 3741
rect 438 3738 457 3741
rect 886 3738 905 3741
rect 1342 3738 1358 3741
rect 1582 3738 1593 3741
rect 1922 3738 1929 3741
rect 2246 3741 2249 3748
rect 3462 3748 3470 3751
rect 3486 3748 3494 3751
rect 3918 3751 3921 3761
rect 4358 3752 4361 3761
rect 4802 3758 4806 3762
rect 3918 3748 3953 3751
rect 4062 3748 4070 3751
rect 4110 3748 4118 3751
rect 4254 3748 4270 3751
rect 4382 3748 4398 3751
rect 4562 3748 4569 3751
rect 4814 3751 4817 3761
rect 4794 3748 4801 3751
rect 4814 3748 4833 3751
rect 4966 3751 4969 3761
rect 4934 3748 4969 3751
rect 5042 3748 5057 3751
rect 2246 3738 2257 3741
rect 2294 3738 2313 3741
rect 2382 3738 2417 3741
rect 2422 3738 2449 3741
rect 2506 3738 2521 3741
rect 2534 3738 2553 3741
rect 2686 3738 2694 3741
rect 2986 3738 3009 3741
rect 3230 3738 3249 3741
rect 3526 3738 3537 3741
rect 4654 3741 4657 3748
rect 4654 3738 4673 3741
rect 886 3728 889 3738
rect 1582 3736 1586 3738
rect 1022 3731 1026 3736
rect 1010 3728 1026 3731
rect 1038 3731 1042 3733
rect 1766 3732 1770 3736
rect 1038 3728 1049 3731
rect 1614 3728 1625 3731
rect 1730 3728 1737 3731
rect 2126 3731 2129 3738
rect 2126 3728 2137 3731
rect 2294 3728 2297 3738
rect 2382 3728 2385 3738
rect 2534 3728 2537 3738
rect 3182 3731 3185 3738
rect 3526 3732 3529 3738
rect 3630 3736 3634 3738
rect 3182 3728 3193 3731
rect 3406 3728 3441 3731
rect 3742 3728 3761 3731
rect 4646 3728 4654 3731
rect 5206 3731 5210 3736
rect 5206 3728 5222 3731
rect 2498 3718 2499 3722
rect 2714 3718 2715 3722
rect 3786 3718 3787 3722
rect 4402 3718 4417 3721
rect 848 3703 850 3707
rect 854 3703 857 3707
rect 861 3703 864 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1885 3703 1888 3707
rect 2888 3703 2890 3707
rect 2894 3703 2897 3707
rect 2901 3703 2904 3707
rect 3920 3703 3922 3707
rect 3926 3703 3929 3707
rect 3933 3703 3936 3707
rect 4936 3703 4938 3707
rect 4942 3703 4945 3707
rect 4949 3703 4952 3707
rect 93 3688 94 3692
rect 2405 3688 2406 3692
rect 3530 3688 3531 3692
rect 166 3668 182 3671
rect 230 3671 233 3681
rect 438 3678 457 3681
rect 654 3678 673 3681
rect 230 3668 249 3671
rect 302 3668 318 3671
rect 758 3671 761 3681
rect 990 3678 1009 3681
rect 1014 3672 1017 3681
rect 742 3668 761 3671
rect 1074 3668 1075 3672
rect 1174 3668 1185 3671
rect 1214 3668 1233 3671
rect 1410 3668 1425 3671
rect 1518 3668 1529 3671
rect 1774 3668 1785 3671
rect 1854 3668 1889 3671
rect 1942 3668 1950 3671
rect 2006 3671 2009 3681
rect 2150 3672 2153 3681
rect 2806 3678 2825 3681
rect 3102 3678 3114 3681
rect 3350 3678 3362 3681
rect 1990 3668 2009 3671
rect 2062 3668 2073 3671
rect 2154 3668 2169 3671
rect 2246 3668 2249 3678
rect 3110 3677 3114 3678
rect 3358 3677 3362 3678
rect 2478 3668 2489 3671
rect 2594 3668 2601 3671
rect 2774 3668 2782 3671
rect 46 3658 54 3661
rect 390 3658 398 3661
rect 582 3661 585 3668
rect 574 3658 585 3661
rect 690 3658 697 3661
rect 1446 3658 1465 3661
rect 1518 3661 1521 3668
rect 1506 3658 1521 3661
rect 1862 3658 1870 3661
rect 2510 3658 2537 3661
rect 2722 3658 2737 3661
rect 2778 3658 2785 3661
rect 2842 3658 2849 3661
rect 2862 3661 2865 3671
rect 2966 3668 2974 3671
rect 2998 3668 3017 3671
rect 3078 3668 3086 3671
rect 3466 3668 3481 3671
rect 3606 3671 3609 3681
rect 4390 3678 4398 3681
rect 4430 3678 4446 3681
rect 3602 3668 3609 3671
rect 2862 3658 2870 3661
rect 2982 3658 2985 3668
rect 3078 3658 3097 3661
rect 3638 3662 3641 3671
rect 4078 3668 4086 3671
rect 4302 3668 4318 3671
rect 4830 3668 4838 3671
rect 5082 3668 5089 3671
rect 3702 3658 3710 3661
rect 3814 3658 3822 3661
rect 3894 3658 3910 3661
rect 3970 3658 3985 3661
rect 4126 3658 4134 3661
rect 4242 3658 4249 3661
rect 4370 3658 4377 3661
rect 4418 3658 4425 3661
rect 5046 3658 5065 3661
rect 5070 3658 5078 3661
rect 5082 3658 5097 3661
rect 5102 3658 5121 3661
rect 5270 3658 5278 3661
rect 1446 3648 1449 3658
rect 1586 3648 1590 3652
rect 1618 3648 1622 3652
rect 1806 3648 1825 3651
rect 2394 3648 2401 3651
rect 2706 3648 2710 3652
rect 2930 3648 2934 3652
rect 4018 3648 4022 3652
rect 4030 3648 4038 3651
rect 4326 3648 4345 3651
rect 5046 3648 5049 3658
rect 5118 3648 5121 3658
rect 5130 3648 5134 3652
rect 1653 3638 1654 3642
rect 4157 3638 4158 3642
rect 3986 3628 3987 3632
rect 878 3618 894 3621
rect 1501 3618 1502 3622
rect 1794 3618 1795 3622
rect 2765 3618 2766 3622
rect 2882 3618 2883 3622
rect 3218 3618 3219 3622
rect 3325 3618 3326 3622
rect 3813 3618 3814 3622
rect 4189 3618 4190 3622
rect 4357 3618 4358 3622
rect 4890 3618 4891 3622
rect 5290 3618 5291 3622
rect 328 3603 330 3607
rect 334 3603 337 3607
rect 341 3603 344 3607
rect 1352 3603 1354 3607
rect 1358 3603 1361 3607
rect 1365 3603 1368 3607
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2397 3603 2400 3607
rect 3400 3603 3402 3607
rect 3406 3603 3409 3607
rect 3413 3603 3416 3607
rect 4424 3603 4426 3607
rect 4430 3603 4433 3607
rect 4437 3603 4440 3607
rect 2978 3588 2979 3592
rect 3477 3588 3478 3592
rect 5149 3588 5150 3592
rect 3989 3578 3990 3582
rect 1021 3568 1022 3572
rect 1194 3568 1195 3572
rect 1770 3568 1771 3572
rect 2834 3568 2835 3572
rect 3173 3568 3174 3572
rect 4557 3568 4558 3572
rect 106 3558 113 3561
rect 562 3558 566 3562
rect 198 3548 206 3551
rect 122 3538 129 3541
rect 278 3538 286 3541
rect 294 3541 297 3551
rect 346 3548 377 3551
rect 798 3551 801 3561
rect 782 3548 801 3551
rect 1022 3548 1038 3551
rect 1094 3548 1102 3551
rect 1206 3551 1209 3561
rect 1206 3548 1225 3551
rect 1278 3548 1286 3551
rect 1366 3551 1369 3561
rect 1346 3548 1353 3551
rect 1366 3548 1401 3551
rect 1406 3548 1422 3551
rect 1518 3548 1537 3551
rect 1550 3548 1558 3551
rect 1614 3548 1622 3551
rect 1534 3542 1537 3548
rect 1814 3542 1817 3551
rect 1838 3548 1846 3551
rect 1894 3548 1902 3551
rect 1966 3548 1977 3551
rect 2166 3548 2174 3551
rect 2250 3548 2257 3551
rect 2306 3548 2313 3551
rect 2550 3551 2553 3561
rect 2594 3558 2598 3562
rect 2686 3561 2689 3568
rect 3670 3566 3674 3568
rect 2542 3548 2553 3551
rect 2646 3551 2649 3561
rect 2686 3558 2698 3561
rect 3542 3558 3550 3561
rect 4018 3558 4022 3562
rect 4490 3558 4494 3562
rect 4522 3558 4526 3562
rect 4686 3558 4694 3561
rect 2694 3556 2698 3558
rect 2630 3548 2649 3551
rect 1974 3542 1977 3548
rect 290 3538 297 3541
rect 574 3538 582 3541
rect 838 3538 862 3541
rect 990 3538 1001 3541
rect 1482 3538 1489 3541
rect 1498 3538 1505 3541
rect 1554 3538 1561 3541
rect 2038 3538 2054 3541
rect 2270 3538 2281 3541
rect 2374 3538 2398 3541
rect 2542 3541 2545 3548
rect 2534 3538 2545 3541
rect 2814 3538 2817 3548
rect 3034 3548 3041 3551
rect 3046 3548 3054 3551
rect 3194 3548 3201 3551
rect 3610 3548 3617 3551
rect 3738 3548 3745 3551
rect 3798 3548 3806 3551
rect 4022 3548 4030 3551
rect 4078 3548 4086 3551
rect 4170 3548 4177 3551
rect 4418 3548 4441 3551
rect 4606 3542 4609 3551
rect 4686 3548 4713 3551
rect 4746 3548 4753 3551
rect 4782 3548 4801 3551
rect 4934 3548 4961 3551
rect 5150 3548 5158 3551
rect 4934 3542 4937 3548
rect 2858 3538 2874 3541
rect 3101 3538 3102 3542
rect 3362 3538 3369 3541
rect 3526 3538 3534 3541
rect 3702 3538 3710 3541
rect 3718 3538 3737 3541
rect 4782 3538 4790 3541
rect 5006 3538 5025 3541
rect 318 3528 337 3531
rect 518 3528 537 3531
rect 878 3528 897 3531
rect 1950 3531 1954 3533
rect 1798 3528 1817 3531
rect 1950 3528 1961 3531
rect 2078 3528 2097 3531
rect 2494 3531 2498 3533
rect 2694 3531 2698 3533
rect 2166 3528 2177 3531
rect 2494 3528 2505 3531
rect 2686 3528 2698 3531
rect 3262 3531 3266 3533
rect 3254 3528 3266 3531
rect 3558 3531 3562 3533
rect 3550 3528 3562 3531
rect 4814 3531 4818 3533
rect 4806 3528 4818 3531
rect 4954 3528 4969 3531
rect 4974 3528 4977 3538
rect 5006 3528 5009 3538
rect 5182 3531 5186 3533
rect 5174 3528 5186 3531
rect 605 3518 606 3522
rect 3666 3518 3667 3522
rect 4725 3518 4726 3522
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 861 3503 864 3507
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1885 3503 1888 3507
rect 2888 3503 2890 3507
rect 2894 3503 2897 3507
rect 2901 3503 2904 3507
rect 3920 3503 3922 3507
rect 3926 3503 3929 3507
rect 3933 3503 3936 3507
rect 4936 3503 4938 3507
rect 4942 3503 4945 3507
rect 4949 3503 4952 3507
rect 1762 3488 1763 3492
rect 2149 3488 2150 3492
rect 2338 3488 2339 3492
rect 2362 3488 2363 3492
rect 2398 3488 2409 3491
rect 3157 3488 3158 3492
rect 4202 3488 4203 3492
rect 4674 3488 4675 3492
rect 22 3468 41 3471
rect 166 3462 169 3471
rect 326 3468 342 3471
rect 306 3458 313 3461
rect 534 3458 553 3461
rect 694 3462 697 3471
rect 1674 3468 1675 3472
rect 1710 3471 1714 3474
rect 1710 3468 1721 3471
rect 1878 3471 1881 3481
rect 2398 3481 2401 3488
rect 2222 3478 2234 3481
rect 2382 3478 2401 3481
rect 2506 3478 2513 3481
rect 2614 3478 2625 3481
rect 2981 3478 2982 3482
rect 3014 3478 3026 3481
rect 2230 3477 2234 3478
rect 2614 3477 2618 3478
rect 3022 3477 3026 3478
rect 3382 3478 3393 3481
rect 3398 3478 3406 3481
rect 3558 3478 3566 3481
rect 3622 3478 3641 3481
rect 3646 3478 3658 3481
rect 4062 3478 4081 3481
rect 4086 3478 4098 3481
rect 4270 3478 4289 3481
rect 3382 3477 3386 3478
rect 3654 3477 3658 3478
rect 4094 3477 4098 3478
rect 1878 3468 1913 3471
rect 2014 3471 2018 3474
rect 2014 3468 2025 3471
rect 2038 3468 2050 3471
rect 2642 3468 2649 3471
rect 3398 3468 3425 3471
rect 3830 3468 3841 3471
rect 758 3458 766 3461
rect 778 3458 785 3461
rect 934 3458 953 3461
rect 1222 3458 1241 3461
rect 1446 3458 1454 3461
rect 1514 3458 1521 3461
rect 1742 3458 1753 3461
rect 1878 3458 1894 3461
rect 2038 3462 2041 3468
rect 2170 3458 2177 3461
rect 2630 3458 2649 3461
rect 2838 3458 2857 3461
rect 2866 3458 2889 3461
rect 2894 3458 2929 3461
rect 2942 3458 2950 3461
rect 3278 3458 3286 3461
rect 3594 3458 3601 3461
rect 3622 3458 3625 3468
rect 3686 3458 3694 3461
rect 3790 3458 3809 3461
rect 4002 3458 4009 3461
rect 4034 3458 4041 3461
rect 4062 3458 4065 3468
rect 4206 3458 4225 3461
rect 4242 3458 4249 3461
rect 4446 3458 4481 3461
rect 4954 3458 4961 3461
rect 5006 3458 5025 3461
rect 5042 3458 5050 3461
rect 5090 3458 5105 3461
rect 5234 3458 5249 3461
rect 534 3448 537 3458
rect 950 3448 953 3458
rect 1238 3448 1241 3458
rect 1750 3452 1753 3458
rect 1578 3448 1582 3452
rect 2838 3448 2841 3458
rect 2926 3448 2929 3458
rect 3806 3448 3809 3458
rect 4206 3448 4209 3458
rect 4446 3457 4450 3458
rect 5006 3448 5009 3458
rect 5046 3457 5050 3458
rect 243 3438 246 3442
rect 1522 3438 1523 3442
rect 1691 3438 1694 3442
rect 2189 3438 2190 3442
rect 2250 3438 2253 3442
rect 3042 3438 3045 3442
rect 4114 3438 4117 3442
rect 5066 3438 5069 3442
rect 458 3418 459 3422
rect 2698 3418 2699 3422
rect 2941 3418 2942 3422
rect 3218 3418 3219 3422
rect 3434 3418 3435 3422
rect 4701 3418 4702 3422
rect 4946 3418 4961 3421
rect 328 3403 330 3407
rect 334 3403 337 3407
rect 341 3403 344 3407
rect 1352 3403 1354 3407
rect 1358 3403 1361 3407
rect 1365 3403 1368 3407
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2397 3403 2400 3407
rect 3400 3403 3402 3407
rect 3406 3403 3409 3407
rect 3413 3403 3416 3407
rect 4424 3403 4426 3407
rect 4430 3403 4433 3407
rect 4437 3403 4440 3407
rect 1549 3388 1550 3392
rect 1794 3388 1795 3392
rect 3709 3388 3710 3392
rect 3885 3388 3886 3392
rect 4565 3388 4566 3392
rect 4690 3388 4691 3392
rect 1517 3378 1518 3382
rect 354 3368 355 3372
rect 1443 3368 1446 3372
rect 4410 3368 4411 3372
rect 4422 3368 4438 3371
rect 4906 3368 4909 3372
rect 198 3358 206 3361
rect 366 3351 369 3361
rect 990 3352 993 3361
rect 1010 3358 1014 3362
rect 1274 3358 1278 3362
rect 338 3348 353 3351
rect 366 3348 385 3351
rect 606 3348 622 3351
rect 866 3348 881 3351
rect 1286 3351 1289 3361
rect 1502 3352 1505 3361
rect 1286 3348 1305 3351
rect 1310 3348 1318 3351
rect 1654 3351 1657 3361
rect 1666 3358 1670 3362
rect 3354 3358 3358 3362
rect 3586 3358 3590 3362
rect 1614 3348 1633 3351
rect 1638 3348 1657 3351
rect 526 3338 545 3341
rect 902 3338 921 3341
rect 1154 3338 1161 3341
rect 1614 3341 1617 3348
rect 1606 3338 1617 3341
rect 1858 3338 1866 3341
rect 2078 3341 2081 3348
rect 2318 3342 2321 3351
rect 2510 3348 2518 3351
rect 2742 3348 2750 3351
rect 2758 3348 2766 3351
rect 3494 3348 3513 3351
rect 3602 3348 3609 3351
rect 3614 3348 3622 3351
rect 3654 3348 3662 3351
rect 3742 3348 3758 3351
rect 3822 3348 3830 3351
rect 3870 3351 3873 3361
rect 3854 3348 3873 3351
rect 3906 3348 3913 3351
rect 4094 3351 4097 3358
rect 4086 3348 4097 3351
rect 4166 3348 4185 3351
rect 4250 3348 4257 3351
rect 4362 3348 4377 3351
rect 4518 3351 4521 3361
rect 4530 3358 4534 3362
rect 4510 3348 4521 3351
rect 4534 3348 4550 3351
rect 4614 3351 4617 3361
rect 4598 3348 4617 3351
rect 4738 3348 4745 3351
rect 4774 3348 4793 3351
rect 4938 3348 4945 3351
rect 2070 3338 2081 3341
rect 2466 3338 2473 3341
rect 3090 3338 3097 3341
rect 3366 3338 3374 3341
rect 3670 3338 3689 3341
rect 3718 3338 3729 3341
rect 3754 3338 3761 3341
rect 3926 3338 3942 3341
rect 4166 3338 4174 3341
rect 4510 3338 4513 3348
rect 4670 3338 4681 3341
rect 4710 3338 4718 3341
rect 4810 3338 4817 3341
rect 4838 3338 4857 3341
rect 526 3328 529 3338
rect 554 3328 561 3331
rect 718 3331 722 3336
rect 706 3328 722 3331
rect 902 3328 905 3338
rect 1574 3328 1582 3331
rect 1982 3328 2001 3331
rect 2302 3328 2321 3331
rect 2454 3331 2458 3333
rect 2454 3328 2465 3331
rect 2498 3328 2499 3332
rect 2646 3328 2665 3331
rect 3110 3331 3114 3333
rect 3102 3328 3114 3331
rect 3478 3331 3482 3333
rect 3478 3328 3489 3331
rect 4198 3331 4202 3333
rect 4194 3328 4202 3331
rect 4722 3328 4729 3331
rect 4798 3328 4806 3331
rect 4854 3328 4857 3338
rect 213 3318 214 3322
rect 1350 3318 1366 3321
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 861 3303 864 3307
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1885 3303 1888 3307
rect 2888 3303 2890 3307
rect 2894 3303 2897 3307
rect 2901 3303 2904 3307
rect 3920 3303 3922 3307
rect 3926 3303 3929 3307
rect 3933 3303 3936 3307
rect 4936 3303 4938 3307
rect 4942 3303 4945 3307
rect 4949 3303 4952 3307
rect 2714 3288 2715 3292
rect 230 3278 242 3281
rect 486 3278 498 3281
rect 858 3278 865 3281
rect 1046 3278 1057 3281
rect 1702 3278 1713 3281
rect 3254 3278 3273 3281
rect 3278 3278 3290 3281
rect 4202 3278 4209 3281
rect 4998 3278 5010 3281
rect 5110 3278 5129 3281
rect 5174 3278 5182 3281
rect 238 3277 242 3278
rect 494 3277 498 3278
rect 1046 3277 1050 3278
rect 1702 3277 1706 3278
rect 3222 3277 3226 3278
rect 3286 3277 3290 3278
rect 4622 3274 4626 3278
rect 5006 3277 5010 3278
rect 2334 3272 2338 3274
rect 214 3268 225 3271
rect 326 3268 354 3271
rect 462 3268 481 3271
rect 1062 3268 1073 3271
rect 1302 3268 1313 3271
rect 1598 3268 1609 3271
rect 1714 3268 1721 3271
rect 1730 3268 1737 3271
rect 2666 3268 2681 3271
rect 2698 3268 2705 3271
rect 4226 3268 4233 3271
rect 4694 3268 4706 3271
rect 4954 3268 4977 3271
rect 5130 3268 5137 3271
rect 702 3258 721 3261
rect 1086 3258 1094 3261
rect 1106 3258 1113 3261
rect 1302 3262 1305 3268
rect 1606 3262 1609 3268
rect 1470 3258 1478 3261
rect 1574 3258 1582 3261
rect 1798 3258 1806 3261
rect 2062 3258 2081 3261
rect 2086 3258 2110 3261
rect 2694 3258 2705 3261
rect 2822 3258 2830 3261
rect 2862 3258 2870 3261
rect 2982 3258 2993 3261
rect 3330 3258 3345 3261
rect 3418 3258 3425 3261
rect 3470 3258 3473 3268
rect 3606 3258 3614 3261
rect 3694 3258 3713 3261
rect 3894 3258 3918 3261
rect 4118 3258 4126 3261
rect 4190 3258 4198 3261
rect 4214 3258 4233 3261
rect 4326 3258 4334 3261
rect 4558 3258 4577 3261
rect 4882 3258 4897 3261
rect 4934 3258 4942 3261
rect 634 3248 638 3252
rect 718 3248 721 3258
rect 1570 3248 1574 3252
rect 2062 3248 2065 3258
rect 2702 3252 2705 3258
rect 2990 3252 2993 3258
rect 2306 3248 2310 3252
rect 3694 3248 3697 3258
rect 4326 3248 4329 3258
rect 4574 3248 4577 3258
rect 4586 3248 4590 3252
rect 4866 3248 4870 3252
rect 733 3238 734 3242
rect 1446 3238 1458 3241
rect 1469 3238 1470 3242
rect 1533 3238 1534 3242
rect 2050 3238 2051 3242
rect 2126 3238 2137 3241
rect 2318 3238 2329 3241
rect 3902 3238 3929 3241
rect 1821 3228 1822 3232
rect 2114 3228 2115 3232
rect 901 3218 902 3222
rect 1125 3218 1126 3222
rect 2861 3218 2862 3222
rect 3389 3218 3390 3222
rect 3429 3218 3430 3222
rect 3789 3218 3790 3222
rect 5194 3218 5195 3222
rect 328 3203 330 3207
rect 334 3203 337 3207
rect 341 3203 344 3207
rect 1352 3203 1354 3207
rect 1358 3203 1361 3207
rect 1365 3203 1368 3207
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2397 3203 2400 3207
rect 3400 3203 3402 3207
rect 3406 3203 3409 3207
rect 3413 3203 3416 3207
rect 4424 3203 4426 3207
rect 4430 3203 4433 3207
rect 4437 3203 4440 3207
rect 1674 3188 1675 3192
rect 2610 3188 2611 3192
rect 4125 3188 4126 3192
rect 5101 3188 5102 3192
rect 1386 3168 1387 3172
rect 2782 3168 2790 3171
rect 4538 3168 4539 3172
rect 3126 3166 3130 3168
rect 614 3151 617 3161
rect 762 3158 766 3162
rect 614 3148 633 3151
rect 766 3148 774 3151
rect 786 3148 793 3151
rect 910 3148 918 3151
rect 1082 3148 1089 3151
rect 1230 3151 1233 3161
rect 1418 3158 1422 3162
rect 1214 3148 1233 3151
rect 1378 3148 1385 3151
rect 1598 3151 1601 3161
rect 2346 3158 2350 3162
rect 2674 3158 2678 3162
rect 2830 3158 2838 3161
rect 1582 3148 1601 3151
rect 1614 3148 1622 3151
rect 1934 3148 1953 3151
rect 2214 3148 2230 3151
rect 2338 3148 2345 3151
rect 2414 3148 2422 3151
rect 2482 3148 2489 3151
rect 2526 3148 2534 3151
rect 2590 3148 2609 3151
rect 2658 3148 2673 3151
rect 3058 3148 3073 3151
rect 3210 3148 3217 3151
rect 3246 3148 3254 3151
rect 3358 3151 3361 3158
rect 3966 3153 3970 3158
rect 734 3138 742 3141
rect 806 3138 814 3141
rect 850 3138 865 3141
rect 1142 3138 1150 3141
rect 1166 3138 1174 3141
rect 1806 3138 1818 3141
rect 1946 3138 1953 3141
rect 2086 3141 2089 3148
rect 3358 3148 3369 3151
rect 3398 3148 3433 3151
rect 3450 3148 3465 3151
rect 3654 3151 3658 3153
rect 3654 3148 3673 3151
rect 3678 3148 3697 3151
rect 3702 3148 3710 3151
rect 3858 3148 3865 3151
rect 3870 3148 3897 3151
rect 4054 3148 4073 3151
rect 4178 3148 4193 3151
rect 4862 3151 4865 3161
rect 4846 3148 4865 3151
rect 4946 3148 4953 3151
rect 5070 3148 5086 3151
rect 5150 3148 5169 3151
rect 5178 3148 5185 3151
rect 2078 3138 2089 3141
rect 2226 3138 2233 3141
rect 2922 3138 2937 3141
rect 3366 3138 3385 3141
rect 3482 3138 3489 3141
rect 3538 3138 3545 3141
rect 3562 3138 3570 3141
rect 3710 3138 3729 3141
rect 3878 3138 3886 3141
rect 3906 3138 3921 3141
rect 4174 3138 4182 3141
rect 438 3128 457 3131
rect 1046 3128 1065 3131
rect 1078 3128 1081 3138
rect 1806 3132 1809 3138
rect 1910 3128 1929 3131
rect 2198 3131 2202 3133
rect 2198 3128 2209 3131
rect 2870 3128 2881 3131
rect 2966 3128 2985 3131
rect 3350 3131 3354 3133
rect 3350 3128 3361 3131
rect 3526 3128 3529 3138
rect 3710 3128 3713 3138
rect 3758 3131 3762 3133
rect 3750 3128 3762 3131
rect 3950 3131 3954 3133
rect 3926 3128 3954 3131
rect 4206 3131 4210 3133
rect 4198 3128 4210 3131
rect 4486 3128 4497 3131
rect 1910 3121 1913 3128
rect 1902 3118 1913 3121
rect 3122 3118 3123 3122
rect 3186 3118 3187 3122
rect 4346 3118 4347 3122
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 861 3103 864 3107
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1885 3103 1888 3107
rect 2888 3103 2890 3107
rect 2894 3103 2897 3107
rect 2901 3103 2904 3107
rect 3920 3103 3922 3107
rect 3926 3103 3929 3107
rect 3933 3103 3936 3107
rect 4936 3103 4938 3107
rect 4942 3103 4945 3107
rect 4949 3103 4952 3107
rect 1358 3088 1374 3091
rect 3934 3088 3953 3091
rect 3934 3082 3937 3088
rect 102 3078 121 3081
rect 190 3078 209 3081
rect 318 3078 337 3081
rect 342 3078 358 3081
rect 582 3071 585 3081
rect 566 3068 585 3071
rect 638 3071 641 3081
rect 790 3078 809 3081
rect 1118 3078 1129 3081
rect 2038 3078 2057 3081
rect 2158 3078 2169 3081
rect 2206 3078 2218 3081
rect 1118 3077 1122 3078
rect 1278 3077 1282 3078
rect 2214 3077 2218 3078
rect 622 3068 641 3071
rect 782 3068 798 3071
rect 1550 3068 1569 3071
rect 1658 3068 1665 3071
rect 1898 3068 1913 3071
rect 2058 3068 2065 3071
rect 2190 3068 2201 3071
rect 2446 3071 2449 3081
rect 2654 3078 2666 3081
rect 2918 3078 2930 3081
rect 3582 3078 3601 3081
rect 4642 3078 4649 3081
rect 4678 3078 4694 3081
rect 2662 3077 2666 3078
rect 2926 3077 2930 3078
rect 3494 3072 3498 3077
rect 3846 3072 3850 3077
rect 4678 3074 4682 3078
rect 2446 3068 2465 3071
rect 2806 3068 2817 3071
rect 3158 3068 3174 3071
rect 3310 3068 3321 3071
rect 3430 3068 3449 3071
rect 1130 3058 1137 3061
rect 1146 3058 1153 3061
rect 1398 3058 1406 3061
rect 1450 3058 1457 3061
rect 1758 3058 1766 3061
rect 1870 3058 1894 3061
rect 2418 3058 2425 3061
rect 2638 3061 2641 3068
rect 2638 3058 2649 3061
rect 2766 3058 2774 3061
rect 2798 3058 2814 3061
rect 2898 3058 2913 3061
rect 3318 3062 3321 3068
rect 3470 3062 3473 3071
rect 3602 3068 3609 3071
rect 4630 3068 4638 3071
rect 5126 3068 5129 3078
rect 5182 3068 5194 3071
rect 5242 3068 5243 3072
rect 3382 3058 3390 3061
rect 3886 3058 3902 3061
rect 4142 3058 4161 3061
rect 4214 3058 4222 3061
rect 4254 3058 4262 3061
rect 4278 3058 4297 3061
rect 4774 3058 4782 3061
rect 5042 3058 5057 3061
rect 1310 3048 1313 3058
rect 1482 3048 1489 3051
rect 3378 3048 3382 3052
rect 3722 3048 3726 3052
rect 3882 3048 3886 3052
rect 3938 3048 3953 3051
rect 4294 3048 4297 3058
rect 531 3038 534 3042
rect 1003 3038 1006 3042
rect 1099 3038 1102 3042
rect 2946 3038 2949 3042
rect 3862 3038 3874 3041
rect 4309 3038 4310 3042
rect 4901 3038 4902 3042
rect 4990 3038 5001 3041
rect 1578 3018 1579 3022
rect 1610 3018 1611 3022
rect 3034 3018 3035 3022
rect 3690 3018 3691 3022
rect 4021 3018 4022 3022
rect 4485 3018 4486 3022
rect 328 3003 330 3007
rect 334 3003 337 3007
rect 341 3003 344 3007
rect 1352 3003 1354 3007
rect 1358 3003 1361 3007
rect 1365 3003 1368 3007
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2397 3003 2400 3007
rect 3400 3003 3402 3007
rect 3406 3003 3409 3007
rect 3413 3003 3416 3007
rect 4424 3003 4426 3007
rect 4430 3003 4433 3007
rect 4437 3003 4440 3007
rect 2730 2968 2733 2972
rect 3675 2968 3678 2972
rect 3918 2968 3926 2971
rect 1078 2966 1082 2968
rect 3438 2966 3442 2968
rect 354 2948 361 2951
rect 378 2948 385 2951
rect 1102 2948 1129 2951
rect 1358 2948 1374 2951
rect 1654 2951 1657 2961
rect 3398 2958 3433 2961
rect 1626 2948 1633 2951
rect 1638 2948 1657 2951
rect 1730 2948 1745 2951
rect 2102 2951 2105 2958
rect 2086 2948 2105 2951
rect 2374 2948 2406 2951
rect 2606 2948 2614 2951
rect 3062 2948 3070 2951
rect 3134 2948 3142 2951
rect 3222 2942 3225 2951
rect 3470 2948 3478 2951
rect 3658 2948 3665 2951
rect 3710 2948 3729 2951
rect 4094 2948 4113 2951
rect 4166 2951 4169 2961
rect 4150 2948 4169 2951
rect 4182 2948 4198 2951
rect 4550 2948 4558 2951
rect 4626 2948 4641 2951
rect 4918 2951 4921 2961
rect 4902 2948 4921 2951
rect 5042 2948 5049 2951
rect 818 2938 826 2941
rect 1330 2938 1337 2941
rect 1606 2938 1625 2941
rect 2022 2938 2041 2941
rect 2054 2938 2073 2941
rect 2210 2938 2217 2941
rect 2518 2938 2545 2941
rect 2662 2938 2681 2941
rect 2694 2938 2702 2941
rect 2798 2938 2810 2941
rect 2954 2938 2969 2941
rect 3086 2938 3094 2941
rect 3602 2938 3610 2941
rect 3722 2938 3729 2941
rect 3966 2938 3985 2941
rect 4214 2938 4226 2941
rect 4566 2938 4574 2941
rect 4826 2938 4833 2941
rect 4946 2938 4958 2941
rect 334 2928 369 2931
rect 630 2928 649 2931
rect 658 2928 665 2931
rect 1141 2928 1142 2932
rect 1286 2928 1297 2931
rect 1414 2928 1433 2931
rect 1566 2931 1570 2933
rect 1566 2928 1577 2931
rect 2054 2928 2057 2938
rect 2110 2931 2114 2933
rect 2102 2928 2114 2931
rect 2294 2928 2313 2931
rect 2394 2928 2409 2931
rect 2414 2928 2433 2931
rect 2554 2928 2558 2932
rect 2678 2928 2681 2938
rect 2902 2928 2921 2931
rect 3238 2928 3246 2931
rect 3694 2931 3698 2933
rect 3694 2928 3705 2931
rect 3966 2928 3969 2938
rect 4222 2936 4226 2938
rect 4326 2928 4334 2931
rect 4582 2931 4586 2933
rect 4574 2928 4586 2931
rect 4814 2931 4818 2933
rect 4814 2928 4825 2931
rect 4858 2928 4859 2932
rect 5134 2928 5137 2938
rect 5142 2928 5161 2931
rect 1085 2918 1086 2922
rect 2902 2921 2905 2928
rect 2894 2918 2905 2921
rect 4205 2918 4206 2922
rect 4973 2918 4974 2922
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 861 2903 864 2907
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1885 2903 1888 2907
rect 2888 2903 2890 2907
rect 2894 2903 2897 2907
rect 2901 2903 2904 2907
rect 3920 2903 3922 2907
rect 3926 2903 3929 2907
rect 3933 2903 3936 2907
rect 4936 2903 4938 2907
rect 4942 2903 4945 2907
rect 4949 2903 4952 2907
rect 862 2888 870 2891
rect 2349 2888 2350 2892
rect 2902 2888 2913 2891
rect 3333 2888 3334 2892
rect 4450 2888 4465 2891
rect 346 2878 361 2881
rect 334 2868 361 2871
rect 358 2862 361 2868
rect 502 2862 505 2871
rect 654 2871 657 2881
rect 910 2878 929 2881
rect 990 2878 1009 2881
rect 1678 2878 1689 2881
rect 1774 2878 1793 2881
rect 1894 2878 1921 2881
rect 2062 2878 2081 2881
rect 1502 2874 1506 2878
rect 1678 2877 1682 2878
rect 1894 2877 1898 2878
rect 2278 2872 2281 2881
rect 2582 2878 2601 2881
rect 2718 2878 2729 2881
rect 2902 2881 2905 2888
rect 2886 2878 2905 2881
rect 3134 2878 3145 2881
rect 3294 2878 3313 2881
rect 3950 2878 3977 2881
rect 4342 2878 4354 2881
rect 2718 2877 2722 2878
rect 3134 2877 3138 2878
rect 3950 2877 3954 2878
rect 4350 2877 4354 2878
rect 654 2868 673 2871
rect 694 2868 713 2871
rect 950 2868 958 2871
rect 1322 2868 1338 2871
rect 1702 2868 1713 2871
rect 2298 2868 2305 2871
rect 2358 2868 2366 2871
rect 2730 2868 2745 2871
rect 2798 2868 2817 2871
rect 3754 2868 3761 2871
rect 3994 2868 4001 2871
rect 4150 2868 4158 2871
rect 4566 2871 4569 2881
rect 4598 2877 4602 2878
rect 4750 2876 4754 2878
rect 4550 2868 4569 2871
rect 4946 2868 4953 2871
rect 5198 2868 5210 2871
rect 222 2858 241 2861
rect 286 2858 305 2861
rect 438 2858 446 2861
rect 518 2858 534 2861
rect 550 2858 558 2861
rect 874 2858 889 2861
rect 1018 2858 1025 2861
rect 1030 2858 1057 2861
rect 1118 2858 1137 2861
rect 1290 2858 1297 2861
rect 1366 2858 1374 2861
rect 1702 2862 1705 2868
rect 1530 2858 1537 2861
rect 1642 2858 1649 2861
rect 2114 2858 2129 2861
rect 2286 2858 2305 2861
rect 2334 2858 2342 2861
rect 2414 2858 2422 2861
rect 2758 2858 2766 2861
rect 2870 2861 2873 2868
rect 2870 2858 2881 2861
rect 3078 2858 3094 2861
rect 3162 2858 3169 2861
rect 3354 2858 3361 2861
rect 3486 2858 3494 2861
rect 3594 2858 3601 2861
rect 3670 2858 3678 2861
rect 3742 2858 3761 2861
rect 3830 2861 3833 2868
rect 3822 2858 3833 2861
rect 3894 2858 3902 2861
rect 4094 2858 4102 2861
rect 4234 2858 4249 2861
rect 4650 2858 4657 2861
rect 4802 2858 4809 2861
rect 4870 2858 4889 2861
rect 5026 2858 5041 2861
rect 222 2848 225 2858
rect 274 2848 278 2852
rect 286 2848 289 2858
rect 362 2848 369 2851
rect 1134 2848 1137 2858
rect 1270 2848 1289 2851
rect 1690 2848 1697 2851
rect 4870 2848 4873 2858
rect 4962 2848 4966 2852
rect 5110 2851 5114 2854
rect 5102 2848 5114 2851
rect 843 2838 846 2842
rect 3658 2838 3661 2842
rect 4309 2838 4310 2842
rect 4778 2828 4779 2832
rect 613 2818 614 2822
rect 722 2818 723 2822
rect 754 2818 755 2822
rect 1058 2818 1059 2822
rect 1549 2818 1550 2822
rect 1930 2818 1931 2822
rect 2162 2818 2163 2822
rect 2789 2818 2790 2822
rect 328 2803 330 2807
rect 334 2803 337 2807
rect 341 2803 344 2807
rect 1352 2803 1354 2807
rect 1358 2803 1361 2807
rect 1365 2803 1368 2807
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2397 2803 2400 2807
rect 3400 2803 3402 2807
rect 3406 2803 3409 2807
rect 3413 2803 3416 2807
rect 4424 2803 4426 2807
rect 4430 2803 4433 2807
rect 4437 2803 4440 2807
rect 709 2788 710 2792
rect 1386 2788 1387 2792
rect 1538 2788 1539 2792
rect 2117 2788 2118 2792
rect 2773 2788 2774 2792
rect 5013 2788 5014 2792
rect 5294 2788 5302 2791
rect 1450 2768 1451 2772
rect 2154 2768 2155 2772
rect 3914 2768 3930 2771
rect 4734 2768 4742 2771
rect 1742 2766 1746 2768
rect 110 2748 129 2751
rect 182 2748 198 2751
rect 390 2751 393 2761
rect 954 2758 958 2762
rect 1082 2758 1086 2762
rect 374 2748 393 2751
rect 654 2748 662 2751
rect 798 2748 806 2751
rect 882 2748 889 2751
rect 934 2751 937 2758
rect 934 2748 945 2751
rect 1074 2748 1081 2751
rect 1150 2748 1158 2751
rect 542 2738 561 2741
rect 874 2738 881 2741
rect 942 2738 945 2748
rect 1398 2751 1401 2761
rect 1398 2748 1417 2751
rect 1462 2751 1465 2761
rect 1442 2748 1449 2751
rect 1462 2748 1481 2751
rect 1670 2751 1674 2753
rect 1670 2748 1686 2751
rect 1702 2751 1705 2761
rect 2562 2758 2569 2761
rect 1702 2748 1713 2751
rect 1758 2751 1761 2758
rect 1758 2748 1769 2751
rect 1834 2748 1841 2751
rect 2098 2748 2105 2751
rect 1574 2738 1577 2748
rect 1710 2742 1713 2748
rect 1714 2738 1721 2741
rect 1766 2738 1769 2748
rect 1842 2738 1849 2741
rect 2038 2741 2041 2748
rect 2062 2741 2065 2748
rect 2030 2738 2041 2741
rect 2054 2738 2065 2741
rect 2270 2738 2273 2748
rect 2410 2748 2417 2751
rect 2450 2748 2457 2751
rect 2546 2748 2553 2751
rect 2634 2748 2641 2751
rect 2750 2748 2758 2751
rect 2902 2748 2918 2751
rect 3054 2748 3062 2751
rect 3902 2751 3905 2761
rect 3902 2748 3937 2751
rect 3954 2748 3961 2751
rect 4014 2751 4017 2761
rect 4138 2758 4142 2762
rect 4218 2758 4222 2762
rect 4014 2748 4033 2751
rect 4222 2748 4230 2751
rect 4302 2751 4305 2761
rect 4690 2758 4694 2762
rect 4734 2758 4745 2761
rect 4334 2756 4338 2758
rect 4286 2748 4305 2751
rect 4378 2748 4393 2751
rect 4490 2748 4505 2751
rect 4546 2748 4553 2751
rect 4714 2748 4721 2751
rect 2430 2738 2438 2741
rect 2630 2738 2638 2741
rect 2794 2738 2801 2741
rect 2838 2738 2846 2741
rect 2982 2738 2990 2741
rect 3110 2738 3126 2741
rect 3198 2738 3206 2741
rect 3486 2738 3505 2741
rect 3950 2738 3958 2741
rect 3986 2738 3993 2741
rect 4014 2738 4022 2741
rect 94 2731 98 2733
rect 94 2728 105 2731
rect 542 2728 545 2738
rect 1542 2731 1545 2738
rect 1534 2728 1545 2731
rect 1862 2728 1897 2731
rect 2734 2731 2738 2733
rect 2734 2728 2745 2731
rect 3502 2728 3505 2738
rect 3622 2731 3626 2733
rect 3662 2732 3666 2736
rect 4478 2732 4481 2742
rect 4670 2738 4681 2741
rect 4742 2738 4745 2758
rect 4766 2751 4769 2761
rect 4926 2761 4929 2768
rect 4926 2758 4937 2761
rect 4942 2758 4958 2761
rect 4762 2748 4769 2751
rect 4998 2751 5001 2761
rect 4982 2748 5001 2751
rect 5062 2751 5065 2761
rect 5046 2748 5065 2751
rect 5078 2748 5086 2751
rect 5138 2748 5153 2751
rect 5238 2748 5249 2751
rect 5238 2742 5241 2748
rect 3622 2728 3633 2731
rect 2045 2718 2046 2722
rect 2181 2718 2182 2722
rect 2469 2718 2470 2722
rect 2829 2718 2830 2722
rect 2938 2718 2939 2722
rect 3902 2718 3910 2721
rect 4602 2718 4603 2722
rect 4754 2718 4755 2722
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 861 2703 864 2707
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1885 2703 1888 2707
rect 2888 2703 2890 2707
rect 2894 2703 2897 2707
rect 2901 2703 2904 2707
rect 3920 2703 3922 2707
rect 3926 2703 3929 2707
rect 3933 2703 3936 2707
rect 4936 2703 4938 2707
rect 4942 2703 4945 2707
rect 4949 2703 4952 2707
rect 141 2688 142 2692
rect 2358 2688 2369 2691
rect 5278 2688 5286 2691
rect 226 2678 233 2681
rect 1026 2678 1042 2681
rect 182 2668 190 2671
rect 210 2668 225 2671
rect 758 2671 761 2678
rect 1038 2674 1042 2678
rect 1054 2678 1065 2681
rect 1854 2678 1873 2681
rect 2058 2678 2065 2681
rect 2154 2678 2166 2681
rect 2358 2681 2361 2688
rect 2346 2678 2361 2681
rect 4062 2678 4074 2681
rect 4526 2678 4545 2681
rect 4662 2678 4673 2681
rect 4974 2678 4986 2681
rect 1054 2677 1058 2678
rect 4070 2677 4074 2678
rect 4662 2677 4666 2678
rect 4982 2677 4986 2678
rect 758 2668 769 2671
rect 858 2668 870 2671
rect 874 2668 881 2671
rect 1686 2668 1697 2671
rect 2002 2668 2009 2671
rect 2734 2668 2745 2671
rect 3034 2668 3041 2671
rect 3082 2668 3089 2671
rect 3346 2668 3361 2671
rect 3478 2668 3489 2671
rect 3670 2668 3681 2671
rect 3730 2668 3737 2671
rect 3902 2668 3910 2671
rect 4170 2668 4177 2671
rect 4366 2668 4377 2671
rect 4386 2668 4393 2671
rect 4674 2668 4681 2671
rect 4954 2668 4969 2671
rect 5182 2668 5194 2671
rect 222 2662 225 2668
rect 162 2658 169 2661
rect 174 2658 182 2661
rect 242 2658 257 2661
rect 270 2658 289 2661
rect 294 2658 302 2661
rect 438 2658 446 2661
rect 1146 2658 1161 2661
rect 1238 2658 1246 2661
rect 1330 2658 1337 2661
rect 1370 2658 1385 2661
rect 1406 2658 1409 2668
rect 1430 2658 1449 2661
rect 1686 2662 1689 2668
rect 1638 2658 1665 2661
rect 1742 2658 1750 2661
rect 2038 2658 2046 2661
rect 2162 2658 2169 2661
rect 2174 2658 2182 2661
rect 2230 2658 2257 2661
rect 2318 2658 2337 2661
rect 2614 2658 2622 2661
rect 2650 2658 2657 2661
rect 2694 2658 2713 2661
rect 2958 2658 2966 2661
rect 3054 2658 3062 2661
rect 3086 2661 3089 2668
rect 3486 2662 3489 2668
rect 3086 2658 3097 2661
rect 3218 2658 3225 2661
rect 3374 2658 3382 2661
rect 3458 2658 3465 2661
rect 3542 2661 3545 2668
rect 3490 2658 3497 2661
rect 3534 2658 3545 2661
rect 3862 2661 3865 2668
rect 3862 2658 3873 2661
rect 3882 2658 3889 2661
rect 3990 2658 3998 2661
rect 4346 2658 4353 2661
rect 4406 2658 4441 2661
rect 4606 2658 4622 2661
rect 4754 2658 4761 2661
rect 4778 2658 4793 2661
rect 4934 2658 4942 2661
rect 5222 2658 5238 2661
rect 154 2648 161 2651
rect 270 2648 273 2658
rect 802 2648 809 2651
rect 1334 2648 1337 2658
rect 1446 2648 1449 2658
rect 2710 2648 2713 2658
rect 2722 2648 2726 2652
rect 4438 2648 4441 2658
rect 4646 2652 4650 2657
rect 4758 2648 4761 2658
rect 4826 2648 4830 2652
rect 922 2638 923 2642
rect 4062 2641 4065 2648
rect 4054 2638 4065 2641
rect 845 2618 846 2622
rect 954 2618 955 2622
rect 1666 2618 1667 2622
rect 2093 2618 2094 2622
rect 2258 2618 2259 2622
rect 4234 2618 4235 2622
rect 4861 2618 4862 2622
rect 4885 2618 4886 2622
rect 328 2603 330 2607
rect 334 2603 337 2607
rect 341 2603 344 2607
rect 1352 2603 1354 2607
rect 1358 2603 1361 2607
rect 1365 2603 1368 2607
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2397 2603 2400 2607
rect 3400 2603 3402 2607
rect 3406 2603 3409 2607
rect 3413 2603 3416 2607
rect 4424 2603 4426 2607
rect 4430 2603 4433 2607
rect 4437 2603 4440 2607
rect 490 2588 491 2592
rect 2282 2588 2283 2592
rect 5269 2588 5270 2592
rect 334 2568 350 2571
rect 1291 2568 1294 2572
rect 1910 2568 1918 2571
rect 4242 2568 4249 2571
rect 114 2558 118 2562
rect 146 2558 150 2562
rect 274 2558 278 2562
rect 286 2551 289 2561
rect 810 2558 814 2562
rect 986 2558 990 2562
rect 286 2548 305 2551
rect 310 2548 318 2551
rect 366 2548 377 2551
rect 374 2542 377 2548
rect 438 2542 441 2551
rect 638 2548 646 2551
rect 814 2548 822 2551
rect 998 2551 1001 2561
rect 1342 2558 1358 2561
rect 1378 2558 1382 2562
rect 998 2548 1017 2551
rect 1022 2548 1041 2551
rect 1106 2548 1113 2551
rect 1174 2548 1182 2551
rect 1254 2548 1262 2551
rect 1346 2548 1377 2551
rect 1518 2548 1526 2551
rect 1574 2548 1582 2551
rect 1606 2548 1622 2551
rect 218 2538 219 2542
rect 318 2538 326 2541
rect 398 2538 425 2541
rect 830 2538 833 2548
rect 1038 2541 1041 2548
rect 1722 2548 1729 2551
rect 2050 2548 2057 2551
rect 2062 2548 2081 2551
rect 2138 2548 2145 2551
rect 2338 2548 2353 2551
rect 2486 2548 2494 2551
rect 2506 2548 2513 2551
rect 2554 2548 2561 2551
rect 2602 2548 2609 2551
rect 2642 2548 2649 2551
rect 2674 2548 2681 2551
rect 2870 2548 2878 2551
rect 3006 2548 3014 2551
rect 3090 2548 3097 2551
rect 3158 2548 3166 2551
rect 3410 2548 3433 2551
rect 3522 2548 3529 2551
rect 3670 2548 3678 2551
rect 4082 2548 4089 2551
rect 4170 2548 4177 2551
rect 4222 2548 4249 2551
rect 4398 2551 4401 2558
rect 4398 2548 4409 2551
rect 4478 2551 4481 2561
rect 4478 2548 4497 2551
rect 4554 2548 4569 2551
rect 4994 2548 5009 2551
rect 5078 2551 5081 2561
rect 5050 2548 5057 2551
rect 5062 2548 5081 2551
rect 5138 2548 5145 2551
rect 5150 2548 5158 2551
rect 5198 2548 5206 2551
rect 1038 2538 1049 2541
rect 1098 2538 1105 2541
rect 1206 2538 1214 2541
rect 1402 2538 1409 2541
rect 1470 2538 1478 2541
rect 1494 2538 1505 2541
rect 2422 2538 2430 2541
rect 2606 2541 2609 2548
rect 2606 2538 2617 2541
rect 2662 2538 2670 2541
rect 1550 2532 1553 2538
rect 1138 2528 1145 2531
rect 1546 2528 1553 2532
rect 2238 2528 2257 2531
rect 2262 2528 2270 2531
rect 2542 2531 2546 2533
rect 2542 2528 2553 2531
rect 2586 2528 2587 2532
rect 2638 2528 2649 2531
rect 2678 2528 2681 2548
rect 2698 2538 2713 2541
rect 2774 2538 2790 2541
rect 2850 2538 2857 2541
rect 2914 2538 2937 2541
rect 2954 2538 2969 2541
rect 3122 2538 3129 2541
rect 3158 2538 3161 2548
rect 3226 2538 3233 2541
rect 3446 2538 3454 2541
rect 3650 2538 3657 2541
rect 3766 2538 3793 2541
rect 4406 2541 4409 2548
rect 4406 2538 4417 2541
rect 4502 2538 4514 2541
rect 4510 2536 4514 2538
rect 2686 2528 2705 2531
rect 4126 2528 4134 2531
rect 4758 2528 4777 2531
rect 1878 2518 1894 2521
rect 2437 2518 2438 2522
rect 4154 2518 4155 2522
rect 4210 2518 4211 2522
rect 4946 2518 4953 2521
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 861 2503 864 2507
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1885 2503 1888 2507
rect 2888 2503 2890 2507
rect 2894 2503 2897 2507
rect 2901 2503 2904 2507
rect 3920 2503 3922 2507
rect 3926 2503 3929 2507
rect 3933 2503 3936 2507
rect 4936 2503 4938 2507
rect 4942 2503 4945 2507
rect 4949 2503 4952 2507
rect 2669 2488 2670 2492
rect 534 2478 553 2481
rect 558 2472 561 2481
rect 342 2468 350 2471
rect 358 2468 377 2471
rect 406 2468 417 2471
rect 438 2468 449 2471
rect 618 2468 625 2471
rect 702 2471 705 2478
rect 1414 2472 1417 2481
rect 1806 2478 1825 2481
rect 694 2468 705 2471
rect 162 2458 169 2461
rect 310 2458 329 2461
rect 358 2461 361 2468
rect 1238 2462 1241 2471
rect 1422 2468 1441 2471
rect 1462 2468 1473 2471
rect 1926 2468 1945 2471
rect 2006 2471 2009 2481
rect 1990 2468 2009 2471
rect 2086 2471 2089 2481
rect 4646 2478 4665 2481
rect 4770 2478 4777 2481
rect 4934 2478 4945 2481
rect 4950 2478 4978 2481
rect 2070 2468 2089 2471
rect 2434 2468 2449 2471
rect 2902 2468 2918 2471
rect 2954 2468 2961 2471
rect 3214 2468 3230 2471
rect 3410 2468 3425 2471
rect 3454 2468 3465 2471
rect 338 2458 361 2461
rect 734 2458 742 2461
rect 826 2458 833 2461
rect 874 2458 881 2461
rect 886 2458 894 2461
rect 1002 2458 1009 2461
rect 1118 2458 1126 2461
rect 1470 2462 1473 2468
rect 3494 2462 3497 2471
rect 3638 2468 3649 2471
rect 3686 2468 3694 2471
rect 4054 2468 4062 2471
rect 4086 2468 4094 2471
rect 4638 2471 4641 2478
rect 4934 2472 4937 2478
rect 4974 2477 4978 2478
rect 5270 2474 5274 2478
rect 4630 2468 4641 2471
rect 4726 2468 4737 2471
rect 4758 2468 4769 2471
rect 4766 2462 4769 2468
rect 1442 2458 1449 2461
rect 1946 2458 1953 2461
rect 1958 2458 1977 2461
rect 2134 2458 2142 2461
rect 2206 2458 2214 2461
rect 2310 2458 2318 2461
rect 3046 2458 3054 2461
rect 3082 2458 3089 2461
rect 3182 2458 3190 2461
rect 3390 2458 3433 2461
rect 3522 2458 3537 2461
rect 3566 2458 3593 2461
rect 3758 2458 3777 2461
rect 3806 2458 3849 2461
rect 3974 2458 3982 2461
rect 4190 2458 4206 2461
rect 4258 2458 4265 2461
rect 4374 2458 4401 2461
rect 4794 2458 4801 2461
rect 4918 2458 4926 2461
rect 5154 2458 5161 2461
rect 114 2448 118 2452
rect 154 2448 161 2451
rect 310 2448 313 2458
rect 1350 2452 1354 2457
rect 5174 2452 5178 2457
rect 666 2448 670 2452
rect 806 2448 825 2451
rect 1258 2448 1262 2452
rect 3882 2448 3886 2452
rect 4618 2448 4622 2452
rect 4802 2448 4806 2452
rect 4342 2442 4346 2444
rect 1066 2438 1067 2442
rect 949 2428 950 2432
rect 2373 2428 2374 2432
rect 2549 2428 2550 2432
rect 578 2418 579 2422
rect 1194 2418 1195 2422
rect 1597 2418 1598 2422
rect 1853 2418 1854 2422
rect 1898 2418 1899 2422
rect 2789 2418 2790 2422
rect 2938 2418 2939 2422
rect 3237 2418 3238 2422
rect 3629 2418 3630 2422
rect 3677 2418 3678 2422
rect 3733 2418 3734 2422
rect 3850 2418 3851 2422
rect 4266 2418 4267 2422
rect 328 2403 330 2407
rect 334 2403 337 2407
rect 341 2403 344 2407
rect 1352 2403 1354 2407
rect 1358 2403 1361 2407
rect 1365 2403 1368 2407
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2397 2403 2400 2407
rect 3400 2403 3402 2407
rect 3406 2403 3409 2407
rect 3413 2403 3416 2407
rect 4424 2403 4426 2407
rect 4430 2403 4433 2407
rect 4437 2403 4440 2407
rect 658 2388 659 2392
rect 746 2388 747 2392
rect 1381 2388 1382 2392
rect 1685 2388 1686 2392
rect 1714 2388 1715 2392
rect 1810 2388 1811 2392
rect 2026 2388 2027 2392
rect 2557 2388 2558 2392
rect 2661 2388 2662 2392
rect 2754 2388 2755 2392
rect 2781 2388 2782 2392
rect 2981 2388 2982 2392
rect 3770 2388 3771 2392
rect 5226 2388 5227 2392
rect 4298 2378 4299 2382
rect 619 2368 622 2372
rect 946 2368 947 2372
rect 2421 2368 2422 2372
rect 686 2358 705 2361
rect 110 2348 126 2351
rect 142 2338 145 2348
rect 374 2348 390 2351
rect 430 2351 434 2353
rect 430 2348 441 2351
rect 438 2342 441 2348
rect 958 2351 961 2361
rect 1138 2358 1142 2362
rect 1170 2358 1174 2362
rect 1342 2358 1369 2361
rect 1494 2358 1502 2361
rect 1778 2358 1785 2361
rect 1934 2353 1938 2358
rect 958 2348 977 2351
rect 1194 2348 1201 2351
rect 1206 2348 1214 2351
rect 1562 2348 1569 2351
rect 1754 2348 1761 2351
rect 1822 2348 1830 2351
rect 1862 2348 1878 2351
rect 1918 2351 1922 2353
rect 1902 2348 1922 2351
rect 2038 2351 2041 2361
rect 2102 2358 2110 2361
rect 3402 2358 3406 2362
rect 2038 2348 2057 2351
rect 2066 2348 2089 2351
rect 2130 2348 2145 2351
rect 2570 2348 2585 2351
rect 2866 2348 2873 2351
rect 2902 2348 2910 2351
rect 2982 2348 2990 2351
rect 3118 2348 3145 2351
rect 3406 2348 3433 2351
rect 3462 2348 3473 2351
rect 3430 2342 3433 2348
rect 478 2338 497 2341
rect 1710 2338 1729 2341
rect 1842 2338 1849 2341
rect 2202 2338 2209 2341
rect 2874 2338 2881 2341
rect 2950 2338 2961 2341
rect 3026 2338 3041 2341
rect 3066 2338 3073 2341
rect 3098 2338 3105 2341
rect 3230 2338 3257 2341
rect 3318 2338 3326 2341
rect 3338 2338 3345 2341
rect 3414 2338 3422 2341
rect 3502 2341 3505 2351
rect 3782 2351 3785 2361
rect 3782 2348 3801 2351
rect 3818 2348 3825 2351
rect 3850 2348 3857 2351
rect 4070 2348 4078 2351
rect 3502 2338 3518 2341
rect 3534 2338 3561 2341
rect 3566 2338 3593 2341
rect 3690 2338 3705 2341
rect 3822 2338 3825 2348
rect 4310 2351 4313 2361
rect 4310 2348 4329 2351
rect 4586 2348 4601 2351
rect 4762 2348 4777 2351
rect 4878 2348 4886 2351
rect 3962 2338 3969 2341
rect 4014 2338 4033 2341
rect 4422 2338 4454 2341
rect 4494 2338 4513 2341
rect 4998 2341 5001 2348
rect 5162 2348 5177 2351
rect 5282 2348 5289 2351
rect 4998 2338 5009 2341
rect 94 2331 98 2333
rect 94 2328 105 2331
rect 170 2328 171 2332
rect 430 2331 434 2333
rect 430 2328 441 2331
rect 494 2328 497 2338
rect 1581 2328 1582 2332
rect 1770 2328 1777 2331
rect 1862 2328 1889 2331
rect 2282 2328 2286 2332
rect 2597 2328 2598 2332
rect 2702 2328 2713 2331
rect 3082 2328 3086 2332
rect 3266 2328 3270 2332
rect 3718 2328 3729 2331
rect 3942 2328 3961 2331
rect 4014 2328 4017 2338
rect 4510 2328 4513 2338
rect 5126 2336 5130 2338
rect 1661 2318 1662 2322
rect 3522 2318 3523 2322
rect 4394 2318 4395 2322
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 861 2303 864 2307
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1885 2303 1888 2307
rect 2888 2303 2890 2307
rect 2894 2303 2897 2307
rect 2901 2303 2904 2307
rect 3920 2303 3922 2307
rect 3926 2303 3929 2307
rect 3933 2303 3936 2307
rect 4936 2303 4938 2307
rect 4942 2303 4945 2307
rect 4949 2303 4952 2307
rect 2701 2288 2702 2292
rect 2886 2288 2894 2291
rect 3309 2288 3310 2292
rect 3602 2288 3603 2292
rect 94 2278 105 2281
rect 94 2277 98 2278
rect 110 2268 121 2271
rect 190 2271 193 2281
rect 438 2278 457 2281
rect 654 2278 665 2281
rect 814 2278 833 2281
rect 1078 2278 1097 2281
rect 654 2277 658 2278
rect 1102 2272 1105 2281
rect 1490 2278 1497 2281
rect 1982 2278 1990 2281
rect 174 2268 193 2271
rect 678 2268 689 2271
rect 118 2262 121 2268
rect 290 2258 297 2261
rect 314 2258 345 2261
rect 678 2262 681 2268
rect 782 2262 785 2271
rect 1010 2268 1017 2271
rect 1070 2268 1078 2271
rect 1354 2268 1377 2271
rect 1422 2268 1430 2271
rect 1506 2268 1513 2271
rect 1870 2268 1905 2271
rect 1922 2268 1937 2271
rect 2182 2271 2185 2281
rect 3926 2278 3934 2281
rect 2182 2268 2201 2271
rect 2442 2268 2449 2271
rect 2498 2268 2505 2271
rect 2678 2268 2694 2271
rect 2790 2268 2809 2271
rect 3110 2268 3118 2271
rect 3142 2268 3150 2271
rect 666 2258 673 2261
rect 814 2258 817 2268
rect 1230 2258 1249 2261
rect 1298 2258 1305 2261
rect 1422 2258 1441 2261
rect 1534 2258 1553 2261
rect 1698 2258 1713 2261
rect 1718 2258 1737 2261
rect 2002 2258 2009 2261
rect 2718 2262 2722 2264
rect 2154 2258 2161 2261
rect 2634 2258 2641 2261
rect 2690 2258 2697 2261
rect 1230 2248 1233 2258
rect 1422 2248 1425 2258
rect 1534 2248 1537 2258
rect 1734 2248 1737 2258
rect 2694 2248 2697 2258
rect 2806 2248 2809 2268
rect 3510 2262 3513 2271
rect 3518 2268 3526 2271
rect 2934 2258 2942 2261
rect 3026 2258 3033 2261
rect 3242 2258 3249 2261
rect 3586 2258 3593 2261
rect 3878 2262 3881 2271
rect 3902 2268 3910 2271
rect 3918 2268 3926 2271
rect 4014 2268 4033 2271
rect 4210 2268 4217 2271
rect 4438 2268 4446 2271
rect 4518 2271 4521 2281
rect 4614 2278 4626 2281
rect 4622 2277 4626 2278
rect 4518 2268 4537 2271
rect 4750 2268 4758 2271
rect 4830 2271 4833 2281
rect 4814 2268 4833 2271
rect 5134 2271 5137 2281
rect 5278 2278 5289 2281
rect 5118 2268 5137 2271
rect 4006 2258 4014 2261
rect 4166 2258 4185 2261
rect 4278 2258 4297 2261
rect 4750 2258 4769 2261
rect 4778 2258 4793 2261
rect 4962 2258 4977 2261
rect 3946 2248 3953 2251
rect 4166 2248 4169 2258
rect 4294 2248 4297 2258
rect 4398 2252 4402 2257
rect 4306 2248 4310 2252
rect 4430 2248 4465 2251
rect 4606 2248 4614 2251
rect 1854 2238 1862 2241
rect 4422 2241 4426 2244
rect 4414 2238 4426 2241
rect 357 2218 358 2222
rect 981 2218 982 2222
rect 1218 2218 1219 2222
rect 1277 2218 1278 2222
rect 1682 2218 1683 2222
rect 2298 2218 2299 2222
rect 2525 2218 2526 2222
rect 3213 2218 3214 2222
rect 3570 2218 3571 2222
rect 3994 2218 3995 2222
rect 328 2203 330 2207
rect 334 2203 337 2207
rect 341 2203 344 2207
rect 1352 2203 1354 2207
rect 1358 2203 1361 2207
rect 1365 2203 1368 2207
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2397 2203 2400 2207
rect 3400 2203 3402 2207
rect 3406 2203 3409 2207
rect 3413 2203 3416 2207
rect 4424 2203 4426 2207
rect 4430 2203 4433 2207
rect 4437 2203 4440 2207
rect 1962 2188 1963 2192
rect 2245 2188 2246 2192
rect 3298 2188 3299 2192
rect 3965 2188 3966 2192
rect 4453 2188 4454 2192
rect 5154 2188 5155 2192
rect 5181 2188 5182 2192
rect 685 2178 686 2182
rect 147 2168 150 2172
rect 357 2168 358 2172
rect 866 2168 881 2171
rect 1206 2168 1218 2171
rect 1554 2168 1555 2172
rect 2306 2168 2307 2172
rect 1214 2166 1218 2168
rect 3862 2166 3866 2168
rect 4174 2166 4178 2168
rect 830 2151 833 2161
rect 842 2158 846 2162
rect 1890 2158 1897 2161
rect 2846 2158 2854 2161
rect 814 2148 833 2151
rect 1006 2148 1014 2151
rect 1098 2148 1105 2151
rect 1150 2148 1158 2151
rect 1362 2148 1374 2151
rect 1578 2148 1585 2151
rect 1650 2148 1657 2151
rect 2034 2148 2041 2151
rect 2134 2148 2142 2151
rect 2166 2148 2174 2151
rect 2258 2148 2265 2151
rect 2522 2148 2529 2151
rect 2566 2148 2574 2151
rect 2662 2148 2670 2151
rect 2790 2148 2801 2151
rect 2902 2148 2918 2151
rect 2998 2148 3017 2151
rect 198 2138 217 2141
rect 198 2128 201 2138
rect 286 2132 289 2142
rect 370 2138 377 2141
rect 694 2138 705 2141
rect 858 2138 870 2141
rect 966 2138 978 2141
rect 1078 2138 1097 2141
rect 1342 2138 1366 2141
rect 1606 2141 1609 2148
rect 1598 2138 1609 2141
rect 1622 2138 1641 2141
rect 1862 2138 1873 2141
rect 1934 2138 1942 2141
rect 2350 2141 2353 2148
rect 2342 2138 2353 2141
rect 2454 2138 2462 2141
rect 2498 2138 2505 2141
rect 2718 2138 2726 2141
rect 2790 2141 2793 2148
rect 3186 2148 3193 2151
rect 3394 2148 3417 2151
rect 3474 2148 3481 2151
rect 3538 2148 3545 2151
rect 3634 2148 3641 2151
rect 3774 2148 3793 2151
rect 3854 2151 3857 2161
rect 4182 2158 4201 2161
rect 3854 2148 3873 2151
rect 3930 2148 3950 2151
rect 4046 2148 4065 2151
rect 4130 2148 4137 2151
rect 4226 2148 4241 2151
rect 4254 2148 4270 2151
rect 4454 2148 4470 2151
rect 4478 2148 4497 2151
rect 4586 2148 4593 2151
rect 4710 2151 4713 2161
rect 4814 2153 4818 2158
rect 4694 2148 4713 2151
rect 2786 2138 2793 2141
rect 2998 2138 3006 2141
rect 3786 2138 3793 2141
rect 3854 2138 3862 2141
rect 4058 2138 4065 2141
rect 4254 2138 4257 2148
rect 5006 2148 5014 2151
rect 5126 2148 5134 2151
rect 390 2131 394 2133
rect 382 2128 394 2131
rect 1094 2128 1097 2138
rect 1326 2131 1330 2133
rect 1326 2128 1337 2131
rect 1658 2128 1665 2131
rect 1870 2131 1873 2138
rect 1870 2128 1886 2131
rect 3758 2131 3762 2133
rect 4078 2131 4082 2133
rect 3758 2128 3769 2131
rect 4070 2128 4082 2131
rect 4285 2128 4286 2132
rect 4326 2131 4330 2133
rect 4318 2128 4330 2131
rect 4878 2128 4897 2131
rect 4994 2128 4995 2132
rect 1221 2118 1222 2122
rect 2477 2118 2478 2122
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 861 2103 864 2107
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1885 2103 1888 2107
rect 2888 2103 2890 2107
rect 2894 2103 2897 2107
rect 2901 2103 2904 2107
rect 3920 2103 3922 2107
rect 3926 2103 3929 2107
rect 3933 2103 3936 2107
rect 4936 2103 4938 2107
rect 4942 2103 4945 2107
rect 4949 2103 4952 2107
rect 342 2088 350 2091
rect 3778 2088 3779 2092
rect 4210 2088 4211 2092
rect 5026 2088 5027 2092
rect 166 2078 177 2081
rect 262 2078 281 2081
rect 446 2078 462 2081
rect 918 2078 929 2081
rect 1134 2078 1153 2081
rect 1366 2081 1369 2088
rect 1342 2078 1369 2081
rect 166 2077 170 2078
rect 446 2074 450 2078
rect 194 2068 201 2071
rect 374 2068 393 2071
rect 430 2071 434 2074
rect 926 2072 929 2078
rect 422 2068 434 2071
rect 610 2068 617 2071
rect 854 2068 862 2071
rect 290 2058 305 2061
rect 398 2061 401 2068
rect 1370 2068 1385 2071
rect 1402 2068 1409 2071
rect 1430 2068 1438 2071
rect 1526 2068 1537 2071
rect 1590 2071 1593 2081
rect 1610 2078 1617 2081
rect 1638 2078 1649 2081
rect 1646 2072 1649 2078
rect 1574 2068 1593 2071
rect 1662 2068 1681 2071
rect 1890 2068 1905 2071
rect 2286 2068 2302 2071
rect 2822 2068 2825 2078
rect 2838 2074 2842 2078
rect 2854 2078 2865 2081
rect 2870 2078 2905 2081
rect 2974 2078 2986 2081
rect 3494 2078 3506 2081
rect 2854 2077 2858 2078
rect 2982 2077 2986 2078
rect 3502 2077 3506 2078
rect 2958 2068 2969 2071
rect 3318 2068 3326 2071
rect 3762 2068 3769 2071
rect 3870 2068 3878 2071
rect 3914 2068 3929 2071
rect 4054 2071 4057 2081
rect 4238 2077 4242 2078
rect 4862 2074 4866 2078
rect 4054 2068 4073 2071
rect 4078 2068 4105 2071
rect 4222 2068 4230 2071
rect 4686 2068 4694 2071
rect 398 2058 417 2061
rect 462 2058 470 2061
rect 586 2058 593 2061
rect 598 2058 614 2061
rect 782 2058 790 2061
rect 846 2058 870 2061
rect 882 2058 889 2061
rect 1298 2058 1305 2061
rect 1350 2058 1358 2061
rect 1466 2058 1473 2061
rect 1478 2058 1505 2061
rect 1550 2058 1558 2061
rect 1630 2061 1633 2068
rect 1622 2058 1633 2061
rect 1646 2058 1654 2061
rect 1874 2058 1902 2061
rect 1922 2058 1929 2061
rect 2034 2058 2041 2061
rect 2362 2058 2369 2061
rect 2798 2058 2814 2061
rect 3138 2058 3145 2061
rect 3186 2058 3201 2061
rect 3218 2058 3225 2061
rect 3250 2058 3257 2061
rect 3478 2061 3481 2068
rect 3478 2058 3489 2061
rect 3830 2058 3857 2061
rect 3862 2058 3870 2061
rect 4166 2058 4185 2061
rect 5086 2062 5089 2071
rect 4422 2058 4457 2061
rect 4574 2058 4593 2061
rect 4878 2058 4886 2061
rect 5162 2058 5177 2061
rect 178 2048 185 2051
rect 634 2048 636 2052
rect 810 2048 814 2052
rect 1942 2048 1945 2058
rect 2502 2052 2506 2054
rect 3798 2048 3817 2051
rect 4166 2048 4169 2058
rect 4346 2048 4350 2052
rect 4422 2048 4425 2058
rect 4574 2048 4577 2058
rect 4630 2048 4633 2058
rect 4650 2048 4654 2052
rect 362 2038 369 2041
rect 1837 2038 1838 2042
rect 1930 2038 1931 2042
rect 1965 2038 1966 2042
rect 2949 2038 2950 2042
rect 3082 2038 3089 2041
rect 3370 2038 3371 2042
rect 3522 2038 3525 2042
rect 4410 2038 4411 2042
rect 5138 2038 5141 2042
rect 1178 2028 1179 2032
rect 3202 2028 3203 2032
rect 781 2018 782 2022
rect 890 2018 891 2022
rect 1517 2018 1518 2022
rect 2725 2018 2726 2022
rect 2749 2018 2750 2022
rect 4482 2018 4483 2022
rect 4725 2018 4726 2022
rect 328 2003 330 2007
rect 334 2003 337 2007
rect 341 2003 344 2007
rect 1352 2003 1354 2007
rect 1358 2003 1361 2007
rect 1365 2003 1368 2007
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2397 2003 2400 2007
rect 3400 2003 3402 2007
rect 3406 2003 3409 2007
rect 3413 2003 3416 2007
rect 4424 2003 4426 2007
rect 4430 2003 4433 2007
rect 4437 2003 4440 2007
rect 301 1988 302 1992
rect 1602 1988 1603 1992
rect 1989 1988 1990 1992
rect 2138 1988 2139 1992
rect 2693 1988 2694 1992
rect 3525 1988 3526 1992
rect 4781 1988 4782 1992
rect 4869 1988 4870 1992
rect 1138 1978 1139 1982
rect 1333 1978 1334 1982
rect 3130 1978 3131 1982
rect 234 1968 235 1972
rect 414 1968 425 1971
rect 731 1968 734 1972
rect 1310 1968 1322 1971
rect 1826 1968 1833 1971
rect 2066 1968 2067 1972
rect 2766 1968 2774 1971
rect 3011 1968 3014 1972
rect 5066 1968 5073 1971
rect 414 1966 418 1968
rect 422 1962 425 1968
rect 390 1958 409 1961
rect 938 1958 945 1961
rect 110 1948 118 1951
rect 178 1948 185 1951
rect 214 1948 233 1951
rect 382 1948 390 1951
rect 566 1948 574 1951
rect 762 1948 769 1951
rect 1150 1951 1153 1961
rect 1318 1952 1321 1961
rect 1454 1958 1466 1961
rect 1890 1958 1897 1961
rect 2818 1958 2825 1961
rect 2842 1958 2849 1961
rect 2866 1958 2873 1961
rect 3050 1958 3054 1962
rect 3082 1958 3086 1962
rect 1462 1956 1466 1958
rect 1150 1948 1169 1951
rect 334 1938 342 1941
rect 526 1938 538 1941
rect 454 1932 458 1936
rect 590 1932 593 1942
rect 782 1938 790 1941
rect 1002 1938 1009 1941
rect 1214 1938 1217 1948
rect 1402 1948 1409 1951
rect 1426 1948 1441 1951
rect 1674 1948 1681 1951
rect 1686 1948 1697 1951
rect 1694 1942 1697 1948
rect 1794 1938 1825 1941
rect 1894 1941 1897 1948
rect 1842 1938 1849 1941
rect 1870 1938 1897 1941
rect 1910 1938 1913 1958
rect 2038 1948 2046 1951
rect 2058 1948 2065 1951
rect 2130 1948 2137 1951
rect 2350 1948 2358 1951
rect 2526 1948 2545 1951
rect 2622 1948 2641 1951
rect 2718 1948 2729 1951
rect 1950 1938 1969 1941
rect 2090 1938 2097 1941
rect 2454 1938 2470 1941
rect 2702 1938 2721 1941
rect 2822 1938 2825 1958
rect 2830 1948 2846 1951
rect 3166 1948 3185 1951
rect 3190 1948 3209 1951
rect 3262 1948 3270 1951
rect 3454 1948 3473 1951
rect 3670 1951 3674 1953
rect 3662 1948 3674 1951
rect 3454 1942 3457 1948
rect 3798 1948 3806 1951
rect 3886 1948 3902 1951
rect 4022 1948 4041 1951
rect 4326 1951 4329 1961
rect 4310 1948 4329 1951
rect 4622 1951 4625 1961
rect 4838 1958 4857 1961
rect 4606 1948 4625 1951
rect 4830 1951 4833 1958
rect 4782 1948 4809 1951
rect 4814 1948 4833 1951
rect 5038 1951 5041 1961
rect 5038 1948 5057 1951
rect 2906 1938 2913 1941
rect 3094 1938 3102 1941
rect 3110 1938 3121 1941
rect 3214 1938 3241 1941
rect 3254 1938 3262 1941
rect 3406 1938 3414 1941
rect 3466 1938 3473 1941
rect 3622 1938 3638 1941
rect 3758 1938 3770 1941
rect 4006 1938 4014 1941
rect 4322 1938 4329 1941
rect 4374 1938 4390 1941
rect 4878 1938 4889 1941
rect 5038 1938 5046 1941
rect 926 1931 930 1933
rect 926 1928 937 1931
rect 1646 1928 1665 1931
rect 2502 1931 2505 1938
rect 2502 1928 2513 1931
rect 2518 1928 2529 1931
rect 2546 1928 2553 1931
rect 2642 1928 2649 1931
rect 2702 1928 2705 1938
rect 2742 1928 2750 1931
rect 4014 1928 4017 1938
rect 4478 1932 4482 1936
rect 4518 1933 4522 1938
rect 4670 1931 4674 1933
rect 4662 1928 4674 1931
rect 4894 1928 4902 1931
rect 2805 1918 2806 1922
rect 2853 1918 2854 1922
rect 3418 1918 3433 1921
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 861 1903 864 1907
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1885 1903 1888 1907
rect 2888 1903 2890 1907
rect 2894 1903 2897 1907
rect 2901 1903 2904 1907
rect 3920 1903 3922 1907
rect 3926 1903 3929 1907
rect 3933 1903 3936 1907
rect 4936 1903 4938 1907
rect 4942 1903 4945 1907
rect 4949 1903 4952 1907
rect 1362 1888 1377 1891
rect 2290 1888 2292 1892
rect 3061 1888 3062 1892
rect 5194 1888 5195 1892
rect 5242 1888 5243 1892
rect 110 1878 129 1881
rect 514 1878 515 1882
rect 998 1878 1009 1881
rect 1550 1878 1558 1881
rect 998 1877 1002 1878
rect 338 1868 361 1871
rect 566 1868 577 1871
rect 882 1868 889 1871
rect 1026 1868 1033 1871
rect 126 1858 129 1868
rect 326 1858 342 1861
rect 1094 1862 1097 1871
rect 1398 1868 1409 1871
rect 1582 1871 1585 1881
rect 1790 1878 1802 1881
rect 2070 1878 2082 1881
rect 2198 1878 2209 1881
rect 2470 1878 2478 1881
rect 3406 1878 3414 1881
rect 1798 1877 1802 1878
rect 2078 1877 2082 1878
rect 2790 1874 2794 1878
rect 1566 1868 1585 1871
rect 1598 1868 1606 1871
rect 1766 1868 1774 1871
rect 1886 1868 1914 1871
rect 2062 1868 2073 1871
rect 2254 1868 2262 1871
rect 2070 1862 2073 1868
rect 3150 1862 3153 1871
rect 3246 1868 3254 1871
rect 3398 1868 3433 1871
rect 3630 1868 3638 1871
rect 3894 1871 3897 1881
rect 4094 1872 4097 1881
rect 4302 1878 4314 1881
rect 4310 1877 4314 1878
rect 5166 1872 5169 1881
rect 3890 1868 3897 1871
rect 4014 1868 4025 1871
rect 4070 1868 4094 1871
rect 4218 1868 4225 1871
rect 4278 1868 4286 1871
rect 4538 1868 4553 1871
rect 4014 1862 4017 1868
rect 774 1858 793 1861
rect 798 1858 806 1861
rect 1014 1858 1033 1861
rect 1126 1858 1134 1861
rect 1286 1858 1305 1861
rect 1718 1858 1737 1861
rect 1766 1858 1785 1861
rect 2326 1858 2353 1861
rect 2358 1858 2393 1861
rect 2478 1858 2505 1861
rect 2750 1858 2766 1861
rect 2838 1858 2857 1861
rect 2862 1858 2878 1861
rect 2926 1858 2942 1861
rect 2982 1858 2990 1861
rect 3014 1858 3033 1861
rect 3042 1858 3054 1861
rect 3266 1858 3273 1861
rect 3330 1858 3345 1861
rect 3630 1858 3649 1861
rect 3758 1858 3777 1861
rect 3822 1858 3830 1861
rect 3862 1858 3881 1861
rect 3902 1858 3910 1861
rect 4278 1858 4297 1861
rect 4438 1858 4473 1861
rect 4622 1861 4625 1871
rect 4862 1868 4870 1871
rect 4902 1868 4913 1871
rect 5066 1868 5073 1871
rect 4622 1858 4630 1861
rect 4714 1858 4721 1861
rect 4806 1861 4809 1868
rect 4910 1862 4913 1868
rect 4762 1858 4769 1861
rect 4782 1858 4801 1861
rect 4806 1858 4825 1861
rect 4998 1858 5006 1861
rect 5054 1858 5073 1861
rect 5106 1858 5113 1861
rect 5170 1858 5177 1861
rect 5254 1858 5273 1861
rect 774 1848 777 1858
rect 1286 1848 1289 1858
rect 2390 1848 2393 1858
rect 2838 1848 2841 1858
rect 2982 1857 2986 1858
rect 3014 1848 3017 1858
rect 3150 1848 3169 1851
rect 3774 1848 3777 1858
rect 3862 1848 3865 1858
rect 4782 1848 4785 1858
rect 4838 1848 4849 1851
rect 1235 1838 1238 1842
rect 1507 1838 1510 1842
rect 1818 1838 1821 1842
rect 2534 1838 2542 1841
rect 3563 1838 3566 1842
rect 4613 1838 4614 1842
rect 4770 1838 4771 1842
rect 1338 1818 1339 1822
rect 2405 1818 2406 1822
rect 4642 1818 4643 1822
rect 328 1803 330 1807
rect 334 1803 337 1807
rect 341 1803 344 1807
rect 1352 1803 1354 1807
rect 1358 1803 1361 1807
rect 1365 1803 1368 1807
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2397 1803 2400 1807
rect 3400 1803 3402 1807
rect 3406 1803 3409 1807
rect 3413 1803 3416 1807
rect 4424 1803 4426 1807
rect 4430 1803 4433 1807
rect 4437 1803 4440 1807
rect 434 1788 435 1792
rect 1541 1788 1542 1792
rect 1994 1788 1995 1792
rect 2026 1788 2027 1792
rect 2506 1788 2507 1792
rect 3506 1788 3507 1792
rect 3914 1788 3915 1792
rect 4682 1788 4683 1792
rect 2165 1778 2166 1782
rect 4277 1778 4278 1782
rect 1894 1768 1922 1771
rect 2765 1768 2766 1772
rect 4594 1768 4597 1772
rect 182 1748 190 1751
rect 446 1751 449 1761
rect 586 1758 590 1762
rect 446 1748 465 1751
rect 374 1741 377 1748
rect 638 1748 654 1751
rect 934 1748 961 1751
rect 1102 1751 1105 1761
rect 1338 1758 1342 1762
rect 1102 1748 1121 1751
rect 1350 1751 1353 1761
rect 1558 1752 1561 1761
rect 2058 1758 2062 1762
rect 2742 1758 2753 1761
rect 2742 1756 2746 1758
rect 1350 1748 1385 1751
rect 1390 1748 1398 1751
rect 1482 1748 1489 1751
rect 1646 1751 1650 1752
rect 1646 1748 1665 1751
rect 1758 1748 1777 1751
rect 366 1738 377 1741
rect 390 1738 398 1741
rect 470 1738 482 1741
rect 758 1738 777 1741
rect 790 1738 806 1741
rect 1414 1738 1425 1741
rect 1614 1738 1622 1741
rect 1774 1738 1777 1748
rect 1914 1748 1929 1751
rect 2050 1748 2057 1751
rect 2346 1748 2353 1751
rect 2998 1751 3001 1761
rect 3182 1758 3190 1761
rect 2998 1748 3017 1751
rect 3242 1748 3257 1751
rect 3318 1751 3321 1761
rect 3318 1748 3337 1751
rect 3522 1748 3537 1751
rect 3542 1742 3545 1751
rect 3582 1748 3601 1751
rect 3742 1748 3750 1751
rect 3814 1748 3830 1751
rect 3886 1748 3894 1751
rect 4054 1748 4062 1751
rect 4126 1748 4145 1751
rect 4262 1751 4265 1761
rect 4734 1752 4738 1753
rect 4246 1748 4265 1751
rect 4350 1748 4377 1751
rect 2174 1738 2193 1741
rect 2394 1738 2402 1741
rect 2606 1738 2625 1741
rect 3074 1738 3081 1741
rect 3086 1738 3094 1741
rect 3486 1738 3497 1741
rect 3582 1738 3590 1741
rect 3598 1738 3606 1741
rect 3702 1738 3714 1741
rect 3938 1738 3953 1741
rect 4198 1741 4201 1748
rect 4546 1748 4561 1751
rect 4618 1748 4633 1751
rect 4698 1748 4705 1751
rect 4854 1751 4857 1761
rect 4838 1748 4857 1751
rect 5102 1748 5121 1751
rect 5178 1748 5193 1751
rect 4190 1738 4201 1741
rect 4318 1738 4329 1741
rect 4410 1738 4418 1741
rect 4613 1738 4614 1742
rect 4990 1738 5001 1741
rect 478 1736 482 1738
rect 222 1731 226 1736
rect 210 1728 226 1731
rect 694 1731 698 1733
rect 346 1728 361 1731
rect 694 1728 705 1731
rect 742 1728 750 1731
rect 774 1728 777 1738
rect 1198 1728 1217 1731
rect 1222 1728 1225 1738
rect 1422 1732 1425 1738
rect 2174 1732 2177 1738
rect 2742 1732 2746 1733
rect 3198 1731 3202 1733
rect 3190 1728 3202 1731
rect 3614 1731 3618 1733
rect 3606 1728 3618 1731
rect 3798 1731 3802 1733
rect 3798 1728 3809 1731
rect 4110 1731 4114 1733
rect 4118 1731 4121 1738
rect 4110 1728 4121 1731
rect 4486 1731 4490 1736
rect 4574 1731 4578 1733
rect 4474 1728 4490 1731
rect 4566 1728 4578 1731
rect 4998 1732 5001 1738
rect 5006 1728 5025 1731
rect 5134 1731 5138 1733
rect 5130 1728 5138 1731
rect 381 1718 382 1722
rect 410 1718 411 1722
rect 1701 1718 1702 1722
rect 2610 1718 2611 1722
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 861 1703 864 1707
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1885 1703 1888 1707
rect 2888 1703 2890 1707
rect 2894 1703 2897 1707
rect 2901 1703 2904 1707
rect 3920 1703 3922 1707
rect 3926 1703 3929 1707
rect 3933 1703 3936 1707
rect 4936 1703 4938 1707
rect 4942 1703 4945 1707
rect 4949 1703 4952 1707
rect 318 1688 334 1691
rect 1862 1688 1873 1691
rect 3106 1688 3107 1692
rect 4274 1688 4275 1692
rect 366 1678 385 1681
rect 1246 1678 1254 1681
rect 1442 1678 1449 1681
rect 1454 1678 1473 1681
rect 1510 1678 1522 1681
rect 1870 1681 1873 1688
rect 1870 1678 1889 1681
rect 1998 1678 2009 1681
rect 1246 1677 1250 1678
rect 338 1668 353 1671
rect 562 1668 569 1671
rect 806 1668 814 1671
rect 886 1668 894 1671
rect 38 1658 46 1661
rect 190 1658 209 1661
rect 402 1658 409 1661
rect 638 1658 646 1661
rect 774 1658 793 1661
rect 802 1658 825 1661
rect 830 1658 865 1661
rect 1110 1662 1113 1671
rect 1134 1668 1142 1671
rect 1262 1668 1270 1671
rect 1422 1671 1425 1678
rect 1518 1677 1522 1678
rect 1422 1668 1433 1671
rect 1734 1668 1745 1671
rect 2126 1671 2129 1681
rect 2590 1678 2601 1681
rect 2670 1678 2689 1681
rect 2762 1678 2778 1681
rect 2590 1677 2594 1678
rect 2774 1674 2778 1678
rect 2790 1678 2801 1681
rect 2958 1678 2974 1681
rect 2790 1677 2794 1678
rect 2958 1674 2962 1678
rect 2118 1668 2129 1671
rect 2598 1668 2609 1671
rect 2802 1668 2809 1671
rect 2886 1668 2913 1671
rect 3062 1671 3065 1681
rect 3254 1678 3270 1681
rect 3342 1678 3361 1681
rect 3494 1678 3506 1681
rect 3806 1678 3817 1681
rect 3254 1674 3258 1678
rect 3502 1677 3506 1678
rect 3806 1677 3810 1678
rect 3062 1668 3081 1671
rect 3174 1668 3185 1671
rect 3210 1668 3217 1671
rect 3414 1668 3422 1671
rect 3470 1668 3478 1671
rect 3982 1671 3986 1674
rect 3834 1668 3841 1671
rect 3982 1668 3993 1671
rect 4134 1671 4138 1674
rect 4134 1668 4145 1671
rect 4214 1668 4222 1671
rect 4310 1671 4313 1681
rect 4358 1678 4374 1681
rect 4542 1678 4554 1681
rect 4358 1674 4362 1678
rect 4550 1677 4554 1678
rect 4294 1668 4313 1671
rect 4670 1671 4673 1681
rect 4782 1672 4786 1674
rect 4654 1668 4673 1671
rect 4678 1668 4686 1671
rect 4918 1671 4921 1678
rect 4998 1674 5002 1678
rect 4918 1668 4930 1671
rect 1378 1658 1401 1661
rect 1510 1661 1513 1668
rect 1502 1658 1513 1661
rect 2126 1662 2129 1668
rect 1654 1658 1662 1661
rect 1978 1658 1985 1661
rect 2110 1658 2118 1661
rect 2262 1658 2270 1661
rect 2298 1658 2305 1661
rect 2458 1658 2465 1661
rect 2598 1662 2601 1668
rect 2926 1658 2946 1661
rect 3418 1658 3441 1661
rect 3470 1658 3489 1661
rect 3686 1658 3694 1661
rect 3702 1658 3710 1661
rect 3822 1658 3841 1661
rect 3926 1658 3934 1661
rect 3998 1658 4017 1661
rect 4078 1658 4094 1661
rect 4150 1658 4169 1661
rect 4254 1658 4257 1668
rect 4518 1658 4526 1661
rect 4530 1658 4537 1661
rect 4594 1658 4609 1661
rect 4734 1658 4753 1661
rect 4826 1658 4841 1661
rect 4882 1658 4889 1661
rect 4958 1658 4974 1661
rect 5038 1658 5057 1661
rect 5082 1658 5090 1661
rect 5130 1658 5145 1661
rect 5238 1658 5249 1661
rect 190 1648 193 1658
rect 774 1648 777 1658
rect 862 1648 865 1658
rect 2942 1657 2946 1658
rect 1706 1648 1710 1652
rect 1890 1648 1897 1651
rect 2906 1648 2913 1651
rect 4014 1648 4017 1658
rect 4166 1648 4169 1658
rect 4750 1648 4753 1658
rect 5054 1648 5057 1658
rect 5086 1657 5090 1658
rect 5238 1652 5241 1658
rect 723 1638 726 1642
rect 1843 1638 1846 1642
rect 2109 1638 2110 1642
rect 2571 1638 2574 1642
rect 2962 1638 2965 1642
rect 3963 1638 3966 1642
rect 762 1628 763 1632
rect 2626 1628 2627 1632
rect 410 1618 411 1622
rect 637 1618 638 1622
rect 1346 1618 1347 1622
rect 4469 1618 4470 1622
rect 328 1603 330 1607
rect 334 1603 337 1607
rect 341 1603 344 1607
rect 1352 1603 1354 1607
rect 1358 1603 1361 1607
rect 1365 1603 1368 1607
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2397 1603 2400 1607
rect 3400 1603 3402 1607
rect 3406 1603 3409 1607
rect 3413 1603 3416 1607
rect 4424 1603 4426 1607
rect 4430 1603 4433 1607
rect 4437 1603 4440 1607
rect 226 1588 227 1592
rect 437 1588 438 1592
rect 626 1588 627 1592
rect 1101 1588 1102 1592
rect 1405 1588 1406 1592
rect 1445 1588 1446 1592
rect 2010 1588 2011 1592
rect 3338 1588 3339 1592
rect 3669 1588 3670 1592
rect 3858 1588 3859 1592
rect 4130 1588 4131 1592
rect 4189 1588 4190 1592
rect 4290 1588 4291 1592
rect 4338 1588 4339 1592
rect 2382 1578 2390 1581
rect 939 1568 942 1572
rect 1165 1568 1166 1572
rect 1718 1568 1729 1571
rect 4405 1568 4406 1572
rect 4930 1568 4937 1571
rect 1718 1562 1721 1568
rect 258 1558 262 1562
rect 1314 1558 1321 1561
rect 138 1548 145 1551
rect 302 1548 310 1551
rect 318 1548 326 1551
rect 346 1548 353 1551
rect 742 1548 758 1551
rect 990 1542 993 1551
rect 1558 1551 1561 1561
rect 1570 1558 1574 1562
rect 1786 1558 1790 1562
rect 1542 1548 1561 1551
rect 1710 1548 1718 1551
rect 1970 1548 1977 1551
rect 1982 1548 2009 1551
rect 282 1538 289 1541
rect 330 1538 353 1541
rect 1006 1538 1014 1541
rect 1070 1538 1078 1541
rect 1198 1538 1206 1541
rect 1326 1541 1329 1548
rect 1326 1538 1337 1541
rect 1766 1538 1769 1548
rect 1938 1538 1945 1541
rect 2030 1541 2033 1548
rect 2194 1548 2201 1551
rect 2258 1548 2265 1551
rect 2326 1548 2334 1551
rect 2454 1551 2457 1561
rect 2454 1548 2473 1551
rect 2478 1548 2486 1551
rect 2518 1551 2521 1561
rect 2502 1548 2521 1551
rect 2574 1551 2577 1561
rect 2678 1553 2682 1558
rect 2558 1548 2577 1551
rect 3022 1548 3033 1551
rect 3078 1551 3081 1561
rect 3350 1558 3369 1561
rect 4830 1552 4833 1561
rect 3050 1548 3057 1551
rect 3062 1548 3081 1551
rect 3154 1548 3169 1551
rect 3670 1548 3686 1551
rect 3966 1548 3982 1551
rect 4038 1548 4057 1551
rect 4134 1548 4142 1551
rect 4418 1548 4449 1551
rect 4454 1548 4462 1551
rect 4486 1548 4494 1551
rect 4518 1548 4526 1551
rect 4554 1548 4561 1551
rect 4666 1548 4673 1551
rect 2030 1538 2041 1541
rect 2290 1538 2298 1541
rect 2486 1538 2494 1541
rect 2906 1538 2913 1541
rect 3318 1538 3329 1541
rect 3526 1541 3529 1548
rect 3518 1538 3529 1541
rect 3614 1538 3625 1541
rect 4138 1538 4145 1541
rect 4166 1538 4169 1548
rect 4906 1548 4926 1551
rect 4978 1548 4993 1551
rect 5146 1548 5153 1551
rect 4262 1538 4281 1541
rect 4634 1538 4641 1541
rect 5078 1538 5086 1541
rect 798 1531 802 1533
rect 958 1531 962 1533
rect 1302 1531 1306 1533
rect 2790 1532 2794 1533
rect 798 1528 809 1531
rect 958 1528 969 1531
rect 974 1528 993 1531
rect 1302 1528 1313 1531
rect 3278 1528 3297 1531
rect 3574 1531 3577 1538
rect 3566 1528 3577 1531
rect 4022 1531 4026 1533
rect 4222 1532 4225 1538
rect 3694 1528 3713 1531
rect 4022 1528 4033 1531
rect 4218 1528 4225 1532
rect 1509 1518 1510 1522
rect 1925 1518 1926 1522
rect 2418 1518 2419 1522
rect 2525 1518 2526 1522
rect 4237 1518 4238 1522
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 861 1503 864 1507
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1885 1503 1888 1507
rect 2888 1503 2890 1507
rect 2894 1503 2897 1507
rect 2901 1503 2904 1507
rect 3920 1503 3922 1507
rect 3926 1503 3929 1507
rect 3933 1503 3936 1507
rect 4936 1503 4938 1507
rect 4942 1503 4945 1507
rect 4949 1503 4952 1507
rect 1997 1488 1998 1492
rect 166 1472 169 1481
rect 1022 1478 1033 1481
rect 1222 1478 1233 1481
rect 2534 1478 2553 1481
rect 2718 1478 2737 1481
rect 2998 1478 3009 1481
rect 1022 1477 1026 1478
rect 1222 1477 1226 1478
rect 2998 1472 3001 1478
rect 3262 1472 3266 1474
rect 190 1468 201 1471
rect 1038 1468 1049 1471
rect 1826 1468 1841 1471
rect 1866 1468 1881 1471
rect 1946 1468 1953 1471
rect 2354 1468 2362 1471
rect 2902 1468 2910 1471
rect 2982 1468 2990 1471
rect 3334 1471 3337 1481
rect 3502 1478 3521 1481
rect 3994 1478 4010 1481
rect 4006 1474 4010 1478
rect 4078 1478 4094 1481
rect 4486 1478 4498 1481
rect 4646 1478 4658 1481
rect 4078 1474 4082 1478
rect 4238 1474 4242 1478
rect 4494 1477 4498 1478
rect 4654 1477 4658 1478
rect 5222 1478 5238 1481
rect 3318 1468 3337 1471
rect 3350 1468 3366 1471
rect 3482 1468 3489 1471
rect 3806 1468 3814 1471
rect 3830 1468 3838 1471
rect 4822 1471 4825 1478
rect 5222 1474 5226 1478
rect 4822 1468 4833 1471
rect 5190 1468 5198 1471
rect 198 1462 201 1468
rect 1046 1462 1049 1468
rect 38 1458 46 1461
rect 326 1458 342 1461
rect 398 1458 417 1461
rect 798 1458 817 1461
rect 966 1458 974 1461
rect 1070 1458 1089 1461
rect 1278 1458 1286 1461
rect 1330 1458 1337 1461
rect 1410 1458 1417 1461
rect 1718 1458 1726 1461
rect 1750 1458 1769 1461
rect 1786 1458 1802 1461
rect 1902 1458 1910 1461
rect 1978 1458 1985 1461
rect 2026 1458 2033 1461
rect 2102 1458 2110 1461
rect 2242 1458 2257 1461
rect 2618 1458 2625 1461
rect 2834 1458 2841 1461
rect 2882 1458 2889 1461
rect 3054 1458 3062 1461
rect 3142 1458 3161 1461
rect 3214 1458 3230 1461
rect 3414 1458 3430 1461
rect 3566 1458 3582 1461
rect 3654 1458 3673 1461
rect 3730 1458 3745 1461
rect 3806 1458 3825 1461
rect 3858 1458 3862 1461
rect 3866 1458 3873 1461
rect 3886 1458 3905 1461
rect 4186 1458 4201 1461
rect 4326 1458 4345 1461
rect 4462 1458 4481 1461
rect 4622 1458 4641 1461
rect 4706 1458 4713 1461
rect 4894 1458 4913 1461
rect 4930 1458 4942 1461
rect 5250 1458 5265 1461
rect 170 1448 177 1451
rect 414 1448 417 1458
rect 1070 1448 1073 1458
rect 1234 1448 1241 1451
rect 1478 1448 1489 1451
rect 1750 1448 1753 1458
rect 2430 1452 2434 1457
rect 2098 1448 2102 1452
rect 2322 1448 2326 1452
rect 2870 1451 2874 1454
rect 2870 1448 2881 1451
rect 3142 1448 3145 1458
rect 3622 1452 3626 1454
rect 3654 1448 3657 1458
rect 3806 1448 3809 1458
rect 3886 1448 3889 1458
rect 4910 1448 4913 1458
rect 4922 1448 4926 1452
rect 1003 1438 1006 1442
rect 4003 1438 4006 1442
rect 4674 1438 4677 1442
rect 1338 1428 1339 1432
rect 4794 1428 4795 1432
rect 429 1418 430 1422
rect 458 1418 459 1422
rect 1429 1418 1430 1422
rect 328 1403 330 1407
rect 334 1403 337 1407
rect 341 1403 344 1407
rect 1352 1403 1354 1407
rect 1358 1403 1361 1407
rect 1365 1403 1368 1407
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2397 1403 2400 1407
rect 3400 1403 3402 1407
rect 3406 1403 3409 1407
rect 3413 1403 3416 1407
rect 4424 1403 4426 1407
rect 4430 1403 4433 1407
rect 4437 1403 4440 1407
rect 314 1388 321 1391
rect 1229 1388 1230 1392
rect 1354 1388 1369 1391
rect 1978 1388 1979 1392
rect 2034 1388 2035 1392
rect 2306 1388 2307 1392
rect 2354 1388 2355 1392
rect 3029 1388 3030 1392
rect 3962 1388 3969 1391
rect 4637 1388 4638 1392
rect 4701 1388 4702 1392
rect 4794 1388 4795 1392
rect 4450 1378 4457 1381
rect 4517 1378 4518 1382
rect 5066 1378 5067 1382
rect 770 1368 771 1372
rect 1037 1368 1038 1372
rect 2162 1368 2163 1372
rect 2194 1368 2195 1372
rect 2570 1368 2571 1372
rect 4842 1368 4845 1372
rect 4930 1368 4931 1372
rect 4954 1368 4970 1371
rect 1102 1366 1106 1368
rect 198 1351 201 1361
rect 294 1358 322 1361
rect 318 1356 322 1358
rect 198 1348 217 1351
rect 286 1348 310 1351
rect 550 1348 558 1351
rect 534 1338 537 1348
rect 782 1351 785 1361
rect 910 1353 914 1358
rect 782 1348 801 1351
rect 1038 1348 1046 1351
rect 1162 1348 1169 1351
rect 1202 1348 1217 1351
rect 1310 1351 1313 1361
rect 1618 1358 1622 1362
rect 1990 1358 2009 1361
rect 2410 1358 2414 1362
rect 2506 1358 2510 1362
rect 3162 1358 3166 1362
rect 3306 1358 3310 1362
rect 3454 1361 3457 1368
rect 3454 1358 3466 1361
rect 3594 1358 3601 1361
rect 3462 1356 3466 1358
rect 1278 1348 1297 1351
rect 1310 1348 1329 1351
rect 814 1338 830 1341
rect 962 1338 969 1341
rect 1278 1341 1281 1348
rect 1182 1338 1193 1341
rect 1270 1338 1281 1341
rect 1342 1338 1358 1341
rect 1598 1338 1601 1348
rect 2086 1348 2094 1351
rect 2154 1348 2161 1351
rect 2242 1348 2249 1351
rect 2366 1348 2398 1351
rect 2466 1348 2473 1351
rect 2490 1348 2505 1351
rect 2522 1348 2537 1351
rect 2654 1348 2662 1351
rect 2674 1348 2681 1351
rect 1666 1338 1673 1341
rect 2018 1338 2025 1341
rect 2278 1338 2297 1341
rect 2838 1338 2850 1341
rect 3142 1338 3145 1348
rect 3298 1348 3305 1351
rect 3506 1348 3521 1351
rect 3726 1348 3734 1351
rect 3998 1348 4006 1351
rect 4018 1348 4025 1351
rect 4310 1348 4329 1351
rect 4374 1348 4382 1351
rect 4394 1348 4401 1351
rect 4602 1348 4609 1351
rect 3286 1338 3297 1341
rect 3454 1338 3466 1341
rect 3574 1338 3601 1341
rect 3610 1338 3617 1341
rect 3782 1338 3790 1341
rect 3942 1338 3958 1341
rect 4094 1338 4102 1341
rect 4214 1338 4233 1341
rect 4734 1341 4737 1348
rect 4942 1351 4945 1361
rect 4942 1348 4977 1351
rect 4982 1348 4990 1351
rect 5014 1348 5030 1351
rect 5182 1351 5185 1361
rect 5302 1356 5306 1358
rect 5142 1348 5161 1351
rect 5166 1348 5185 1351
rect 4710 1338 4729 1341
rect 4734 1338 4745 1341
rect 5142 1341 5145 1348
rect 5134 1338 5145 1341
rect 3462 1336 3466 1338
rect 926 1331 930 1333
rect 926 1328 937 1331
rect 942 1328 961 1331
rect 1550 1331 1554 1333
rect 1550 1328 1561 1331
rect 1846 1328 1862 1331
rect 2918 1331 2922 1336
rect 2906 1328 2922 1331
rect 3434 1328 3446 1331
rect 3706 1328 3713 1331
rect 3718 1328 3726 1331
rect 4198 1331 4202 1333
rect 4198 1328 4209 1331
rect 4342 1331 4346 1333
rect 4334 1328 4346 1331
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 861 1303 864 1307
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1885 1303 1888 1307
rect 2888 1303 2890 1307
rect 2894 1303 2897 1307
rect 2901 1303 2904 1307
rect 3920 1303 3922 1307
rect 3926 1303 3929 1307
rect 3933 1303 3936 1307
rect 4936 1303 4938 1307
rect 4942 1303 4945 1307
rect 4949 1303 4952 1307
rect 310 1288 321 1291
rect 2765 1288 2766 1292
rect 3234 1288 3235 1292
rect 310 1281 313 1288
rect 294 1278 313 1281
rect 630 1278 641 1281
rect 774 1278 793 1281
rect 1850 1278 1857 1281
rect 1938 1278 1945 1282
rect 2414 1278 2433 1281
rect 2662 1278 2673 1281
rect 3110 1278 3122 1281
rect 418 1268 425 1271
rect 534 1268 546 1271
rect 598 1268 601 1278
rect 630 1277 634 1278
rect 1942 1272 1945 1278
rect 2662 1277 2666 1278
rect 3118 1277 3122 1278
rect 2646 1272 2650 1277
rect 822 1268 833 1271
rect 138 1258 145 1261
rect 206 1261 209 1268
rect 822 1262 825 1268
rect 950 1262 953 1271
rect 1438 1268 1457 1271
rect 1918 1268 1926 1271
rect 2502 1268 2513 1271
rect 2678 1268 2689 1271
rect 2710 1268 2718 1271
rect 2854 1268 2862 1271
rect 3086 1268 3094 1271
rect 3258 1268 3273 1271
rect 3310 1271 3313 1281
rect 3430 1278 3457 1281
rect 4230 1278 4241 1281
rect 4862 1278 4881 1281
rect 3430 1277 3434 1278
rect 4230 1277 4234 1278
rect 3310 1268 3329 1271
rect 3734 1268 3742 1271
rect 162 1258 169 1261
rect 198 1258 209 1261
rect 230 1258 238 1261
rect 286 1258 294 1261
rect 478 1258 486 1261
rect 686 1258 702 1261
rect 1062 1258 1081 1261
rect 1326 1258 1345 1261
rect 1398 1261 1401 1268
rect 1362 1258 1385 1261
rect 1390 1258 1401 1261
rect 1670 1258 1689 1261
rect 1998 1258 2006 1261
rect 2262 1258 2281 1261
rect 2458 1258 2473 1261
rect 2546 1258 2553 1261
rect 2710 1258 2729 1261
rect 2746 1258 2753 1261
rect 2926 1258 2945 1261
rect 3758 1262 3761 1271
rect 4106 1268 4121 1271
rect 4258 1268 4265 1271
rect 4882 1268 4889 1271
rect 3374 1258 3382 1261
rect 3462 1258 3481 1261
rect 3646 1258 3662 1261
rect 3734 1258 3753 1261
rect 3854 1258 3873 1261
rect 4038 1258 4049 1261
rect 4246 1258 4262 1261
rect 4318 1258 4326 1261
rect 5062 1258 5081 1261
rect 5154 1258 5169 1261
rect 5238 1258 5246 1261
rect 1078 1248 1081 1258
rect 1326 1248 1329 1258
rect 1686 1248 1689 1258
rect 2250 1248 2254 1252
rect 2262 1248 2265 1258
rect 2710 1248 2713 1258
rect 2942 1248 2945 1258
rect 3046 1252 3050 1257
rect 3734 1248 3737 1258
rect 3854 1248 3857 1258
rect 4038 1257 4042 1258
rect 4022 1252 4026 1257
rect 5078 1248 5081 1258
rect 5222 1252 5226 1257
rect 1022 1242 1026 1244
rect 173 1238 174 1242
rect 723 1238 726 1242
rect 2026 1238 2027 1242
rect 4970 1238 4973 1242
rect 3909 1218 3910 1222
rect 328 1203 330 1207
rect 334 1203 337 1207
rect 341 1203 344 1207
rect 1352 1203 1354 1207
rect 1358 1203 1361 1207
rect 1365 1203 1368 1207
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2397 1203 2400 1207
rect 3400 1203 3402 1207
rect 3406 1203 3409 1207
rect 3413 1203 3416 1207
rect 4424 1203 4426 1207
rect 4430 1203 4433 1207
rect 4437 1203 4440 1207
rect 642 1188 643 1192
rect 805 1188 806 1192
rect 842 1188 843 1192
rect 1013 1188 1014 1192
rect 1386 1188 1387 1192
rect 1506 1188 1507 1192
rect 2125 1188 2126 1192
rect 2570 1188 2571 1192
rect 3034 1188 3035 1192
rect 3549 1188 3550 1192
rect 4149 1188 4150 1192
rect 4333 1188 4334 1192
rect 4725 1188 4726 1192
rect 3125 1178 3126 1182
rect 4637 1178 4638 1182
rect 149 1168 150 1172
rect 234 1168 235 1172
rect 922 1168 923 1172
rect 1195 1168 1198 1172
rect 1691 1168 1694 1172
rect 2722 1168 2729 1171
rect 4499 1168 4502 1172
rect 4518 1168 4526 1171
rect 4670 1168 4697 1171
rect 4885 1168 4886 1172
rect 4670 1162 4673 1168
rect 442 1158 446 1162
rect 562 1158 569 1161
rect 694 1158 713 1161
rect 934 1158 942 1161
rect 1262 1158 1281 1161
rect 1290 1158 1294 1162
rect 1450 1158 1454 1162
rect 2178 1158 2183 1162
rect 2458 1158 2462 1162
rect 94 1156 98 1158
rect 38 1148 46 1151
rect 106 1148 113 1151
rect 150 1148 158 1151
rect 218 1148 233 1151
rect 250 1148 257 1151
rect 394 1148 406 1151
rect 426 1148 441 1151
rect 494 1148 510 1151
rect 618 1148 625 1151
rect 722 1148 729 1151
rect 786 1148 793 1151
rect 1354 1148 1385 1151
rect 1518 1148 1526 1151
rect 1550 1148 1558 1151
rect 1778 1148 1785 1151
rect 1494 1146 1498 1148
rect 2058 1148 2065 1151
rect 2126 1148 2153 1151
rect 2190 1148 2206 1151
rect 2470 1151 2473 1161
rect 3426 1158 3433 1161
rect 3514 1158 3518 1162
rect 4538 1158 4542 1162
rect 5114 1158 5118 1162
rect 2470 1148 2489 1151
rect 2738 1148 2745 1151
rect 2922 1148 2929 1151
rect 3250 1148 3257 1151
rect 3282 1148 3289 1151
rect 3462 1148 3481 1151
rect 3662 1151 3666 1153
rect 3598 1148 3617 1151
rect 3646 1148 3666 1151
rect 3778 1148 3785 1151
rect 3914 1148 3921 1151
rect 4022 1148 4030 1151
rect 4082 1148 4097 1151
rect 722 1138 737 1141
rect 950 1138 961 1141
rect 1478 1138 1486 1141
rect 1526 1138 1545 1141
rect 1554 1138 1569 1141
rect 2526 1138 2534 1141
rect 2606 1138 2614 1141
rect 2738 1138 2745 1141
rect 2818 1138 2825 1141
rect 2918 1138 2937 1141
rect 3950 1138 3958 1141
rect 4326 1141 4329 1151
rect 4386 1148 4393 1151
rect 4462 1148 4470 1151
rect 4694 1148 4713 1151
rect 4898 1148 4913 1151
rect 5050 1148 5065 1151
rect 5258 1148 5273 1151
rect 4310 1138 4329 1141
rect 4558 1138 4561 1148
rect 4582 1138 4590 1141
rect 4813 1138 4814 1142
rect 4942 1138 4977 1141
rect 550 1131 554 1133
rect 550 1128 561 1131
rect 750 1128 769 1131
rect 1094 1128 1113 1131
rect 1710 1131 1714 1133
rect 1710 1128 1721 1131
rect 1966 1131 1970 1136
rect 2526 1132 2529 1138
rect 1954 1128 1970 1131
rect 2074 1128 2081 1131
rect 2294 1128 2305 1131
rect 2710 1131 2714 1133
rect 2710 1128 2721 1131
rect 2918 1131 2921 1138
rect 2914 1128 2921 1131
rect 2982 1128 2993 1131
rect 3862 1131 3866 1133
rect 4326 1132 4329 1138
rect 3854 1128 3866 1131
rect 4774 1131 4778 1133
rect 4766 1128 4778 1131
rect 4974 1128 4977 1138
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 861 1103 864 1107
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1885 1103 1888 1107
rect 2888 1103 2890 1107
rect 2894 1103 2897 1107
rect 2901 1103 2904 1107
rect 3920 1103 3922 1107
rect 3926 1103 3929 1107
rect 3933 1103 3936 1107
rect 4936 1103 4938 1107
rect 4942 1103 4945 1107
rect 4949 1103 4952 1107
rect 957 1088 958 1092
rect 981 1088 982 1092
rect 1878 1088 1894 1091
rect 4085 1088 4086 1092
rect 4138 1088 4139 1092
rect 94 1078 105 1081
rect 622 1078 641 1081
rect 1278 1078 1289 1081
rect 1322 1078 1323 1082
rect 62 1068 65 1078
rect 94 1077 98 1078
rect 1278 1077 1282 1078
rect 122 1068 129 1071
rect 330 1068 345 1071
rect 1454 1068 1457 1078
rect 1566 1074 1570 1078
rect 1582 1078 1593 1081
rect 1598 1078 1617 1081
rect 1926 1078 1945 1081
rect 1982 1078 2001 1081
rect 3626 1078 3633 1081
rect 1582 1077 1586 1078
rect 1618 1068 1625 1071
rect 1742 1068 1750 1071
rect 2102 1071 2106 1074
rect 2102 1068 2113 1071
rect 2214 1068 2222 1071
rect 2538 1068 2545 1071
rect 3014 1068 3022 1071
rect 3358 1068 3377 1071
rect 3506 1068 3513 1071
rect 3558 1068 3569 1071
rect 3598 1068 3617 1071
rect 3722 1068 3737 1071
rect 3922 1068 3945 1071
rect 3966 1068 3974 1071
rect 4030 1071 4033 1081
rect 4286 1078 4302 1081
rect 4854 1078 4873 1081
rect 4286 1074 4290 1078
rect 4014 1068 4033 1071
rect 110 1058 118 1061
rect 278 1058 294 1061
rect 338 1058 353 1061
rect 650 1058 657 1061
rect 886 1058 902 1061
rect 1070 1061 1073 1068
rect 1070 1058 1081 1061
rect 1638 1058 1646 1061
rect 1670 1058 1678 1061
rect 2350 1058 2369 1061
rect 2678 1058 2697 1061
rect 2742 1058 2761 1061
rect 2842 1058 2849 1061
rect 3014 1058 3033 1061
rect 3262 1058 3281 1061
rect 3306 1058 3313 1061
rect 3318 1058 3337 1061
rect 3710 1058 3718 1061
rect 3910 1058 3945 1061
rect 4058 1058 4073 1061
rect 4110 1058 4118 1061
rect 4210 1058 4217 1061
rect 4262 1058 4274 1061
rect 4374 1058 4393 1061
rect 4470 1058 4486 1061
rect 4542 1058 4550 1061
rect 4582 1058 4601 1061
rect 4702 1058 4721 1061
rect 5250 1058 5265 1061
rect 1290 1048 1297 1051
rect 2114 1048 2121 1051
rect 2350 1048 2353 1058
rect 2694 1048 2697 1058
rect 2758 1048 2761 1058
rect 3262 1048 3265 1058
rect 3334 1048 3337 1058
rect 3942 1048 3945 1058
rect 4270 1057 4274 1058
rect 4390 1048 4393 1058
rect 4582 1048 4585 1058
rect 4718 1048 4721 1058
rect 950 1042 954 1044
rect 694 1038 702 1041
rect 966 1041 969 1048
rect 974 1041 978 1044
rect 966 1038 978 1041
rect 1259 1038 1262 1042
rect 1563 1038 1566 1042
rect 306 1018 307 1022
rect 2957 1018 2958 1022
rect 328 1003 330 1007
rect 334 1003 337 1007
rect 341 1003 344 1007
rect 1352 1003 1354 1007
rect 1358 1003 1361 1007
rect 1365 1003 1368 1007
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2397 1003 2400 1007
rect 3400 1003 3402 1007
rect 3406 1003 3409 1007
rect 3413 1003 3416 1007
rect 4424 1003 4426 1007
rect 4430 1003 4433 1007
rect 4437 1003 4440 1007
rect 226 988 227 992
rect 453 988 454 992
rect 818 988 819 992
rect 1653 988 1654 992
rect 1685 988 1686 992
rect 2754 988 2755 992
rect 2810 988 2811 992
rect 3450 988 3451 992
rect 4170 988 4171 992
rect 4405 988 4406 992
rect 197 978 198 982
rect 690 968 691 972
rect 957 968 958 972
rect 2037 968 2038 972
rect 2586 968 2593 971
rect 2722 968 2723 972
rect 2946 968 2949 972
rect 3858 968 3861 972
rect 114 958 118 962
rect 126 951 129 961
rect 326 958 334 961
rect 126 948 145 951
rect 282 948 289 951
rect 390 948 398 951
rect 830 951 833 961
rect 830 948 849 951
rect 1070 951 1073 961
rect 1070 948 1089 951
rect 1134 951 1137 961
rect 1134 948 1153 951
rect 1246 951 1249 961
rect 1230 948 1249 951
rect 1322 948 1337 951
rect 1810 948 1817 951
rect 1902 948 1910 951
rect 2202 948 2209 951
rect 2246 948 2257 951
rect 2650 948 2657 951
rect 2822 951 2825 961
rect 3174 961 3177 968
rect 2922 958 2930 961
rect 3166 958 3177 961
rect 2926 956 2930 958
rect 2822 948 2841 951
rect 2902 948 2910 951
rect 2970 948 2985 951
rect 3158 948 3169 951
rect 530 938 531 942
rect 670 938 681 941
rect 854 938 870 941
rect 930 938 937 941
rect 1378 938 1401 941
rect 1478 941 1481 948
rect 2246 942 2249 948
rect 1470 938 1481 941
rect 1710 938 1729 941
rect 1846 938 1874 941
rect 1990 938 2009 941
rect 2274 938 2281 941
rect 2446 938 2454 941
rect 2598 941 2601 948
rect 3514 948 3521 951
rect 3750 951 3753 961
rect 4226 958 4233 961
rect 3750 948 3769 951
rect 3778 948 3793 951
rect 3890 948 3897 951
rect 4174 948 4182 951
rect 4190 948 4198 951
rect 4338 948 4353 951
rect 4414 948 4449 951
rect 2598 938 2609 941
rect 2794 938 2801 941
rect 2846 938 2854 941
rect 3282 938 3289 941
rect 3478 938 3486 941
rect 4142 938 4161 941
rect 4262 938 4265 948
rect 4414 938 4417 948
rect 4694 948 4702 951
rect 4774 948 4782 951
rect 4822 948 4830 951
rect 5010 948 5017 951
rect 5202 948 5209 951
rect 4782 938 4793 941
rect 4894 938 4913 941
rect 598 928 617 931
rect 782 931 786 936
rect 770 928 786 931
rect 901 928 902 932
rect 1446 928 1465 931
rect 1470 928 1473 938
rect 1694 928 1702 931
rect 1726 928 1729 938
rect 1990 928 1993 938
rect 2150 931 2154 933
rect 2142 928 2154 931
rect 2454 928 2473 931
rect 2574 931 2578 933
rect 2574 928 2585 931
rect 2670 928 2681 931
rect 2854 928 2857 938
rect 2862 928 2881 931
rect 3038 931 3042 933
rect 3030 928 3042 931
rect 3182 931 3186 933
rect 3438 931 3441 938
rect 3174 928 3186 931
rect 3422 928 3441 931
rect 3486 928 3505 931
rect 3582 928 3601 931
rect 4102 928 4121 931
rect 4126 928 4134 931
rect 4158 928 4161 938
rect 4302 936 4306 938
rect 4590 932 4594 936
rect 4502 928 4510 931
rect 4910 928 4913 938
rect 4958 931 4962 933
rect 4954 928 4962 931
rect 3422 921 3425 928
rect 3414 918 3425 921
rect 848 903 850 907
rect 854 903 857 907
rect 861 903 864 907
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1885 903 1888 907
rect 2888 903 2890 907
rect 2894 903 2897 907
rect 2901 903 2904 907
rect 3920 903 3922 907
rect 3926 903 3929 907
rect 3933 903 3936 907
rect 4936 903 4938 907
rect 4942 903 4945 907
rect 4949 903 4952 907
rect 933 888 934 892
rect 1382 888 1393 891
rect 2378 888 2393 891
rect 2765 888 2766 892
rect 4242 888 4243 892
rect 126 878 145 881
rect 694 878 713 881
rect 1390 881 1393 888
rect 1390 878 1406 881
rect 382 874 386 878
rect 586 868 593 871
rect 1426 868 1433 871
rect 1654 871 1657 881
rect 1922 878 1937 881
rect 1942 878 1961 881
rect 2622 878 2633 881
rect 2678 878 2694 881
rect 2678 874 2682 878
rect 1638 868 1657 871
rect 1750 868 1761 871
rect 1910 868 1926 871
rect 2134 868 2153 871
rect 2346 868 2353 871
rect 2546 868 2561 871
rect 2782 871 2785 881
rect 2790 878 2809 881
rect 3238 878 3249 881
rect 3382 878 3401 881
rect 3238 877 3242 878
rect 2778 868 2785 871
rect 286 858 302 861
rect 622 858 641 861
rect 826 858 833 861
rect 846 858 881 861
rect 1070 858 1089 861
rect 1222 858 1241 861
rect 1414 858 1433 861
rect 1690 858 1697 861
rect 1774 858 1793 861
rect 1958 858 1961 868
rect 2198 858 2206 861
rect 2366 858 2374 861
rect 2542 858 2550 861
rect 2714 858 2721 861
rect 2918 858 2934 861
rect 3006 861 3009 871
rect 3498 868 3505 871
rect 3742 868 3761 871
rect 3822 871 3825 881
rect 4310 878 4329 881
rect 4518 878 4537 881
rect 4542 878 4550 881
rect 4710 878 4729 881
rect 3822 868 3841 871
rect 4037 868 4038 872
rect 4114 868 4121 871
rect 4294 868 4302 871
rect 4546 868 4561 871
rect 4566 868 4585 871
rect 5070 871 5073 881
rect 5126 878 5145 881
rect 5222 878 5238 881
rect 5222 874 5226 878
rect 5070 868 5089 871
rect 5094 868 5113 871
rect 5190 868 5198 871
rect 3006 858 3017 861
rect 3134 858 3142 861
rect 3294 858 3310 861
rect 3510 858 3529 861
rect 3534 858 3542 861
rect 3582 858 3590 861
rect 3770 858 3777 861
rect 3930 858 3945 861
rect 4102 858 4121 861
rect 4174 858 4193 861
rect 4350 858 4358 861
rect 4566 858 4569 868
rect 4682 858 4689 861
rect 5094 862 5097 868
rect 4942 858 4977 861
rect 5250 858 5265 861
rect 638 848 641 858
rect 846 848 849 858
rect 866 848 873 851
rect 1070 848 1073 858
rect 1238 848 1241 858
rect 3014 852 3017 858
rect 3350 857 3354 858
rect 2226 848 2230 852
rect 3774 848 3777 858
rect 3866 848 3870 852
rect 4190 848 4193 858
rect 4282 848 4286 852
rect 926 842 930 844
rect 323 838 326 842
rect 834 838 835 842
rect 1603 838 1606 842
rect 2491 838 2494 842
rect 3331 838 3334 842
rect 3789 838 3790 842
rect 909 828 910 832
rect 170 818 171 822
rect 342 818 350 821
rect 533 818 534 822
rect 653 818 654 822
rect 1058 818 1059 822
rect 1698 818 1699 822
rect 328 803 330 807
rect 334 803 337 807
rect 341 803 344 807
rect 1352 803 1354 807
rect 1358 803 1361 807
rect 1365 803 1368 807
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2397 803 2400 807
rect 3400 803 3402 807
rect 3406 803 3409 807
rect 3413 803 3416 807
rect 4424 803 4426 807
rect 4430 803 4433 807
rect 4437 803 4440 807
rect 749 788 750 792
rect 973 788 974 792
rect 1221 788 1222 792
rect 1245 788 1246 792
rect 1389 788 1390 792
rect 1837 788 1838 792
rect 2277 788 2278 792
rect 2357 788 2358 792
rect 2450 788 2451 792
rect 4965 788 4966 792
rect 1115 768 1118 772
rect 1890 768 1897 771
rect 2563 768 2566 772
rect 2877 768 2878 772
rect 3594 768 3597 772
rect 3694 768 3705 771
rect 4810 768 4811 772
rect 142 748 150 751
rect 210 748 217 751
rect 354 748 361 751
rect 398 748 414 751
rect 474 748 481 751
rect 570 748 577 751
rect 658 748 673 751
rect 974 748 982 751
rect 1014 751 1017 761
rect 1146 758 1153 761
rect 1014 748 1033 751
rect 1370 748 1377 751
rect 1446 748 1465 751
rect 1578 748 1585 751
rect 1750 751 1753 761
rect 2306 758 2310 762
rect 1734 748 1753 751
rect 1854 748 1865 751
rect 1870 748 1886 751
rect 1854 742 1857 748
rect 2074 748 2081 751
rect 2238 748 2249 751
rect 2290 748 2297 751
rect 2330 748 2337 751
rect 2358 748 2382 751
rect 2462 751 2465 761
rect 3094 761 3097 768
rect 3086 758 3097 761
rect 3442 758 3446 762
rect 2462 748 2481 751
rect 2526 748 2542 751
rect 2642 748 2649 751
rect 2246 742 2249 748
rect 10 738 17 741
rect 490 738 497 741
rect 1446 738 1454 741
rect 1774 738 1782 741
rect 2014 738 2033 741
rect 2062 738 2070 741
rect 2294 738 2297 748
rect 2774 748 2782 751
rect 2786 748 2793 751
rect 2878 748 2902 751
rect 3006 748 3033 751
rect 3454 751 3457 761
rect 3966 752 3969 761
rect 4050 758 4054 762
rect 4598 756 4602 758
rect 3454 748 3473 751
rect 3618 748 3633 751
rect 3686 748 3694 751
rect 4002 748 4009 751
rect 4054 748 4062 751
rect 4134 748 4153 751
rect 4242 748 4257 751
rect 4326 748 4334 751
rect 4434 748 4454 751
rect 2846 738 2854 741
rect 3406 738 3422 741
rect 3486 738 3494 741
rect 4006 738 4009 748
rect 4722 748 4737 751
rect 4782 748 4793 751
rect 5030 751 5033 761
rect 5030 748 5049 751
rect 5134 751 5137 761
rect 5146 758 5150 762
rect 5118 748 5137 751
rect 5150 748 5158 751
rect 4790 742 4793 748
rect 4134 738 4142 741
rect 4438 738 4446 741
rect 4974 738 4993 741
rect 5098 738 5105 741
rect 334 728 353 731
rect 438 728 457 731
rect 710 731 713 738
rect 1486 736 1490 738
rect 710 728 721 731
rect 790 728 809 731
rect 1242 728 1249 731
rect 1478 731 1482 733
rect 1470 728 1482 731
rect 2014 728 2017 738
rect 2102 728 2121 731
rect 2582 731 2586 733
rect 2582 728 2593 731
rect 2686 731 2690 736
rect 2686 728 2702 731
rect 3102 731 3106 733
rect 4510 732 4514 736
rect 3094 728 3106 731
rect 3526 728 3545 731
rect 4678 731 4682 733
rect 4670 728 4682 731
rect 334 721 337 728
rect 326 718 337 721
rect 386 718 387 722
rect 848 703 850 707
rect 854 703 857 707
rect 861 703 864 707
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1885 703 1888 707
rect 2888 703 2890 707
rect 2894 703 2897 707
rect 2901 703 2904 707
rect 3920 703 3922 707
rect 3926 703 3929 707
rect 3933 703 3936 707
rect 4936 703 4938 707
rect 4942 703 4945 707
rect 4949 703 4952 707
rect 738 688 739 692
rect 1181 688 1182 692
rect 3890 688 3897 691
rect 4442 688 4449 691
rect 4934 688 4942 691
rect 646 678 665 681
rect 1334 678 1345 681
rect 2102 678 2114 681
rect 1334 677 1338 678
rect 2110 677 2114 678
rect 142 668 153 671
rect 686 668 697 671
rect 1422 668 1441 671
rect 1830 668 1841 671
rect 1870 668 1897 671
rect 2142 668 2145 678
rect 2318 674 2322 678
rect 2606 672 2609 681
rect 2614 678 2633 681
rect 3158 678 3177 681
rect 2478 668 2497 671
rect 2634 668 2641 671
rect 54 658 62 661
rect 94 658 113 661
rect 122 658 129 661
rect 310 658 345 661
rect 450 658 457 661
rect 1018 658 1025 661
rect 1110 658 1118 661
rect 1406 658 1425 661
rect 1462 658 1481 661
rect 1550 658 1558 661
rect 1722 658 1729 661
rect 1894 661 1897 668
rect 1894 658 1910 661
rect 1918 658 1937 661
rect 2286 658 2294 661
rect 2710 662 2713 671
rect 2846 662 2849 671
rect 2894 668 2918 671
rect 3318 671 3321 681
rect 4078 678 4089 681
rect 4550 678 4569 681
rect 4838 678 4849 681
rect 3318 668 3337 671
rect 3538 668 3553 671
rect 3814 671 3818 674
rect 4086 672 4089 678
rect 4838 677 4842 678
rect 3814 668 3825 671
rect 2806 658 2822 661
rect 2914 658 2937 661
rect 3102 658 3110 661
rect 3122 658 3129 661
rect 3350 658 3358 661
rect 3410 658 3425 661
rect 3454 661 3457 668
rect 3454 658 3465 661
rect 3470 658 3478 661
rect 3698 658 3705 661
rect 3830 658 3849 661
rect 4046 658 4054 661
rect 4058 658 4065 661
rect 4158 658 4177 661
rect 4402 658 4409 661
rect 4498 658 4505 661
rect 4602 658 4609 661
rect 4622 661 4625 671
rect 4622 658 4630 661
rect 4734 658 4742 661
rect 4782 658 4790 661
rect 4854 658 4873 661
rect 5022 658 5041 661
rect 5122 658 5129 661
rect 5170 658 5177 661
rect 94 648 97 658
rect 342 648 345 658
rect 390 651 393 658
rect 382 648 393 651
rect 1462 648 1465 658
rect 1934 648 1937 658
rect 2806 657 2810 658
rect 2126 652 2130 657
rect 1946 648 1950 652
rect 2970 648 2974 652
rect 3078 651 3082 654
rect 3078 648 3089 651
rect 3098 648 3102 652
rect 3674 648 3678 652
rect 3846 648 3849 658
rect 4034 648 4038 652
rect 4046 648 4049 658
rect 4174 648 4177 658
rect 4934 648 4942 651
rect 5038 648 5041 658
rect 958 642 962 644
rect 274 638 275 642
rect 318 638 334 641
rect 1174 642 1178 644
rect 2221 638 2222 642
rect 4309 638 4310 642
rect 5190 638 5201 641
rect 29 618 30 622
rect 82 618 83 622
rect 242 618 243 622
rect 357 618 358 622
rect 1037 618 1038 622
rect 1786 618 1787 622
rect 2669 618 2670 622
rect 2938 618 2939 622
rect 3549 618 3550 622
rect 4002 618 4003 622
rect 4093 618 4094 622
rect 4189 618 4190 622
rect 4213 618 4214 622
rect 328 603 330 607
rect 334 603 337 607
rect 341 603 344 607
rect 1352 603 1354 607
rect 1358 603 1361 607
rect 1365 603 1368 607
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2397 603 2400 607
rect 3400 603 3402 607
rect 3406 603 3409 607
rect 3413 603 3416 607
rect 4424 603 4426 607
rect 4430 603 4433 607
rect 4437 603 4440 607
rect 498 588 499 592
rect 810 588 811 592
rect 914 588 915 592
rect 1282 588 1283 592
rect 1818 588 1819 592
rect 1842 588 1843 592
rect 2005 588 2006 592
rect 2037 588 2038 592
rect 2398 588 2406 591
rect 2493 588 2494 592
rect 3186 588 3187 592
rect 3522 588 3523 592
rect 3581 588 3582 592
rect 5106 588 5107 592
rect 1677 578 1678 582
rect 874 568 882 571
rect 878 566 882 568
rect 1610 568 1611 572
rect 2202 568 2205 572
rect 2398 568 2426 571
rect 2437 568 2438 572
rect 2906 568 2913 571
rect 4002 568 4003 572
rect 4226 568 4229 572
rect 5210 568 5217 571
rect 510 558 529 561
rect 894 561 897 568
rect 886 558 897 561
rect 302 548 310 551
rect 906 548 913 551
rect 1098 548 1113 551
rect 1318 548 1334 551
rect 1342 548 1366 551
rect 1526 551 1529 561
rect 1526 548 1545 551
rect 1626 548 1633 551
rect 1662 551 1665 561
rect 1854 558 1862 561
rect 1646 548 1665 551
rect 62 532 65 542
rect 314 538 321 541
rect 478 538 489 541
rect 1630 538 1633 548
rect 1798 548 1809 551
rect 2006 548 2022 551
rect 2150 551 2153 561
rect 2122 548 2129 551
rect 2134 548 2153 551
rect 2166 548 2174 551
rect 2282 548 2289 551
rect 1806 542 1809 548
rect 1950 538 1969 541
rect 2114 538 2121 541
rect 2302 538 2305 548
rect 2450 548 2457 551
rect 2494 548 2502 551
rect 2630 542 2633 551
rect 3046 551 3049 561
rect 3198 558 3209 561
rect 5118 558 5129 561
rect 3030 548 3049 551
rect 3538 548 3545 551
rect 3582 548 3590 551
rect 3726 551 3730 553
rect 3710 548 3730 551
rect 3830 548 3849 551
rect 4250 548 4265 551
rect 4346 548 4361 551
rect 4558 548 4566 551
rect 4810 548 4825 551
rect 5182 551 5185 561
rect 5162 548 5169 551
rect 5182 548 5201 551
rect 2782 538 2801 541
rect 2878 538 2894 541
rect 3042 538 3049 541
rect 3478 538 3497 541
rect 3678 538 3686 541
rect 3886 538 3889 548
rect 3910 538 3918 541
rect 4030 538 4041 541
rect 4534 538 4553 541
rect 286 531 290 533
rect 462 531 466 533
rect 286 528 297 531
rect 462 528 473 531
rect 766 531 770 533
rect 766 528 777 531
rect 942 528 961 531
rect 1174 531 1178 533
rect 1950 532 1953 538
rect 1154 528 1161 531
rect 1166 528 1178 531
rect 2606 528 2609 538
rect 2614 528 2633 531
rect 2782 528 2785 538
rect 2837 528 2838 532
rect 2926 531 2930 533
rect 2918 528 2930 531
rect 3478 528 3481 538
rect 3506 528 3513 531
rect 3822 528 3825 538
rect 3950 531 3953 538
rect 3942 528 3953 531
rect 4030 532 4033 538
rect 4158 528 4177 531
rect 4430 531 4434 536
rect 4430 528 4446 531
rect 4534 528 4537 538
rect 4622 531 4626 533
rect 4766 531 4770 533
rect 4614 528 4626 531
rect 4758 528 4770 531
rect 4798 532 4801 542
rect 5066 538 5073 541
rect 5078 538 5086 541
rect 5182 538 5190 541
rect 4950 528 4958 531
rect 848 503 850 507
rect 854 503 857 507
rect 861 503 864 507
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1885 503 1888 507
rect 2888 503 2890 507
rect 2894 503 2897 507
rect 2901 503 2904 507
rect 3920 503 3922 507
rect 3926 503 3929 507
rect 3933 503 3936 507
rect 4936 503 4938 507
rect 4942 503 4945 507
rect 4949 503 4952 507
rect 661 488 662 492
rect 765 488 766 492
rect 1261 488 1262 492
rect 2461 488 2462 492
rect 94 478 105 481
rect 94 477 98 478
rect 110 468 121 471
rect 334 471 337 481
rect 346 478 361 481
rect 510 478 529 481
rect 998 478 1010 481
rect 1126 478 1145 481
rect 1218 478 1234 481
rect 1538 478 1554 481
rect 1742 478 1750 481
rect 1006 477 1010 478
rect 1230 474 1234 478
rect 1550 474 1554 478
rect 1774 474 1778 478
rect 334 468 369 471
rect 706 468 721 471
rect 974 468 982 471
rect 118 462 121 468
rect 38 458 46 461
rect 158 458 166 461
rect 458 458 465 461
rect 778 458 793 461
rect 974 458 993 461
rect 1126 458 1129 468
rect 1278 461 1281 471
rect 1434 468 1435 472
rect 1878 471 1881 481
rect 1878 468 1913 471
rect 1922 468 1929 471
rect 2038 468 2049 471
rect 2070 468 2078 471
rect 2134 468 2145 471
rect 2378 468 2390 471
rect 2478 471 2482 474
rect 2670 472 2673 481
rect 2678 478 2697 481
rect 3518 478 3526 481
rect 3518 477 3522 478
rect 2470 468 2482 471
rect 2942 468 2958 471
rect 3222 468 3233 471
rect 3386 468 3393 471
rect 3546 468 3553 471
rect 3798 471 3801 481
rect 3794 468 3801 471
rect 3814 468 3841 471
rect 4014 471 4017 481
rect 4342 478 4361 481
rect 4254 472 4258 477
rect 3998 468 4017 471
rect 4146 468 4153 471
rect 4398 468 4417 471
rect 4458 468 4465 471
rect 4714 468 4721 471
rect 1274 458 1281 461
rect 1334 458 1353 461
rect 1510 458 1526 461
rect 1686 458 1713 461
rect 1718 458 1734 461
rect 1750 458 1762 461
rect 2002 458 2009 461
rect 2146 458 2153 461
rect 2302 458 2321 461
rect 2406 458 2414 461
rect 2694 458 2697 468
rect 2758 458 2766 461
rect 2942 461 2945 468
rect 2934 458 2945 461
rect 3046 458 3054 461
rect 3094 458 3102 461
rect 3182 458 3201 461
rect 3222 461 3225 468
rect 3210 458 3225 461
rect 3246 458 3254 461
rect 3406 458 3422 461
rect 3526 458 3529 468
rect 3574 458 3593 461
rect 3666 458 3673 461
rect 3714 458 3721 461
rect 3726 458 3745 461
rect 3846 458 3865 461
rect 3870 458 3889 461
rect 3894 458 3926 461
rect 3942 458 3961 461
rect 3974 458 3982 461
rect 4210 458 4217 461
rect 4222 458 4242 461
rect 4418 458 4425 461
rect 4478 458 4497 461
rect 4578 458 4585 461
rect 4734 458 4742 461
rect 5102 462 5105 471
rect 5118 468 5137 471
rect 4894 458 4913 461
rect 4982 458 4998 461
rect 5062 458 5078 461
rect 5138 458 5145 461
rect 1758 457 1762 458
rect 2302 448 2305 458
rect 2434 448 2438 452
rect 2834 448 2838 452
rect 2866 448 2870 452
rect 3182 448 3185 458
rect 3266 448 3270 452
rect 3362 448 3366 452
rect 3562 448 3566 452
rect 3574 448 3577 458
rect 3742 448 3745 458
rect 3958 448 3961 458
rect 4238 457 4242 458
rect 4494 448 4497 458
rect 4526 452 4530 454
rect 4790 452 4794 457
rect 4894 448 4897 458
rect 654 442 658 444
rect 758 442 762 444
rect 1227 438 1230 442
rect 1254 441 1258 444
rect 1246 438 1258 441
rect 3533 428 3534 432
rect 477 418 478 422
rect 805 418 806 422
rect 2357 418 2358 422
rect 3301 418 3302 422
rect 3330 418 3331 422
rect 3973 418 3974 422
rect 328 403 330 407
rect 334 403 337 407
rect 341 403 344 407
rect 1352 403 1354 407
rect 1358 403 1361 407
rect 1365 403 1368 407
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2397 403 2400 407
rect 3400 403 3402 407
rect 3406 403 3409 407
rect 3413 403 3416 407
rect 4424 403 4426 407
rect 4430 403 4433 407
rect 4437 403 4440 407
rect 933 388 934 392
rect 1565 388 1566 392
rect 3013 388 3014 392
rect 3642 388 3643 392
rect 3669 388 3670 392
rect 3730 388 3731 392
rect 3794 388 3795 392
rect 3826 388 3827 392
rect 3930 388 3945 391
rect 4541 388 4542 392
rect 4666 388 4667 392
rect 4962 388 4963 392
rect 5146 388 5147 392
rect 5181 388 5182 392
rect 5237 388 5238 392
rect 5293 388 5294 392
rect 3554 378 3555 382
rect 1366 368 1374 371
rect 3098 368 3101 372
rect 110 348 126 351
rect 258 348 273 351
rect 206 341 209 348
rect 206 338 218 341
rect 310 341 313 348
rect 310 338 321 341
rect 398 341 401 348
rect 686 348 702 351
rect 918 351 921 361
rect 902 348 921 351
rect 934 348 942 351
rect 958 348 977 351
rect 1190 348 1198 351
rect 1278 351 1281 361
rect 1354 358 1358 362
rect 1594 358 1598 362
rect 1262 348 1281 351
rect 1294 348 1318 351
rect 1326 348 1334 351
rect 1478 351 1482 353
rect 1346 348 1353 351
rect 1478 348 1497 351
rect 1522 348 1529 351
rect 1566 348 1582 351
rect 1646 351 1649 361
rect 1790 361 1793 368
rect 1782 358 1793 361
rect 3874 358 3878 362
rect 1630 348 1649 351
rect 1802 348 1809 351
rect 1814 348 1822 351
rect 1834 348 1841 351
rect 374 338 393 341
rect 398 338 417 341
rect 430 338 449 341
rect 1202 338 1209 341
rect 1854 338 1878 341
rect 1934 338 1937 348
rect 2142 348 2150 351
rect 2278 351 2282 353
rect 2262 348 2282 351
rect 2466 348 2473 351
rect 2762 348 2769 351
rect 3046 348 3054 351
rect 3178 348 3185 351
rect 3222 348 3230 351
rect 3582 348 3593 351
rect 3598 348 3606 351
rect 3786 348 3793 351
rect 3878 348 3894 351
rect 3986 348 4001 351
rect 3582 342 3585 348
rect 2454 338 2462 341
rect 2682 338 2689 341
rect 3422 338 3450 341
rect 3710 338 3713 348
rect 4158 351 4161 361
rect 4158 348 4177 351
rect 4230 348 4238 351
rect 4610 348 4617 351
rect 4946 348 4961 351
rect 5038 351 5042 353
rect 5034 348 5042 351
rect 5082 348 5097 351
rect 3778 338 3785 341
rect 3886 338 3905 341
rect 4366 338 4385 341
rect 4550 338 4562 341
rect 214 336 218 338
rect 166 331 170 333
rect 166 328 177 331
rect 374 328 377 338
rect 430 328 433 338
rect 782 331 786 333
rect 774 328 786 331
rect 1174 331 1178 333
rect 1174 328 1185 331
rect 2042 328 2049 331
rect 2102 328 2121 331
rect 2486 331 2490 333
rect 2478 328 2490 331
rect 2598 328 2601 338
rect 2606 328 2625 331
rect 2662 328 2681 331
rect 3078 331 3082 333
rect 3070 328 3082 331
rect 3197 328 3198 332
rect 3238 331 3242 333
rect 3230 328 3242 331
rect 3602 328 3609 331
rect 3614 328 3633 331
rect 3842 328 3849 331
rect 4382 328 4385 338
rect 4558 336 4562 338
rect 4566 336 4570 338
rect 4902 328 4921 331
rect 4926 328 4942 331
rect 5038 331 5042 333
rect 5006 328 5025 331
rect 5030 328 5042 331
rect 848 303 850 307
rect 854 303 857 307
rect 861 303 864 307
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1885 303 1888 307
rect 2888 303 2890 307
rect 2894 303 2897 307
rect 2901 303 2904 307
rect 3920 303 3922 307
rect 3926 303 3929 307
rect 3933 303 3936 307
rect 4936 303 4938 307
rect 4942 303 4945 307
rect 4949 303 4952 307
rect 30 271 33 281
rect 86 278 105 281
rect 478 278 497 281
rect 742 278 753 281
rect 838 278 873 281
rect 1102 278 1121 281
rect 14 268 33 271
rect 46 268 70 271
rect 298 268 314 271
rect 458 268 465 271
rect 566 268 569 278
rect 742 277 746 278
rect 770 268 777 271
rect 1094 268 1102 271
rect 1302 271 1305 281
rect 1598 278 1617 281
rect 1806 278 1817 281
rect 1286 268 1305 271
rect 1546 268 1553 271
rect 1746 268 1761 271
rect 1766 268 1774 271
rect 2006 271 2009 281
rect 2150 278 2158 281
rect 2454 278 2465 281
rect 2934 278 2953 281
rect 3490 278 3491 282
rect 3598 278 3609 281
rect 3730 278 3737 281
rect 3158 272 3161 278
rect 3598 277 3602 278
rect 1990 268 2009 271
rect 2962 268 2970 271
rect 3158 268 3162 272
rect 3702 268 3710 271
rect 4030 271 4033 281
rect 4310 278 4321 281
rect 4434 278 4449 281
rect 4854 278 4866 281
rect 5246 278 5265 281
rect 4310 277 4314 278
rect 4630 274 4634 278
rect 4862 277 4866 278
rect 4014 268 4033 271
rect 4101 268 4102 272
rect 4326 268 4345 271
rect 4574 268 4585 271
rect 4702 268 4710 271
rect 4738 268 4745 271
rect 4842 268 4849 271
rect 286 258 302 261
rect 542 258 558 261
rect 758 258 777 261
rect 918 258 926 261
rect 1758 258 1761 268
rect 1830 258 1854 261
rect 2186 258 2193 261
rect 2434 258 2441 261
rect 2870 258 2881 261
rect 3078 258 3097 261
rect 3302 258 3321 261
rect 3626 258 3633 261
rect 3674 258 3689 261
rect 3782 258 3798 261
rect 3846 258 3865 261
rect 3878 258 3886 261
rect 4106 258 4121 261
rect 4310 258 4318 261
rect 4454 258 4473 261
rect 4550 258 4558 261
rect 4794 258 4801 261
rect 4830 258 4849 261
rect 4914 258 4921 261
rect 2650 248 2657 251
rect 2666 248 2670 252
rect 2698 248 2702 252
rect 3094 248 3097 258
rect 3106 248 3110 252
rect 3266 248 3270 252
rect 3318 248 3321 258
rect 3330 248 3334 252
rect 3778 248 3782 252
rect 3862 248 3865 258
rect 4310 257 4314 258
rect 3874 248 3878 252
rect 4170 248 4174 252
rect 1974 242 1978 244
rect 3654 242 3658 244
rect 906 238 909 242
rect 1515 238 1518 242
rect 3930 238 3933 242
rect 269 218 270 222
rect 429 218 430 222
rect 838 218 854 221
rect 3234 218 3235 222
rect 3813 218 3814 222
rect 328 203 330 207
rect 334 203 337 207
rect 341 203 344 207
rect 1352 203 1354 207
rect 1358 203 1361 207
rect 1365 203 1368 207
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2397 203 2400 207
rect 3400 203 3402 207
rect 3406 203 3409 207
rect 3413 203 3416 207
rect 4424 203 4426 207
rect 4430 203 4433 207
rect 4437 203 4440 207
rect 722 188 723 192
rect 1533 188 1534 192
rect 3546 188 3547 192
rect 3570 188 3571 192
rect 3658 188 3659 192
rect 3853 188 3854 192
rect 4958 188 4966 191
rect 5005 188 5006 192
rect 5277 188 5278 192
rect 147 168 150 172
rect 339 168 342 172
rect 3379 168 3382 172
rect 4794 168 4797 172
rect 3670 158 3678 161
rect 4058 158 4065 161
rect 322 148 329 151
rect 1030 148 1038 151
rect 1142 148 1150 151
rect 1654 148 1662 151
rect 1810 148 1817 151
rect 1854 148 1886 151
rect 1910 142 1913 151
rect 2018 148 2025 151
rect 2086 148 2094 151
rect 2174 148 2190 151
rect 2258 148 2265 151
rect 2302 148 2310 151
rect 2366 148 2374 151
rect 2634 148 2641 151
rect 2682 148 2697 151
rect 3050 148 3057 151
rect 3726 148 3734 151
rect 1042 138 1049 141
rect 1666 138 1673 141
rect 2098 138 2105 141
rect 2454 138 2462 141
rect 2718 138 2737 141
rect 2870 138 2889 141
rect 3134 138 3153 141
rect 3446 138 3465 141
rect 3550 141 3553 148
rect 4818 148 4833 151
rect 5110 148 5118 151
rect 3550 138 3561 141
rect 3682 138 3689 141
rect 3874 138 3881 141
rect 3894 138 3913 141
rect 4074 138 4081 141
rect 4490 138 4498 141
rect 4614 138 4633 141
rect 4862 138 4874 141
rect 5062 138 5070 141
rect 366 128 385 131
rect 422 128 441 131
rect 566 128 585 131
rect 1014 131 1018 133
rect 1014 128 1025 131
rect 1198 131 1202 133
rect 1198 128 1209 131
rect 1246 128 1265 131
rect 1486 128 1505 131
rect 1638 131 1642 133
rect 1638 128 1649 131
rect 1990 131 1994 136
rect 1978 128 1994 131
rect 2078 128 2081 138
rect 2230 131 2234 133
rect 2230 128 2241 131
rect 2622 131 2626 133
rect 2326 128 2345 131
rect 2622 128 2633 131
rect 2666 128 2667 132
rect 2718 128 2721 138
rect 2870 128 2873 138
rect 3038 131 3042 133
rect 3038 128 3049 131
rect 3134 128 3137 138
rect 3446 128 3449 138
rect 3502 128 3521 131
rect 3598 128 3617 131
rect 3894 128 3897 138
rect 4190 131 4194 136
rect 4178 128 4194 131
rect 4614 128 4617 138
rect 4726 128 4745 131
rect 366 121 369 128
rect 358 118 369 121
rect 2290 118 2291 122
rect 3714 118 3715 122
rect 848 103 850 107
rect 854 103 857 107
rect 861 103 864 107
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1885 103 1888 107
rect 2888 103 2890 107
rect 2894 103 2897 107
rect 2901 103 2904 107
rect 3920 103 3922 107
rect 3926 103 3929 107
rect 3933 103 3936 107
rect 4936 103 4938 107
rect 4942 103 4945 107
rect 4949 103 4952 107
rect 2358 88 2366 91
rect 190 78 209 81
rect 614 78 625 81
rect 658 78 659 82
rect 850 78 865 81
rect 870 78 889 81
rect 1038 78 1057 81
rect 1158 78 1169 81
rect 1202 78 1203 82
rect 1430 78 1442 81
rect 614 77 618 78
rect 1158 77 1162 78
rect 1438 77 1442 78
rect 110 68 121 71
rect 1526 68 1538 71
rect 1654 71 1657 81
rect 2166 78 2178 81
rect 2174 77 2178 78
rect 2190 74 2194 78
rect 2470 78 2478 81
rect 2514 78 2515 82
rect 2566 78 2585 81
rect 2590 78 2602 81
rect 2470 77 2474 78
rect 2598 77 2602 78
rect 2902 78 2910 81
rect 2614 74 2618 78
rect 1654 68 1673 71
rect 1774 68 1786 71
rect 2262 68 2274 71
rect 2378 68 2386 71
rect 2686 68 2698 71
rect 3238 71 3241 81
rect 3598 78 3617 81
rect 3750 78 3769 81
rect 3902 78 3921 81
rect 3926 78 3942 81
rect 4118 78 4137 81
rect 3222 68 3241 71
rect 3622 68 3634 71
rect 4098 68 4105 71
rect 4398 71 4401 81
rect 4502 78 4514 81
rect 4510 77 4514 78
rect 4526 78 4542 81
rect 4662 78 4674 81
rect 4526 74 4530 78
rect 4670 77 4674 78
rect 5278 72 5282 77
rect 4382 68 4401 71
rect 4638 68 4646 71
rect 118 62 121 68
rect 190 58 193 68
rect 950 58 966 61
rect 1102 58 1110 61
rect 1170 58 1177 61
rect 1362 58 1377 61
rect 2046 58 2062 61
rect 2158 58 2166 61
rect 2482 58 2489 61
rect 2526 58 2542 61
rect 2566 58 2569 68
rect 3234 58 3241 61
rect 3622 62 3625 68
rect 4050 58 4057 61
rect 4310 58 4326 61
rect 4478 58 4497 61
rect 4554 58 4569 61
rect 4638 58 4657 61
rect 4722 58 4729 61
rect 5166 52 5170 54
rect 626 48 633 51
rect 328 3 330 7
rect 334 3 337 7
rect 341 3 344 7
rect 1352 3 1354 7
rect 1358 3 1361 7
rect 1365 3 1368 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2397 3 2400 7
rect 3400 3 3402 7
rect 3406 3 3409 7
rect 3413 3 3416 7
rect 4424 3 4426 7
rect 4430 3 4433 7
rect 4437 3 4440 7
<< m2contact >>
rect 850 5103 854 5107
rect 857 5103 861 5107
rect 1874 5103 1878 5107
rect 1881 5103 1885 5107
rect 2890 5103 2894 5107
rect 2897 5103 2901 5107
rect 3922 5103 3926 5107
rect 3929 5103 3933 5107
rect 4938 5103 4942 5107
rect 4945 5103 4949 5107
rect 518 5088 522 5092
rect 646 5088 650 5092
rect 806 5088 810 5092
rect 950 5088 954 5092
rect 1134 5088 1138 5092
rect 1462 5088 1466 5092
rect 1542 5088 1546 5092
rect 2302 5088 2306 5092
rect 2622 5088 2626 5092
rect 4142 5088 4146 5092
rect 286 5078 290 5082
rect 310 5078 314 5082
rect 326 5078 330 5082
rect 390 5078 394 5082
rect 542 5078 546 5082
rect 630 5078 634 5082
rect 694 5078 698 5082
rect 702 5078 706 5082
rect 814 5078 818 5082
rect 1126 5078 1130 5082
rect 1230 5078 1234 5082
rect 1726 5078 1730 5082
rect 2422 5078 2426 5082
rect 2454 5078 2458 5082
rect 2470 5078 2474 5082
rect 2526 5078 2530 5082
rect 3566 5078 3570 5082
rect 4238 5078 4242 5082
rect 4486 5078 4490 5082
rect 4494 5078 4498 5082
rect 38 5068 42 5072
rect 118 5068 122 5072
rect 150 5068 154 5072
rect 174 5068 178 5072
rect 190 5068 194 5072
rect 326 5068 330 5072
rect 382 5068 386 5072
rect 406 5068 410 5072
rect 446 5068 450 5072
rect 510 5068 514 5072
rect 558 5068 562 5072
rect 622 5068 626 5072
rect 646 5068 650 5072
rect 710 5068 714 5072
rect 726 5068 730 5072
rect 750 5068 754 5072
rect 798 5068 802 5072
rect 838 5068 842 5072
rect 854 5068 858 5072
rect 894 5068 898 5072
rect 910 5068 914 5072
rect 926 5068 930 5072
rect 1054 5068 1058 5072
rect 1182 5068 1186 5072
rect 1230 5068 1234 5072
rect 1246 5068 1250 5072
rect 1278 5068 1282 5072
rect 1342 5068 1346 5072
rect 1534 5068 1538 5072
rect 1582 5068 1586 5072
rect 1670 5068 1674 5072
rect 1742 5068 1746 5072
rect 1822 5068 1826 5072
rect 1934 5068 1938 5072
rect 2126 5068 2130 5072
rect 2222 5068 2226 5072
rect 2318 5068 2322 5072
rect 2414 5068 2418 5072
rect 2438 5068 2442 5072
rect 2486 5068 2490 5072
rect 2502 5068 2506 5072
rect 2542 5068 2546 5072
rect 2638 5068 2642 5072
rect 2750 5068 2754 5072
rect 2766 5068 2770 5072
rect 2790 5068 2794 5072
rect 2894 5068 2898 5072
rect 3038 5068 3042 5072
rect 3054 5068 3058 5072
rect 3070 5068 3074 5072
rect 3110 5068 3114 5072
rect 3150 5068 3154 5072
rect 3190 5068 3194 5072
rect 3206 5068 3210 5072
rect 3446 5068 3450 5072
rect 3918 5068 3922 5072
rect 3966 5068 3970 5072
rect 4038 5068 4042 5072
rect 4070 5068 4074 5072
rect 4222 5068 4226 5072
rect 4406 5068 4410 5072
rect 4590 5068 4594 5072
rect 4686 5068 4690 5072
rect 4782 5068 4786 5072
rect 4862 5068 4866 5072
rect 4982 5068 4986 5072
rect 5014 5068 5018 5072
rect 5022 5068 5026 5072
rect 5054 5068 5058 5072
rect 5222 5068 5226 5072
rect 5230 5068 5234 5072
rect 46 5058 50 5062
rect 142 5058 146 5062
rect 174 5058 178 5062
rect 206 5059 210 5063
rect 350 5058 354 5062
rect 374 5058 378 5062
rect 438 5058 442 5062
rect 462 5058 466 5062
rect 494 5058 498 5062
rect 502 5058 506 5062
rect 534 5058 538 5062
rect 566 5058 570 5062
rect 590 5058 594 5062
rect 654 5058 658 5062
rect 726 5058 730 5062
rect 750 5058 754 5062
rect 782 5058 786 5062
rect 878 5058 882 5062
rect 1038 5059 1042 5063
rect 1070 5058 1074 5062
rect 1118 5058 1122 5062
rect 1190 5058 1194 5062
rect 1254 5058 1258 5062
rect 1278 5058 1282 5062
rect 1374 5059 1378 5063
rect 1406 5058 1410 5062
rect 1470 5058 1474 5062
rect 1558 5058 1562 5062
rect 1566 5058 1570 5062
rect 1806 5058 1810 5062
rect 1846 5058 1850 5062
rect 1966 5058 1970 5062
rect 1982 5058 1986 5062
rect 2054 5058 2058 5062
rect 2086 5059 2090 5063
rect 2150 5058 2154 5062
rect 2246 5058 2250 5062
rect 2342 5058 2346 5062
rect 2446 5058 2450 5062
rect 2478 5058 2482 5062
rect 2510 5058 2514 5062
rect 2558 5059 2562 5063
rect 2662 5058 2666 5062
rect 2742 5058 2746 5062
rect 2774 5058 2778 5062
rect 2814 5058 2818 5062
rect 2918 5058 2922 5062
rect 2942 5058 2946 5062
rect 2950 5058 2954 5062
rect 3022 5059 3026 5063
rect 3062 5058 3066 5062
rect 3142 5058 3146 5062
rect 3158 5058 3162 5062
rect 3166 5058 3170 5062
rect 3174 5058 3178 5062
rect 3198 5058 3202 5062
rect 3262 5058 3266 5062
rect 3342 5058 3346 5062
rect 3366 5058 3370 5062
rect 3470 5058 3474 5062
rect 3494 5058 3498 5062
rect 3534 5058 3538 5062
rect 3550 5058 3554 5062
rect 3558 5058 3562 5062
rect 3582 5058 3586 5062
rect 3630 5058 3634 5062
rect 3654 5058 3658 5062
rect 3702 5058 3706 5062
rect 3710 5058 3714 5062
rect 3726 5058 3730 5062
rect 3734 5058 3738 5062
rect 3766 5059 3770 5063
rect 3798 5058 3802 5062
rect 3838 5058 3842 5062
rect 3942 5058 3946 5062
rect 4078 5058 4082 5062
rect 4206 5059 4210 5063
rect 4286 5058 4290 5062
rect 4310 5058 4314 5062
rect 4398 5058 4402 5062
rect 4574 5059 4578 5063
rect 4670 5059 4674 5063
rect 4766 5059 4770 5063
rect 4902 5058 4906 5062
rect 4926 5058 4930 5062
rect 4990 5058 4994 5062
rect 5046 5058 5050 5062
rect 5094 5058 5098 5062
rect 5110 5058 5114 5062
rect 5238 5058 5242 5062
rect 118 5048 122 5052
rect 158 5048 162 5052
rect 294 5048 298 5052
rect 454 5048 458 5052
rect 486 5048 490 5052
rect 598 5048 602 5052
rect 606 5048 610 5052
rect 742 5048 746 5052
rect 758 5048 762 5052
rect 782 5048 786 5052
rect 822 5048 826 5052
rect 830 5048 834 5052
rect 838 5048 842 5052
rect 862 5048 866 5052
rect 918 5048 922 5052
rect 942 5048 946 5052
rect 1078 5048 1082 5052
rect 1094 5048 1098 5052
rect 1270 5048 1274 5052
rect 3086 5048 3090 5052
rect 3126 5048 3130 5052
rect 3182 5048 3186 5052
rect 102 5038 106 5042
rect 470 5038 474 5042
rect 582 5038 586 5042
rect 590 5038 594 5042
rect 734 5038 738 5042
rect 2190 5038 2194 5042
rect 3214 5038 3218 5042
rect 3422 5038 3426 5042
rect 5006 5038 5010 5042
rect 5030 5038 5034 5042
rect 5254 5038 5258 5042
rect 5302 5038 5306 5042
rect 462 5028 466 5032
rect 2958 5028 2962 5032
rect 4470 5028 4474 5032
rect 390 5018 394 5022
rect 542 5018 546 5022
rect 574 5018 578 5022
rect 614 5018 618 5022
rect 934 5018 938 5022
rect 1262 5018 1266 5022
rect 1654 5018 1658 5022
rect 1902 5018 1906 5022
rect 2014 5018 2018 5022
rect 2022 5018 2026 5022
rect 2206 5018 2210 5022
rect 2398 5018 2402 5022
rect 2718 5018 2722 5022
rect 3686 5018 3690 5022
rect 3862 5018 3866 5022
rect 3982 5018 3986 5022
rect 4134 5018 4138 5022
rect 4246 5018 4250 5022
rect 4358 5018 4362 5022
rect 4470 5018 4474 5022
rect 4502 5018 4506 5022
rect 4510 5018 4514 5022
rect 4606 5018 4610 5022
rect 4702 5018 4706 5022
rect 4806 5018 4810 5022
rect 4958 5018 4962 5022
rect 4990 5018 4994 5022
rect 5046 5018 5050 5022
rect 5150 5018 5154 5022
rect 5166 5018 5170 5022
rect 5238 5018 5242 5022
rect 330 5003 334 5007
rect 337 5003 341 5007
rect 1354 5003 1358 5007
rect 1361 5003 1365 5007
rect 2386 5003 2390 5007
rect 2393 5003 2397 5007
rect 3402 5003 3406 5007
rect 3409 5003 3413 5007
rect 4426 5003 4430 5007
rect 4433 5003 4437 5007
rect 6 4988 10 4992
rect 158 4988 162 4992
rect 222 4988 226 4992
rect 502 4988 506 4992
rect 662 4988 666 4992
rect 734 4988 738 4992
rect 1342 4988 1346 4992
rect 1438 4988 1442 4992
rect 1558 4988 1562 4992
rect 1654 4988 1658 4992
rect 1942 4988 1946 4992
rect 2134 4988 2138 4992
rect 2350 4988 2354 4992
rect 2454 4988 2458 4992
rect 2518 4988 2522 4992
rect 3630 4988 3634 4992
rect 3702 4988 3706 4992
rect 4342 4988 4346 4992
rect 4566 4988 4570 4992
rect 4782 4988 4786 4992
rect 278 4978 282 4982
rect 958 4978 962 4982
rect 166 4968 170 4972
rect 286 4968 290 4972
rect 478 4968 482 4972
rect 534 4968 538 4972
rect 742 4968 746 4972
rect 830 4968 834 4972
rect 878 4968 882 4972
rect 1222 4968 1226 4972
rect 1350 4968 1354 4972
rect 1550 4968 1554 4972
rect 2046 4968 2050 4972
rect 2318 4968 2322 4972
rect 2854 4968 2858 4972
rect 3230 4968 3234 4972
rect 3246 4968 3250 4972
rect 3286 4968 3290 4972
rect 3430 4968 3434 4972
rect 3446 4968 3450 4972
rect 3526 4968 3530 4972
rect 3542 4968 3546 4972
rect 3822 4968 3826 4972
rect 3846 4968 3850 4972
rect 102 4958 106 4962
rect 150 4958 154 4962
rect 254 4958 258 4962
rect 270 4958 274 4962
rect 326 4958 330 4962
rect 430 4958 434 4962
rect 462 4958 466 4962
rect 518 4958 522 4962
rect 622 4958 626 4962
rect 638 4958 642 4962
rect 702 4958 706 4962
rect 726 4958 730 4962
rect 790 4958 794 4962
rect 846 4958 850 4962
rect 894 4958 898 4962
rect 902 4958 906 4962
rect 950 4958 954 4962
rect 982 4958 986 4962
rect 1014 4958 1018 4962
rect 1046 4958 1050 4962
rect 1062 4958 1066 4962
rect 1294 4958 1298 4962
rect 1918 4958 1922 4962
rect 38 4948 42 4952
rect 70 4947 74 4951
rect 110 4948 114 4952
rect 118 4948 122 4952
rect 134 4948 138 4952
rect 158 4948 162 4952
rect 182 4948 186 4952
rect 214 4948 218 4952
rect 246 4948 250 4952
rect 278 4948 282 4952
rect 310 4948 314 4952
rect 374 4948 378 4952
rect 422 4948 426 4952
rect 446 4948 450 4952
rect 470 4948 474 4952
rect 494 4948 498 4952
rect 534 4948 538 4952
rect 574 4948 578 4952
rect 598 4948 602 4952
rect 622 4948 626 4952
rect 694 4948 698 4952
rect 734 4948 738 4952
rect 790 4948 794 4952
rect 830 4948 834 4952
rect 846 4948 850 4952
rect 974 4948 978 4952
rect 1046 4948 1050 4952
rect 1134 4947 1138 4951
rect 1174 4948 1178 4952
rect 1198 4948 1202 4952
rect 1230 4948 1234 4952
rect 1278 4948 1282 4952
rect 1310 4948 1314 4952
rect 1334 4948 1338 4952
rect 1342 4948 1346 4952
rect 1414 4948 1418 4952
rect 1430 4948 1434 4952
rect 1454 4948 1458 4952
rect 1494 4948 1498 4952
rect 1510 4948 1514 4952
rect 1590 4948 1594 4952
rect 1614 4948 1618 4952
rect 1710 4948 1714 4952
rect 1734 4948 1738 4952
rect 1806 4948 1810 4952
rect 2070 4958 2074 4962
rect 2222 4958 2226 4962
rect 2422 4958 2426 4962
rect 2574 4958 2578 4962
rect 2630 4958 2634 4962
rect 2662 4958 2666 4962
rect 2934 4958 2938 4962
rect 3006 4958 3010 4962
rect 1942 4948 1946 4952
rect 1998 4947 2002 4951
rect 2086 4948 2090 4952
rect 2126 4948 2130 4952
rect 2150 4948 2154 4952
rect 2158 4948 2162 4952
rect 2174 4948 2178 4952
rect 2198 4948 2202 4952
rect 2206 4948 2210 4952
rect 2254 4947 2258 4951
rect 2326 4948 2330 4952
rect 2358 4948 2362 4952
rect 2390 4948 2394 4952
rect 2446 4948 2450 4952
rect 2478 4948 2482 4952
rect 2486 4948 2490 4952
rect 2510 4948 2514 4952
rect 2534 4948 2538 4952
rect 2542 4948 2546 4952
rect 2558 4948 2562 4952
rect 2582 4948 2586 4952
rect 2614 4948 2618 4952
rect 2638 4948 2642 4952
rect 2694 4947 2698 4951
rect 2798 4948 2802 4952
rect 2862 4948 2866 4952
rect 2926 4948 2930 4952
rect 2958 4948 2962 4952
rect 2990 4948 2994 4952
rect 3046 4948 3050 4952
rect 3078 4947 3082 4951
rect 3110 4948 3114 4952
rect 3118 4948 3122 4952
rect 3150 4948 3154 4952
rect 3190 4948 3194 4952
rect 3262 4948 3266 4952
rect 3270 4948 3274 4952
rect 3558 4958 3562 4962
rect 3646 4958 3650 4962
rect 3662 4958 3666 4962
rect 3678 4958 3682 4962
rect 4158 4958 4162 4962
rect 3302 4948 3306 4952
rect 3350 4948 3354 4952
rect 3374 4948 3378 4952
rect 3462 4948 3466 4952
rect 3494 4947 3498 4951
rect 3542 4948 3546 4952
rect 3558 4948 3562 4952
rect 3574 4948 3578 4952
rect 3590 4948 3594 4952
rect 3630 4948 3634 4952
rect 3662 4948 3666 4952
rect 3694 4948 3698 4952
rect 3718 4948 3722 4952
rect 3726 4948 3730 4952
rect 3758 4947 3762 4951
rect 3790 4948 3794 4952
rect 3886 4948 3890 4952
rect 3974 4948 3978 4952
rect 4070 4948 4074 4952
rect 4094 4948 4098 4952
rect 4142 4948 4146 4952
rect 4494 4958 4498 4962
rect 4510 4958 4514 4962
rect 4174 4948 4178 4952
rect 4182 4948 4186 4952
rect 4230 4948 4234 4952
rect 4254 4948 4258 4952
rect 4294 4948 4298 4952
rect 4334 4948 4338 4952
rect 4358 4948 4362 4952
rect 4366 4948 4370 4952
rect 4430 4948 4434 4952
rect 4478 4948 4482 4952
rect 4518 4948 4522 4952
rect 4558 4948 4562 4952
rect 4582 4948 4586 4952
rect 4590 4948 4594 4952
rect 4606 4948 4610 4952
rect 4718 4948 4722 4952
rect 4774 4948 4778 4952
rect 4806 4948 4810 4952
rect 4838 4947 4842 4951
rect 4870 4948 4874 4952
rect 4910 4948 4914 4952
rect 5022 4948 5026 4952
rect 5038 4948 5042 4952
rect 5078 4948 5082 4952
rect 5102 4948 5106 4952
rect 5174 4948 5178 4952
rect 126 4938 130 4942
rect 190 4938 194 4942
rect 222 4938 226 4942
rect 238 4938 242 4942
rect 302 4938 306 4942
rect 350 4938 354 4942
rect 366 4938 370 4942
rect 398 4938 402 4942
rect 414 4938 418 4942
rect 454 4938 458 4942
rect 542 4938 546 4942
rect 550 4938 554 4942
rect 566 4938 570 4942
rect 606 4938 610 4942
rect 614 4938 618 4942
rect 646 4938 650 4942
rect 694 4938 698 4942
rect 718 4938 722 4942
rect 758 4938 762 4942
rect 774 4938 778 4942
rect 782 4938 786 4942
rect 814 4938 818 4942
rect 822 4938 826 4942
rect 870 4938 874 4942
rect 918 4938 922 4942
rect 934 4938 938 4942
rect 982 4938 986 4942
rect 990 4938 994 4942
rect 1006 4938 1010 4942
rect 1038 4938 1042 4942
rect 1150 4938 1154 4942
rect 1166 4938 1170 4942
rect 1222 4938 1226 4942
rect 1270 4938 1274 4942
rect 1406 4938 1410 4942
rect 1486 4938 1490 4942
rect 1902 4938 1906 4942
rect 1950 4938 1954 4942
rect 1982 4938 1986 4942
rect 2094 4938 2098 4942
rect 2238 4938 2242 4942
rect 2334 4938 2338 4942
rect 2406 4938 2410 4942
rect 2470 4938 2474 4942
rect 2486 4938 2490 4942
rect 2550 4938 2554 4942
rect 2646 4938 2650 4942
rect 2702 4938 2706 4942
rect 2774 4938 2778 4942
rect 2790 4938 2794 4942
rect 2870 4938 2874 4942
rect 2942 4938 2946 4942
rect 2958 4938 2962 4942
rect 3166 4938 3170 4942
rect 3254 4938 3258 4942
rect 3310 4938 3314 4942
rect 3550 4938 3554 4942
rect 3582 4938 3586 4942
rect 3614 4938 3618 4942
rect 3622 4938 3626 4942
rect 3654 4938 3658 4942
rect 3766 4938 3770 4942
rect 3870 4938 3874 4942
rect 3982 4938 3986 4942
rect 4134 4938 4138 4942
rect 4190 4938 4194 4942
rect 4302 4938 4306 4942
rect 4406 4938 4410 4942
rect 4454 4938 4458 4942
rect 4478 4938 4482 4942
rect 4526 4938 4530 4942
rect 4638 4938 4642 4942
rect 4654 4938 4658 4942
rect 4694 4938 4698 4942
rect 4742 4938 4746 4942
rect 4798 4938 4802 4942
rect 4822 4938 4826 4942
rect 4974 4938 4978 4942
rect 5014 4938 5018 4942
rect 5110 4938 5114 4942
rect 5150 4938 5154 4942
rect 5302 4938 5306 4942
rect 134 4928 138 4932
rect 206 4928 210 4932
rect 254 4928 258 4932
rect 342 4928 346 4932
rect 382 4928 386 4932
rect 470 4928 474 4932
rect 510 4928 514 4932
rect 550 4928 554 4932
rect 758 4928 762 4932
rect 926 4928 930 4932
rect 1246 4928 1250 4932
rect 1382 4928 1386 4932
rect 1398 4928 1402 4932
rect 1894 4928 1898 4932
rect 1958 4928 1962 4932
rect 2070 4928 2074 4932
rect 2110 4928 2114 4932
rect 2190 4928 2194 4932
rect 2222 4928 2226 4932
rect 2390 4928 2394 4932
rect 2422 4928 2426 4932
rect 2430 4928 2434 4932
rect 2598 4928 2602 4932
rect 2662 4928 2666 4932
rect 2878 4928 2882 4932
rect 2894 4928 2898 4932
rect 2910 4928 2914 4932
rect 2966 4928 2970 4932
rect 3126 4928 3130 4932
rect 3230 4928 3234 4932
rect 4318 4928 4322 4932
rect 4542 4928 4546 4932
rect 4758 4928 4762 4932
rect 5006 4928 5010 4932
rect 5078 4928 5082 4932
rect 198 4918 202 4922
rect 358 4918 362 4922
rect 406 4918 410 4922
rect 430 4918 434 4922
rect 582 4918 586 4922
rect 950 4918 954 4922
rect 1070 4918 1074 4922
rect 1326 4918 1330 4922
rect 1862 4918 1866 4922
rect 1878 4918 1882 4922
rect 2062 4918 2066 4922
rect 2102 4918 2106 4922
rect 2574 4918 2578 4922
rect 2590 4918 2594 4922
rect 2630 4918 2634 4922
rect 2758 4918 2762 4922
rect 2974 4918 2978 4922
rect 3318 4918 3322 4922
rect 3414 4918 3418 4922
rect 3830 4918 3834 4922
rect 4030 4918 4034 4922
rect 4038 4918 4042 4922
rect 4198 4918 4202 4922
rect 4310 4918 4314 4922
rect 4374 4918 4378 4922
rect 4534 4918 4538 4922
rect 4902 4918 4906 4922
rect 4998 4918 5002 4922
rect 5038 4918 5042 4922
rect 5230 4918 5234 4922
rect 5246 4918 5250 4922
rect 850 4903 854 4907
rect 857 4903 861 4907
rect 1874 4903 1878 4907
rect 1881 4903 1885 4907
rect 2890 4903 2894 4907
rect 2897 4903 2901 4907
rect 3922 4903 3926 4907
rect 3929 4903 3933 4907
rect 4938 4903 4942 4907
rect 4945 4903 4949 4907
rect 190 4888 194 4892
rect 502 4888 506 4892
rect 534 4888 538 4892
rect 566 4888 570 4892
rect 630 4888 634 4892
rect 694 4888 698 4892
rect 758 4888 762 4892
rect 782 4888 786 4892
rect 870 4888 874 4892
rect 942 4888 946 4892
rect 998 4888 1002 4892
rect 1014 4888 1018 4892
rect 1054 4888 1058 4892
rect 1270 4888 1274 4892
rect 1422 4888 1426 4892
rect 1430 4888 1434 4892
rect 1470 4888 1474 4892
rect 1862 4888 1866 4892
rect 1998 4888 2002 4892
rect 2558 4888 2562 4892
rect 2662 4888 2666 4892
rect 2854 4888 2858 4892
rect 3014 4888 3018 4892
rect 3230 4888 3234 4892
rect 3286 4888 3290 4892
rect 3590 4888 3594 4892
rect 3654 4888 3658 4892
rect 3782 4888 3786 4892
rect 4006 4888 4010 4892
rect 4094 4888 4098 4892
rect 4206 4888 4210 4892
rect 4278 4888 4282 4892
rect 4326 4888 4330 4892
rect 4646 4888 4650 4892
rect 4966 4888 4970 4892
rect 5086 4888 5090 4892
rect 102 4878 106 4882
rect 118 4878 122 4882
rect 166 4878 170 4882
rect 574 4878 578 4882
rect 638 4878 642 4882
rect 678 4878 682 4882
rect 766 4878 770 4882
rect 814 4878 818 4882
rect 862 4878 866 4882
rect 918 4878 922 4882
rect 126 4868 130 4872
rect 182 4868 186 4872
rect 246 4868 250 4872
rect 390 4868 394 4872
rect 454 4868 458 4872
rect 494 4868 498 4872
rect 510 4868 514 4872
rect 542 4868 546 4872
rect 558 4868 562 4872
rect 574 4868 578 4872
rect 622 4868 626 4872
rect 638 4868 642 4872
rect 694 4868 698 4872
rect 734 4868 738 4872
rect 774 4868 778 4872
rect 806 4868 810 4872
rect 854 4868 858 4872
rect 950 4868 954 4872
rect 1006 4878 1010 4882
rect 1046 4878 1050 4882
rect 1238 4878 1242 4882
rect 1350 4878 1354 4882
rect 1478 4878 1482 4882
rect 1590 4878 1594 4882
rect 2030 4878 2034 4882
rect 2166 4878 2170 4882
rect 2414 4878 2418 4882
rect 2494 4878 2498 4882
rect 2566 4878 2570 4882
rect 2654 4878 2658 4882
rect 2670 4878 2674 4882
rect 2774 4878 2778 4882
rect 2982 4878 2986 4882
rect 3134 4878 3138 4882
rect 3166 4878 3170 4882
rect 3318 4878 3322 4882
rect 4038 4878 4042 4882
rect 4102 4878 4106 4882
rect 4110 4878 4114 4882
rect 4126 4878 4130 4882
rect 4142 4878 4146 4882
rect 4246 4878 4250 4882
rect 4262 4878 4266 4882
rect 974 4868 978 4872
rect 1078 4868 1082 4872
rect 1166 4868 1170 4872
rect 1174 4868 1178 4872
rect 1214 4868 1218 4872
rect 1230 4868 1234 4872
rect 1254 4868 1258 4872
rect 1390 4868 1394 4872
rect 38 4858 42 4862
rect 70 4859 74 4863
rect 102 4858 106 4862
rect 134 4858 138 4862
rect 174 4858 178 4862
rect 206 4858 210 4862
rect 230 4858 234 4862
rect 294 4858 298 4862
rect 318 4858 322 4862
rect 342 4858 346 4862
rect 374 4858 378 4862
rect 430 4858 434 4862
rect 462 4858 466 4862
rect 486 4858 490 4862
rect 518 4858 522 4862
rect 550 4858 554 4862
rect 582 4858 586 4862
rect 662 4858 666 4862
rect 678 4858 682 4862
rect 702 4858 706 4862
rect 742 4858 746 4862
rect 782 4858 786 4862
rect 798 4858 802 4862
rect 862 4858 866 4862
rect 878 4858 882 4862
rect 886 4858 890 4862
rect 926 4858 930 4862
rect 1446 4866 1450 4870
rect 1454 4868 1458 4872
rect 4294 4878 4298 4882
rect 4446 4878 4450 4882
rect 4486 4878 4490 4882
rect 4678 4878 4682 4882
rect 4870 4878 4874 4882
rect 5046 4878 5050 4882
rect 5054 4878 5058 4882
rect 1502 4868 1506 4872
rect 1654 4868 1658 4872
rect 1726 4868 1730 4872
rect 1742 4868 1746 4872
rect 1910 4868 1914 4872
rect 1990 4868 1994 4872
rect 2046 4868 2050 4872
rect 2238 4868 2242 4872
rect 2302 4868 2306 4872
rect 2582 4868 2586 4872
rect 2678 4868 2682 4872
rect 2862 4868 2866 4872
rect 2958 4868 2962 4872
rect 2966 4868 2970 4872
rect 2990 4868 2994 4872
rect 3022 4868 3026 4872
rect 3070 4868 3074 4872
rect 3118 4868 3122 4872
rect 3246 4868 3250 4872
rect 3278 4868 3282 4872
rect 3326 4868 3330 4872
rect 3398 4868 3402 4872
rect 3502 4868 3506 4872
rect 3566 4868 3570 4872
rect 3622 4868 3626 4872
rect 3630 4868 3634 4872
rect 3662 4868 3666 4872
rect 3694 4868 3698 4872
rect 3742 4868 3746 4872
rect 3750 4868 3754 4872
rect 3806 4868 3810 4872
rect 3926 4868 3930 4872
rect 3958 4868 3962 4872
rect 3982 4868 3986 4872
rect 3998 4868 4002 4872
rect 4046 4868 4050 4872
rect 4086 4868 4090 4872
rect 4286 4868 4290 4872
rect 4310 4868 4314 4872
rect 4406 4868 4410 4872
rect 4574 4868 4578 4872
rect 4718 4868 4722 4872
rect 4974 4868 4978 4872
rect 5030 4868 5034 4872
rect 5070 4868 5074 4872
rect 5166 4868 5170 4872
rect 5182 4868 5186 4872
rect 5254 4868 5258 4872
rect 982 4858 986 4862
rect 1022 4858 1026 4862
rect 1030 4858 1034 4862
rect 1078 4858 1082 4862
rect 1094 4858 1098 4862
rect 1126 4858 1130 4862
rect 1182 4858 1186 4862
rect 1222 4858 1226 4862
rect 1326 4858 1330 4862
rect 1406 4858 1410 4862
rect 1462 4858 1466 4862
rect 1582 4858 1586 4862
rect 1662 4858 1666 4862
rect 1766 4858 1770 4862
rect 1846 4858 1850 4862
rect 1854 4858 1858 4862
rect 1878 4858 1882 4862
rect 1982 4858 1986 4862
rect 2014 4858 2018 4862
rect 2070 4858 2074 4862
rect 2150 4858 2154 4862
rect 2158 4858 2162 4862
rect 2182 4858 2186 4862
rect 2222 4859 2226 4863
rect 2326 4858 2330 4862
rect 2350 4858 2354 4862
rect 2430 4858 2434 4862
rect 2454 4858 2458 4862
rect 2462 4858 2466 4862
rect 2502 4858 2506 4862
rect 2614 4858 2618 4862
rect 2622 4858 2626 4862
rect 2630 4858 2634 4862
rect 2646 4858 2650 4862
rect 2742 4858 2746 4862
rect 2782 4858 2786 4862
rect 2894 4858 2898 4862
rect 2902 4858 2906 4862
rect 2926 4858 2930 4862
rect 2998 4858 3002 4862
rect 3030 4858 3034 4862
rect 3078 4858 3082 4862
rect 3086 4858 3090 4862
rect 3166 4859 3170 4863
rect 3198 4858 3202 4862
rect 3262 4858 3266 4862
rect 3270 4858 3274 4862
rect 3302 4858 3306 4862
rect 3334 4858 3338 4862
rect 3382 4858 3386 4862
rect 3438 4858 3442 4862
rect 3462 4858 3466 4862
rect 3510 4858 3514 4862
rect 3542 4858 3546 4862
rect 3550 4858 3554 4862
rect 3574 4858 3578 4862
rect 3614 4858 3618 4862
rect 3630 4858 3634 4862
rect 3670 4858 3674 4862
rect 3734 4858 3738 4862
rect 3758 4858 3762 4862
rect 3798 4858 3802 4862
rect 3846 4858 3850 4862
rect 3870 4858 3874 4862
rect 3934 4858 3938 4862
rect 3974 4858 3978 4862
rect 3990 4858 3994 4862
rect 4022 4858 4026 4862
rect 4054 4858 4058 4862
rect 4078 4858 4082 4862
rect 4126 4858 4130 4862
rect 4150 4858 4154 4862
rect 4190 4858 4194 4862
rect 4214 4858 4218 4862
rect 4222 4858 4226 4862
rect 4230 4858 4234 4862
rect 4238 4858 4242 4862
rect 4270 4858 4274 4862
rect 4302 4858 4306 4862
rect 4318 4858 4322 4862
rect 4382 4858 4386 4862
rect 4422 4858 4426 4862
rect 4494 4858 4498 4862
rect 4606 4858 4610 4862
rect 4614 4858 4618 4862
rect 4630 4858 4634 4862
rect 4686 4858 4690 4862
rect 4694 4858 4698 4862
rect 4790 4858 4794 4862
rect 4878 4858 4882 4862
rect 5006 4858 5010 4862
rect 5014 4858 5018 4862
rect 5022 4858 5026 4862
rect 5078 4858 5082 4862
rect 5142 4858 5146 4862
rect 5262 4858 5266 4862
rect 5286 4858 5290 4862
rect 150 4848 154 4852
rect 166 4848 170 4852
rect 214 4848 218 4852
rect 270 4848 274 4852
rect 310 4848 314 4852
rect 358 4848 362 4852
rect 414 4848 418 4852
rect 422 4848 426 4852
rect 478 4848 482 4852
rect 526 4848 530 4852
rect 606 4848 610 4852
rect 646 4848 650 4852
rect 814 4848 818 4852
rect 998 4848 1002 4852
rect 1086 4848 1090 4852
rect 1118 4848 1122 4852
rect 1150 4848 1154 4852
rect 1182 4848 1186 4852
rect 1198 4848 1202 4852
rect 1206 4848 1210 4852
rect 2438 4848 2442 4852
rect 3014 4848 3018 4852
rect 3054 4848 3058 4852
rect 3590 4848 3594 4852
rect 3614 4848 3618 4852
rect 3654 4848 3658 4852
rect 3670 4848 3674 4852
rect 3694 4848 3698 4852
rect 3710 4848 3714 4852
rect 3774 4848 3778 4852
rect 3950 4848 3954 4852
rect 4070 4848 4074 4852
rect 5278 4848 5282 4852
rect 254 4838 258 4842
rect 286 4838 290 4842
rect 326 4838 330 4842
rect 398 4838 402 4842
rect 438 4838 442 4842
rect 1102 4838 1106 4842
rect 1134 4838 1138 4842
rect 3350 4838 3354 4842
rect 3494 4838 3498 4842
rect 3526 4838 3530 4842
rect 3598 4838 3602 4842
rect 3902 4838 3906 4842
rect 5302 4838 5306 4842
rect 1030 4828 1034 4832
rect 6 4818 10 4822
rect 102 4818 106 4822
rect 134 4818 138 4822
rect 278 4818 282 4822
rect 318 4818 322 4822
rect 430 4818 434 4822
rect 462 4818 466 4822
rect 870 4818 874 4822
rect 1094 4818 1098 4822
rect 1126 4818 1130 4822
rect 1158 4818 1162 4822
rect 1238 4818 1242 4822
rect 1510 4818 1514 4822
rect 1630 4818 1634 4822
rect 1838 4818 1842 4822
rect 1966 4818 1970 4822
rect 2142 4818 2146 4822
rect 2286 4818 2290 4822
rect 2638 4818 2642 4822
rect 2982 4818 2986 4822
rect 3030 4818 3034 4822
rect 3374 4818 3378 4822
rect 3734 4818 3738 4822
rect 4054 4818 4058 4822
rect 4134 4818 4138 4822
rect 4166 4818 4170 4822
rect 4254 4818 4258 4822
rect 4430 4818 4434 4822
rect 4550 4818 4554 4822
rect 4734 4818 4738 4822
rect 5046 4818 5050 4822
rect 5054 4818 5058 4822
rect 5086 4818 5090 4822
rect 5238 4818 5242 4822
rect 5262 4818 5266 4822
rect 330 4803 334 4807
rect 337 4803 341 4807
rect 1354 4803 1358 4807
rect 1361 4803 1365 4807
rect 2386 4803 2390 4807
rect 2393 4803 2397 4807
rect 3402 4803 3406 4807
rect 3409 4803 3413 4807
rect 4426 4803 4430 4807
rect 4433 4803 4437 4807
rect 110 4788 114 4792
rect 150 4788 154 4792
rect 326 4788 330 4792
rect 374 4788 378 4792
rect 422 4788 426 4792
rect 502 4788 506 4792
rect 518 4788 522 4792
rect 646 4788 650 4792
rect 654 4788 658 4792
rect 774 4788 778 4792
rect 974 4788 978 4792
rect 1502 4788 1506 4792
rect 1862 4788 1866 4792
rect 2190 4788 2194 4792
rect 3478 4788 3482 4792
rect 3582 4788 3586 4792
rect 4022 4788 4026 4792
rect 4118 4788 4122 4792
rect 622 4778 626 4782
rect 798 4778 802 4782
rect 142 4768 146 4772
rect 382 4768 386 4772
rect 414 4768 418 4772
rect 662 4768 666 4772
rect 814 4768 818 4772
rect 910 4768 914 4772
rect 1022 4768 1026 4772
rect 1382 4768 1386 4772
rect 2102 4768 2106 4772
rect 2830 4768 2834 4772
rect 4582 4768 4586 4772
rect 78 4758 82 4762
rect 126 4758 130 4762
rect 190 4758 194 4762
rect 206 4758 210 4762
rect 230 4758 234 4762
rect 366 4758 370 4762
rect 398 4758 402 4762
rect 430 4758 434 4762
rect 534 4758 538 4762
rect 614 4758 618 4762
rect 734 4758 738 4762
rect 758 4758 762 4762
rect 846 4758 850 4762
rect 982 4758 986 4762
rect 1038 4758 1042 4762
rect 1046 4758 1050 4762
rect 1158 4758 1162 4762
rect 1166 4758 1170 4762
rect 1246 4758 1250 4762
rect 1318 4758 1322 4762
rect 1334 4758 1338 4762
rect 2158 4758 2162 4762
rect 2254 4758 2258 4762
rect 3046 4758 3050 4762
rect 3702 4758 3706 4762
rect 118 4748 122 4752
rect 142 4748 146 4752
rect 166 4748 170 4752
rect 190 4748 194 4752
rect 230 4748 234 4752
rect 6 4738 10 4742
rect 54 4738 58 4742
rect 62 4738 66 4742
rect 78 4738 82 4742
rect 158 4738 162 4742
rect 190 4738 194 4742
rect 214 4738 218 4742
rect 262 4747 266 4751
rect 390 4748 394 4752
rect 422 4748 426 4752
rect 462 4748 466 4752
rect 486 4748 490 4752
rect 518 4748 522 4752
rect 542 4748 546 4752
rect 590 4748 594 4752
rect 598 4748 602 4752
rect 606 4748 610 4752
rect 670 4748 674 4752
rect 678 4748 682 4752
rect 734 4748 738 4752
rect 798 4748 802 4752
rect 814 4748 818 4752
rect 830 4748 834 4752
rect 854 4748 858 4752
rect 918 4748 922 4752
rect 950 4748 954 4752
rect 974 4748 978 4752
rect 982 4748 986 4752
rect 998 4748 1002 4752
rect 1030 4748 1034 4752
rect 1078 4748 1082 4752
rect 1102 4748 1106 4752
rect 1142 4748 1146 4752
rect 1174 4748 1178 4752
rect 1182 4748 1186 4752
rect 1198 4748 1202 4752
rect 1206 4748 1210 4752
rect 1238 4748 1242 4752
rect 1262 4748 1266 4752
rect 1278 4748 1282 4752
rect 1294 4748 1298 4752
rect 246 4738 250 4742
rect 342 4738 346 4742
rect 438 4738 442 4742
rect 470 4738 474 4742
rect 494 4738 498 4742
rect 510 4738 514 4742
rect 550 4738 554 4742
rect 558 4738 562 4742
rect 566 4738 570 4742
rect 1446 4747 1450 4751
rect 1486 4748 1490 4752
rect 1510 4748 1514 4752
rect 1518 4748 1522 4752
rect 1534 4748 1538 4752
rect 1558 4748 1562 4752
rect 1566 4748 1570 4752
rect 1574 4748 1578 4752
rect 1622 4748 1626 4752
rect 1654 4748 1658 4752
rect 590 4738 594 4742
rect 638 4738 642 4742
rect 702 4738 706 4742
rect 750 4738 754 4742
rect 790 4738 794 4742
rect 822 4738 826 4742
rect 886 4740 890 4744
rect 894 4738 898 4742
rect 942 4738 946 4742
rect 1006 4738 1010 4742
rect 1054 4738 1058 4742
rect 1070 4738 1074 4742
rect 1110 4738 1114 4742
rect 1134 4738 1138 4742
rect 1190 4738 1194 4742
rect 1270 4738 1274 4742
rect 1286 4738 1290 4742
rect 1302 4738 1306 4742
rect 1334 4738 1338 4742
rect 1342 4738 1346 4742
rect 1366 4738 1370 4742
rect 1462 4738 1466 4742
rect 1582 4738 1586 4742
rect 1646 4738 1650 4742
rect 1686 4748 1690 4752
rect 1694 4748 1698 4752
rect 1806 4748 1810 4752
rect 1854 4748 1858 4752
rect 1878 4748 1882 4752
rect 1886 4748 1890 4752
rect 1942 4748 1946 4752
rect 1966 4748 1970 4752
rect 2046 4748 2050 4752
rect 2070 4747 2074 4751
rect 2118 4748 2122 4752
rect 2142 4748 2146 4752
rect 2166 4748 2170 4752
rect 2214 4748 2218 4752
rect 2222 4748 2226 4752
rect 2278 4748 2282 4752
rect 2294 4748 2298 4752
rect 2334 4748 2338 4752
rect 2350 4748 2354 4752
rect 2414 4748 2418 4752
rect 2478 4748 2482 4752
rect 2542 4748 2546 4752
rect 2550 4748 2554 4752
rect 2606 4748 2610 4752
rect 2638 4748 2642 4752
rect 2718 4748 2722 4752
rect 2790 4748 2794 4752
rect 2878 4748 2882 4752
rect 2902 4748 2906 4752
rect 2926 4748 2930 4752
rect 2990 4748 2994 4752
rect 3070 4748 3074 4752
rect 3094 4748 3098 4752
rect 3102 4748 3106 4752
rect 3174 4747 3178 4751
rect 3206 4748 3210 4752
rect 3302 4747 3306 4751
rect 3414 4747 3418 4751
rect 3446 4748 3450 4752
rect 3518 4748 3522 4752
rect 3638 4748 3642 4752
rect 3686 4748 3690 4752
rect 3814 4758 3818 4762
rect 3862 4758 3866 4762
rect 3902 4758 3906 4762
rect 3974 4758 3978 4762
rect 4414 4758 4418 4762
rect 4510 4758 4514 4762
rect 4550 4758 4554 4762
rect 5006 4758 5010 4762
rect 5190 4758 5194 4762
rect 3726 4748 3730 4752
rect 3774 4748 3778 4752
rect 3846 4748 3850 4752
rect 3870 4748 3874 4752
rect 3942 4748 3946 4752
rect 3958 4748 3962 4752
rect 4038 4748 4042 4752
rect 4046 4748 4050 4752
rect 4094 4748 4098 4752
rect 4102 4748 4106 4752
rect 4134 4748 4138 4752
rect 4142 4748 4146 4752
rect 4150 4748 4154 4752
rect 4158 4748 4162 4752
rect 4182 4748 4186 4752
rect 4214 4748 4218 4752
rect 4294 4748 4298 4752
rect 4430 4748 4434 4752
rect 4454 4748 4458 4752
rect 4494 4748 4498 4752
rect 4566 4748 4570 4752
rect 4574 4748 4578 4752
rect 4638 4748 4642 4752
rect 4678 4748 4682 4752
rect 4710 4748 4714 4752
rect 4742 4748 4746 4752
rect 4758 4748 4762 4752
rect 4806 4748 4810 4752
rect 4910 4748 4914 4752
rect 4918 4748 4922 4752
rect 4998 4748 5002 4752
rect 5022 4748 5026 4752
rect 5102 4747 5106 4751
rect 5134 4748 5138 4752
rect 5166 4748 5170 4752
rect 5246 4748 5250 4752
rect 1678 4738 1682 4742
rect 1726 4738 1730 4742
rect 1830 4738 1834 4742
rect 1902 4738 1906 4742
rect 2126 4738 2130 4742
rect 2134 4738 2138 4742
rect 2206 4738 2210 4742
rect 2358 4738 2362 4742
rect 2422 4738 2426 4742
rect 2454 4738 2458 4742
rect 2614 4738 2618 4742
rect 2630 4738 2634 4742
rect 2742 4738 2746 4742
rect 2854 4738 2858 4742
rect 2870 4738 2874 4742
rect 2958 4738 2962 4742
rect 2982 4738 2986 4742
rect 3062 4738 3066 4742
rect 3158 4738 3162 4742
rect 3270 4738 3274 4742
rect 3470 4738 3474 4742
rect 3494 4738 3498 4742
rect 3542 4738 3546 4742
rect 3662 4738 3666 4742
rect 3678 4738 3682 4742
rect 3734 4738 3738 4742
rect 3766 4738 3770 4742
rect 3838 4738 3842 4742
rect 3878 4738 3882 4742
rect 3950 4738 3954 4742
rect 3998 4738 4002 4742
rect 4006 4738 4010 4742
rect 4086 4738 4090 4742
rect 4190 4738 4194 4742
rect 4318 4738 4322 4742
rect 4334 4738 4338 4742
rect 4398 4738 4402 4742
rect 4462 4738 4466 4742
rect 4486 4738 4490 4742
rect 4518 4738 4522 4742
rect 4630 4738 4634 4742
rect 4686 4738 4690 4742
rect 4750 4738 4754 4742
rect 4998 4738 5002 4742
rect 5030 4738 5034 4742
rect 5118 4738 5122 4742
rect 5134 4738 5138 4742
rect 5158 4738 5162 4742
rect 5222 4738 5226 4742
rect 5270 4738 5274 4742
rect 86 4728 90 4732
rect 630 4728 634 4732
rect 694 4728 698 4732
rect 902 4728 906 4732
rect 926 4728 930 4732
rect 958 4728 962 4732
rect 1094 4728 1098 4732
rect 1126 4728 1130 4732
rect 1158 4728 1162 4732
rect 1598 4728 1602 4732
rect 1606 4728 1610 4732
rect 1638 4728 1642 4732
rect 1678 4728 1682 4732
rect 1782 4728 1786 4732
rect 2182 4728 2186 4732
rect 2278 4728 2282 4732
rect 2438 4728 2442 4732
rect 2470 4728 2474 4732
rect 2558 4728 2562 4732
rect 2598 4728 2602 4732
rect 2854 4728 2858 4732
rect 2886 4728 2890 4732
rect 2902 4728 2906 4732
rect 2942 4728 2946 4732
rect 3302 4728 3306 4732
rect 3598 4728 3602 4732
rect 4062 4728 4066 4732
rect 4214 4728 4218 4732
rect 4230 4728 4234 4732
rect 4478 4728 4482 4732
rect 4702 4728 4706 4732
rect 4726 4728 4730 4732
rect 4974 4728 4978 4732
rect 38 4718 42 4722
rect 110 4718 114 4722
rect 206 4718 210 4722
rect 366 4718 370 4722
rect 446 4718 450 4722
rect 734 4718 738 4722
rect 854 4718 858 4722
rect 934 4718 938 4722
rect 1014 4718 1018 4722
rect 1086 4718 1090 4722
rect 1118 4718 1122 4722
rect 1222 4718 1226 4722
rect 1246 4718 1250 4722
rect 1550 4718 1554 4722
rect 1590 4718 1594 4722
rect 1998 4718 2002 4722
rect 2006 4718 2010 4722
rect 2102 4718 2106 4722
rect 2158 4718 2162 4722
rect 2230 4718 2234 4722
rect 2286 4718 2290 4722
rect 2390 4718 2394 4722
rect 2430 4718 2434 4722
rect 2534 4718 2538 4722
rect 2662 4718 2666 4722
rect 2846 4718 2850 4722
rect 2934 4718 2938 4722
rect 3110 4718 3114 4722
rect 3366 4718 3370 4722
rect 3574 4718 3578 4722
rect 3710 4718 3714 4722
rect 3830 4718 3834 4722
rect 3862 4718 3866 4722
rect 3886 4718 3890 4722
rect 3990 4718 3994 4722
rect 4078 4718 4082 4722
rect 4222 4718 4226 4722
rect 4238 4718 4242 4722
rect 4470 4718 4474 4722
rect 4510 4718 4514 4722
rect 4694 4718 4698 4722
rect 4766 4718 4770 4722
rect 4966 4718 4970 4722
rect 4982 4718 4986 4722
rect 5006 4718 5010 4722
rect 5038 4718 5042 4722
rect 850 4703 854 4707
rect 857 4703 861 4707
rect 1874 4703 1878 4707
rect 1881 4703 1885 4707
rect 2890 4703 2894 4707
rect 2897 4703 2901 4707
rect 3922 4703 3926 4707
rect 3929 4703 3933 4707
rect 4938 4703 4942 4707
rect 4945 4703 4949 4707
rect 94 4688 98 4692
rect 222 4688 226 4692
rect 238 4688 242 4692
rect 438 4688 442 4692
rect 590 4688 594 4692
rect 670 4688 674 4692
rect 686 4688 690 4692
rect 934 4688 938 4692
rect 958 4688 962 4692
rect 1182 4688 1186 4692
rect 1262 4688 1266 4692
rect 1358 4688 1362 4692
rect 1382 4688 1386 4692
rect 1438 4688 1442 4692
rect 1646 4688 1650 4692
rect 1742 4688 1746 4692
rect 1894 4688 1898 4692
rect 2022 4688 2026 4692
rect 2150 4688 2154 4692
rect 2270 4688 2274 4692
rect 2422 4688 2426 4692
rect 2454 4688 2458 4692
rect 2942 4688 2946 4692
rect 3182 4688 3186 4692
rect 3286 4688 3290 4692
rect 3518 4688 3522 4692
rect 3638 4688 3642 4692
rect 3734 4688 3738 4692
rect 4342 4688 4346 4692
rect 4422 4688 4426 4692
rect 4526 4688 4530 4692
rect 4630 4688 4634 4692
rect 4726 4688 4730 4692
rect 4910 4688 4914 4692
rect 5070 4688 5074 4692
rect 134 4678 138 4682
rect 158 4678 162 4682
rect 38 4668 42 4672
rect 126 4668 130 4672
rect 366 4678 370 4682
rect 422 4678 426 4682
rect 214 4668 218 4672
rect 286 4668 290 4672
rect 318 4668 322 4672
rect 710 4678 714 4682
rect 822 4678 826 4682
rect 878 4678 882 4682
rect 886 4678 890 4682
rect 966 4678 970 4682
rect 1102 4678 1106 4682
rect 1174 4678 1178 4682
rect 1318 4678 1322 4682
rect 486 4668 490 4672
rect 502 4668 506 4672
rect 606 4668 610 4672
rect 742 4668 746 4672
rect 766 4668 770 4672
rect 798 4668 802 4672
rect 830 4668 834 4672
rect 894 4668 898 4672
rect 950 4668 954 4672
rect 966 4668 970 4672
rect 998 4668 1002 4672
rect 1022 4668 1026 4672
rect 1134 4668 1138 4672
rect 1142 4668 1146 4672
rect 1206 4668 1210 4672
rect 1238 4668 1242 4672
rect 1246 4668 1250 4672
rect 1270 4668 1274 4672
rect 1310 4668 1314 4672
rect 1342 4678 1346 4682
rect 1366 4678 1370 4682
rect 1462 4678 1466 4682
rect 1566 4678 1570 4682
rect 1798 4678 1802 4682
rect 1990 4678 1994 4682
rect 2110 4678 2114 4682
rect 2118 4678 2122 4682
rect 1398 4668 1402 4672
rect 1454 4668 1458 4672
rect 1534 4668 1538 4672
rect 1662 4668 1666 4672
rect 1758 4668 1762 4672
rect 1774 4668 1778 4672
rect 1814 4668 1818 4672
rect 1918 4668 1922 4672
rect 1990 4668 1994 4672
rect 2062 4668 2066 4672
rect 2078 4668 2082 4672
rect 2094 4668 2098 4672
rect 2190 4668 2194 4672
rect 2286 4668 2290 4672
rect 2294 4668 2298 4672
rect 2310 4678 2314 4682
rect 2358 4678 2362 4682
rect 2438 4678 2442 4682
rect 2462 4678 2466 4682
rect 2542 4678 2546 4682
rect 2558 4678 2562 4682
rect 2494 4668 2498 4672
rect 2654 4678 2658 4682
rect 2934 4678 2938 4682
rect 2982 4678 2986 4682
rect 3150 4678 3154 4682
rect 3238 4678 3242 4682
rect 3318 4678 3322 4682
rect 3326 4678 3330 4682
rect 3350 4678 3354 4682
rect 3550 4678 3554 4682
rect 3670 4678 3674 4682
rect 3758 4678 3762 4682
rect 3798 4678 3802 4682
rect 3854 4678 3858 4682
rect 4054 4678 4058 4682
rect 4126 4678 4130 4682
rect 4366 4678 4370 4682
rect 2582 4668 2586 4672
rect 2606 4668 2610 4672
rect 2654 4668 2658 4672
rect 2702 4668 2706 4672
rect 2814 4668 2818 4672
rect 2862 4668 2866 4672
rect 3070 4668 3074 4672
rect 3142 4668 3146 4672
rect 3190 4668 3194 4672
rect 3230 4668 3234 4672
rect 3374 4668 3378 4672
rect 3406 4668 3410 4672
rect 3422 4668 3426 4672
rect 3462 4668 3466 4672
rect 3606 4668 3610 4672
rect 3614 4668 3618 4672
rect 3958 4668 3962 4672
rect 4014 4668 4018 4672
rect 4206 4668 4210 4672
rect 4518 4678 4522 4682
rect 4534 4678 4538 4682
rect 4686 4678 4690 4682
rect 4382 4668 4386 4672
rect 4390 4668 4394 4672
rect 4550 4668 4554 4672
rect 4574 4668 4578 4672
rect 4638 4668 4642 4672
rect 4854 4678 4858 4682
rect 4990 4678 4994 4682
rect 4710 4668 4714 4672
rect 4894 4668 4898 4672
rect 5046 4668 5050 4672
rect 5062 4668 5066 4672
rect 5086 4678 5090 4682
rect 5270 4678 5274 4682
rect 5102 4668 5106 4672
rect 5190 4668 5194 4672
rect 5262 4668 5266 4672
rect 46 4658 50 4662
rect 102 4658 106 4662
rect 150 4658 154 4662
rect 198 4658 202 4662
rect 214 4658 218 4662
rect 278 4658 282 4662
rect 334 4659 338 4663
rect 406 4658 410 4662
rect 526 4658 530 4662
rect 622 4658 626 4662
rect 654 4658 658 4662
rect 686 4658 690 4662
rect 758 4658 762 4662
rect 774 4658 778 4662
rect 830 4658 834 4662
rect 918 4658 922 4662
rect 942 4658 946 4662
rect 990 4658 994 4662
rect 1038 4658 1042 4662
rect 1070 4658 1074 4662
rect 1102 4658 1106 4662
rect 1110 4658 1114 4662
rect 1126 4658 1130 4662
rect 1158 4658 1162 4662
rect 1198 4658 1202 4662
rect 1230 4658 1234 4662
rect 1246 4658 1250 4662
rect 1278 4658 1282 4662
rect 1302 4658 1306 4662
rect 1318 4658 1322 4662
rect 1398 4658 1402 4662
rect 1414 4658 1418 4662
rect 1566 4659 1570 4663
rect 1598 4658 1602 4662
rect 1678 4659 1682 4663
rect 1710 4658 1714 4662
rect 1750 4658 1754 4662
rect 1782 4658 1786 4662
rect 1830 4659 1834 4663
rect 2006 4658 2010 4662
rect 2014 4658 2018 4662
rect 2038 4658 2042 4662
rect 2070 4658 2074 4662
rect 2086 4658 2090 4662
rect 2166 4658 2170 4662
rect 2174 4658 2178 4662
rect 2214 4658 2218 4662
rect 2278 4658 2282 4662
rect 2326 4658 2330 4662
rect 2366 4658 2370 4662
rect 2462 4658 2466 4662
rect 2486 4658 2490 4662
rect 2518 4658 2522 4662
rect 2534 4658 2538 4662
rect 2574 4658 2578 4662
rect 2590 4658 2594 4662
rect 2622 4659 2626 4663
rect 2726 4658 2730 4662
rect 2806 4658 2810 4662
rect 2838 4658 2842 4662
rect 2846 4658 2850 4662
rect 2870 4658 2874 4662
rect 2926 4658 2930 4662
rect 2950 4658 2954 4662
rect 2990 4658 2994 4662
rect 3102 4658 3106 4662
rect 3110 4658 3114 4662
rect 3118 4658 3122 4662
rect 3166 4658 3170 4662
rect 3198 4658 3202 4662
rect 3222 4658 3226 4662
rect 3254 4658 3258 4662
rect 3262 4658 3266 4662
rect 3270 4658 3274 4662
rect 3342 4658 3346 4662
rect 3366 4658 3370 4662
rect 3382 4658 3386 4662
rect 3398 4658 3402 4662
rect 3438 4658 3442 4662
rect 3470 4658 3474 4662
rect 3494 4658 3498 4662
rect 3502 4658 3506 4662
rect 3566 4658 3570 4662
rect 3622 4658 3626 4662
rect 3678 4658 3682 4662
rect 3742 4658 3746 4662
rect 3750 4658 3754 4662
rect 3822 4658 3826 4662
rect 3862 4658 3866 4662
rect 3990 4658 3994 4662
rect 3998 4658 4002 4662
rect 4006 4658 4010 4662
rect 4038 4658 4042 4662
rect 4110 4658 4114 4662
rect 4222 4659 4226 4663
rect 4278 4659 4282 4663
rect 4350 4658 4354 4662
rect 4406 4658 4410 4662
rect 4454 4658 4458 4662
rect 4478 4658 4482 4662
rect 4518 4658 4522 4662
rect 4566 4659 4570 4663
rect 4638 4658 4642 4662
rect 4670 4658 4674 4662
rect 4702 4658 4706 4662
rect 4718 4658 4722 4662
rect 4766 4658 4770 4662
rect 4782 4658 4786 4662
rect 4846 4658 4850 4662
rect 4870 4658 4874 4662
rect 4886 4658 4890 4662
rect 4902 4658 4906 4662
rect 4982 4658 4986 4662
rect 5038 4658 5042 4662
rect 5054 4658 5058 4662
rect 5102 4658 5106 4662
rect 5118 4658 5122 4662
rect 5142 4658 5146 4662
rect 5150 4658 5154 4662
rect 5166 4658 5170 4662
rect 5190 4658 5194 4662
rect 5246 4658 5250 4662
rect 102 4648 106 4652
rect 230 4648 234 4652
rect 262 4648 266 4652
rect 470 4648 474 4652
rect 590 4648 594 4652
rect 614 4648 618 4652
rect 646 4648 650 4652
rect 678 4648 682 4652
rect 718 4648 722 4652
rect 790 4648 794 4652
rect 822 4648 826 4652
rect 854 4648 858 4652
rect 934 4648 938 4652
rect 974 4648 978 4652
rect 1006 4648 1010 4652
rect 1030 4648 1034 4652
rect 1062 4648 1066 4652
rect 1206 4648 1210 4652
rect 1286 4648 1290 4652
rect 1406 4648 1410 4652
rect 2054 4648 2058 4652
rect 2854 4648 2858 4652
rect 3206 4648 3210 4652
rect 3334 4648 3338 4652
rect 3454 4648 3458 4652
rect 3486 4648 3490 4652
rect 3590 4648 3594 4652
rect 3638 4648 3642 4652
rect 4614 4648 4618 4652
rect 4662 4648 4666 4652
rect 5022 4648 5026 4652
rect 406 4638 410 4642
rect 614 4638 618 4642
rect 662 4638 666 4642
rect 694 4638 698 4642
rect 838 4638 842 4642
rect 1046 4638 1050 4642
rect 1078 4638 1082 4642
rect 1102 4638 1106 4642
rect 1414 4638 1418 4642
rect 1422 4638 1426 4642
rect 1878 4638 1882 4642
rect 3366 4638 3370 4642
rect 4030 4638 4034 4642
rect 622 4628 626 4632
rect 1014 4628 1018 4632
rect 182 4618 186 4622
rect 398 4618 402 4622
rect 582 4618 586 4622
rect 670 4618 674 4622
rect 702 4618 706 4622
rect 1038 4618 1042 4622
rect 1070 4618 1074 4622
rect 1230 4618 1234 4622
rect 1302 4618 1306 4622
rect 1478 4618 1482 4622
rect 1742 4618 1746 4622
rect 1894 4618 1898 4622
rect 1974 4618 1978 4622
rect 2110 4618 2114 4622
rect 2270 4618 2274 4622
rect 2478 4618 2482 4622
rect 2510 4618 2514 4622
rect 2686 4618 2690 4622
rect 2910 4618 2914 4622
rect 3046 4618 3050 4622
rect 3222 4618 3226 4622
rect 3254 4618 3258 4622
rect 3390 4618 3394 4622
rect 3438 4618 3442 4622
rect 3470 4618 3474 4622
rect 3566 4618 3570 4622
rect 3822 4618 3826 4622
rect 3934 4618 3938 4622
rect 4158 4618 4162 4622
rect 4646 4618 4650 4622
rect 4726 4618 4730 4622
rect 4830 4618 4834 4622
rect 5038 4618 5042 4622
rect 5206 4618 5210 4622
rect 330 4603 334 4607
rect 337 4603 341 4607
rect 1354 4603 1358 4607
rect 1361 4603 1365 4607
rect 2386 4603 2390 4607
rect 2393 4603 2397 4607
rect 3402 4603 3406 4607
rect 3409 4603 3413 4607
rect 4426 4603 4430 4607
rect 4433 4603 4437 4607
rect 94 4588 98 4592
rect 190 4588 194 4592
rect 214 4588 218 4592
rect 318 4588 322 4592
rect 622 4588 626 4592
rect 638 4588 642 4592
rect 902 4588 906 4592
rect 1278 4588 1282 4592
rect 1302 4588 1306 4592
rect 1422 4588 1426 4592
rect 1742 4588 1746 4592
rect 2518 4588 2522 4592
rect 2638 4588 2642 4592
rect 4046 4588 4050 4592
rect 4222 4588 4226 4592
rect 5142 4588 5146 4592
rect 582 4578 586 4582
rect 86 4568 90 4572
rect 126 4568 130 4572
rect 150 4568 154 4572
rect 182 4568 186 4572
rect 222 4568 226 4572
rect 246 4568 250 4572
rect 310 4568 314 4572
rect 590 4568 594 4572
rect 614 4568 618 4572
rect 1110 4568 1114 4572
rect 1118 4568 1122 4572
rect 1310 4568 1314 4572
rect 3294 4568 3298 4572
rect 3422 4568 3426 4572
rect 3614 4568 3618 4572
rect 4974 4568 4978 4572
rect 14 4558 18 4562
rect 54 4558 58 4562
rect 102 4558 106 4562
rect 110 4558 114 4562
rect 166 4558 170 4562
rect 198 4558 202 4562
rect 262 4558 266 4562
rect 294 4558 298 4562
rect 326 4558 330 4562
rect 470 4558 474 4562
rect 510 4558 514 4562
rect 606 4558 610 4562
rect 94 4548 98 4552
rect 126 4548 130 4552
rect 190 4548 194 4552
rect 214 4548 218 4552
rect 246 4548 250 4552
rect 278 4548 282 4552
rect 294 4548 298 4552
rect 310 4548 314 4552
rect 350 4548 354 4552
rect 374 4548 378 4552
rect 406 4548 410 4552
rect 446 4548 450 4552
rect 526 4548 530 4552
rect 550 4548 554 4552
rect 566 4548 570 4552
rect 598 4548 602 4552
rect 742 4558 746 4562
rect 918 4558 922 4562
rect 942 4558 946 4562
rect 1046 4558 1050 4562
rect 1126 4558 1130 4562
rect 1150 4558 1154 4562
rect 1158 4558 1162 4562
rect 1190 4558 1194 4562
rect 1222 4558 1226 4562
rect 1238 4558 1242 4562
rect 1294 4558 1298 4562
rect 1326 4558 1330 4562
rect 1414 4558 1418 4562
rect 1430 4558 1434 4562
rect 1614 4558 1618 4562
rect 1774 4558 1778 4562
rect 1782 4558 1786 4562
rect 1950 4558 1954 4562
rect 2390 4558 2394 4562
rect 2790 4558 2794 4562
rect 2878 4558 2882 4562
rect 638 4548 642 4552
rect 678 4548 682 4552
rect 686 4548 690 4552
rect 766 4548 770 4552
rect 806 4548 810 4552
rect 814 4548 818 4552
rect 902 4548 906 4552
rect 950 4548 954 4552
rect 1030 4548 1034 4552
rect 1118 4548 1122 4552
rect 1174 4548 1178 4552
rect 1182 4548 1186 4552
rect 1206 4548 1210 4552
rect 1262 4548 1266 4552
rect 1278 4548 1282 4552
rect 1318 4548 1322 4552
rect 1350 4548 1354 4552
rect 1374 4548 1378 4552
rect 1406 4548 1410 4552
rect 1438 4548 1442 4552
rect 1454 4548 1458 4552
rect 1470 4548 1474 4552
rect 1478 4548 1482 4552
rect 1502 4548 1506 4552
rect 1542 4547 1546 4551
rect 1574 4548 1578 4552
rect 1654 4547 1658 4551
rect 1726 4548 1730 4552
rect 1862 4548 1866 4552
rect 1926 4548 1930 4552
rect 1958 4548 1962 4552
rect 2038 4548 2042 4552
rect 2110 4548 2114 4552
rect 2134 4548 2138 4552
rect 2190 4548 2194 4552
rect 2222 4548 2226 4552
rect 2262 4548 2266 4552
rect 2286 4548 2290 4552
rect 2350 4548 2354 4552
rect 2358 4548 2362 4552
rect 2454 4548 2458 4552
rect 2502 4548 2506 4552
rect 2510 4548 2514 4552
rect 2534 4548 2538 4552
rect 2574 4547 2578 4551
rect 2606 4548 2610 4552
rect 2678 4548 2682 4552
rect 2686 4548 2690 4552
rect 2758 4548 2762 4552
rect 2766 4548 2770 4552
rect 2774 4548 2778 4552
rect 2798 4548 2802 4552
rect 2814 4548 2818 4552
rect 2846 4548 2850 4552
rect 2958 4548 2962 4552
rect 3014 4548 3018 4552
rect 3046 4547 3050 4551
rect 3150 4548 3154 4552
rect 3182 4547 3186 4551
rect 3214 4548 3218 4552
rect 3270 4548 3274 4552
rect 3278 4548 3282 4552
rect 3318 4558 3322 4562
rect 3510 4558 3514 4562
rect 3806 4558 3810 4562
rect 3822 4558 3826 4562
rect 3838 4558 3842 4562
rect 3870 4558 3874 4562
rect 4062 4558 4066 4562
rect 4078 4558 4082 4562
rect 4134 4558 4138 4562
rect 4206 4558 4210 4562
rect 4262 4558 4266 4562
rect 4630 4558 4634 4562
rect 4638 4558 4642 4562
rect 4694 4558 4698 4562
rect 4726 4558 4730 4562
rect 4998 4558 5002 4562
rect 5126 4558 5130 4562
rect 3318 4548 3322 4552
rect 3358 4547 3362 4551
rect 3446 4548 3450 4552
rect 3462 4548 3466 4552
rect 3478 4548 3482 4552
rect 3526 4548 3530 4552
rect 3574 4548 3578 4552
rect 3662 4548 3666 4552
rect 3686 4548 3690 4552
rect 3694 4548 3698 4552
rect 3702 4548 3706 4552
rect 3734 4548 3738 4552
rect 3774 4548 3778 4552
rect 3790 4548 3794 4552
rect 3822 4548 3826 4552
rect 3854 4548 3858 4552
rect 3870 4548 3874 4552
rect 3886 4548 3890 4552
rect 3902 4548 3906 4552
rect 3950 4548 3954 4552
rect 3982 4547 3986 4551
rect 4054 4548 4058 4552
rect 4086 4548 4090 4552
rect 4118 4548 4122 4552
rect 4150 4548 4154 4552
rect 4166 4548 4170 4552
rect 4198 4548 4202 4552
rect 4222 4548 4226 4552
rect 4262 4548 4266 4552
rect 4286 4548 4290 4552
rect 4374 4547 4378 4551
rect 4430 4548 4434 4552
rect 4454 4548 4458 4552
rect 4486 4548 4490 4552
rect 4502 4548 4506 4552
rect 4550 4548 4554 4552
rect 4614 4548 4618 4552
rect 4654 4548 4658 4552
rect 4686 4548 4690 4552
rect 4718 4548 4722 4552
rect 4734 4548 4738 4552
rect 4742 4548 4746 4552
rect 4774 4548 4778 4552
rect 4806 4548 4810 4552
rect 4814 4548 4818 4552
rect 4822 4548 4826 4552
rect 4854 4548 4858 4552
rect 4878 4548 4882 4552
rect 4910 4547 4914 4551
rect 5014 4548 5018 4552
rect 5054 4548 5058 4552
rect 5118 4548 5122 4552
rect 5142 4548 5146 4552
rect 5182 4548 5186 4552
rect 5206 4548 5210 4552
rect 5254 4548 5258 4552
rect 22 4538 26 4542
rect 30 4538 34 4542
rect 46 4538 50 4542
rect 70 4538 74 4542
rect 142 4538 146 4542
rect 238 4538 242 4542
rect 270 4538 274 4542
rect 382 4538 386 4542
rect 438 4538 442 4542
rect 470 4538 474 4542
rect 502 4538 506 4542
rect 518 4538 522 4542
rect 534 4538 538 4542
rect 542 4538 546 4542
rect 574 4538 578 4542
rect 614 4538 618 4542
rect 710 4538 714 4542
rect 758 4538 762 4542
rect 806 4538 810 4542
rect 830 4538 834 4542
rect 862 4538 866 4542
rect 926 4538 930 4542
rect 942 4538 946 4542
rect 958 4538 962 4542
rect 1022 4538 1026 4542
rect 1062 4538 1066 4542
rect 1078 4538 1082 4542
rect 1134 4538 1138 4542
rect 1182 4538 1186 4542
rect 1214 4538 1218 4542
rect 1246 4538 1250 4542
rect 1358 4538 1362 4542
rect 1430 4538 1434 4542
rect 1462 4538 1466 4542
rect 1502 4538 1506 4542
rect 1526 4538 1530 4542
rect 1662 4538 1666 4542
rect 1758 4538 1762 4542
rect 1790 4538 1794 4542
rect 1806 4538 1810 4542
rect 1878 4538 1882 4542
rect 1910 4538 1914 4542
rect 1934 4538 1938 4542
rect 2222 4538 2226 4542
rect 2326 4538 2330 4542
rect 2366 4538 2370 4542
rect 2470 4538 2474 4542
rect 2558 4538 2562 4542
rect 2806 4538 2810 4542
rect 2982 4538 2986 4542
rect 3030 4538 3034 4542
rect 3222 4538 3226 4542
rect 3230 4538 3234 4542
rect 3262 4538 3266 4542
rect 3326 4538 3330 4542
rect 3342 4538 3346 4542
rect 3470 4538 3474 4542
rect 3502 4538 3506 4542
rect 3534 4538 3538 4542
rect 3550 4538 3554 4542
rect 3598 4538 3602 4542
rect 3654 4538 3658 4542
rect 3710 4538 3714 4542
rect 3782 4538 3786 4542
rect 3814 4538 3818 4542
rect 3846 4538 3850 4542
rect 3878 4538 3882 4542
rect 3910 4538 3914 4542
rect 3926 4538 3930 4542
rect 3966 4538 3970 4542
rect 4054 4538 4058 4542
rect 4110 4538 4114 4542
rect 4142 4538 4146 4542
rect 4174 4538 4178 4542
rect 4230 4538 4234 4542
rect 4270 4538 4274 4542
rect 4286 4538 4290 4542
rect 4358 4538 4362 4542
rect 4494 4538 4498 4542
rect 4574 4538 4578 4542
rect 4590 4538 4594 4542
rect 4606 4538 4610 4542
rect 4694 4538 4698 4542
rect 4718 4538 4722 4542
rect 4758 4538 4762 4542
rect 4798 4538 4802 4542
rect 4846 4538 4850 4542
rect 4894 4538 4898 4542
rect 5022 4538 5026 4542
rect 5030 4538 5034 4542
rect 5078 4538 5082 4542
rect 5110 4538 5114 4542
rect 5158 4538 5162 4542
rect 5174 4538 5178 4542
rect 5190 4538 5194 4542
rect 5262 4538 5266 4542
rect 366 4528 370 4532
rect 398 4528 402 4532
rect 422 4528 426 4532
rect 430 4528 434 4532
rect 438 4528 442 4532
rect 462 4528 466 4532
rect 662 4528 666 4532
rect 702 4528 706 4532
rect 782 4528 786 4532
rect 822 4528 826 4532
rect 974 4528 978 4532
rect 990 4528 994 4532
rect 1070 4528 1074 4532
rect 1246 4528 1250 4532
rect 1382 4528 1386 4532
rect 1974 4528 1978 4532
rect 2174 4528 2178 4532
rect 2206 4528 2210 4532
rect 2382 4528 2386 4532
rect 2742 4528 2746 4532
rect 2862 4528 2866 4532
rect 2998 4528 3002 4532
rect 3246 4528 3250 4532
rect 3446 4528 3450 4532
rect 3670 4528 3674 4532
rect 3726 4528 3730 4532
rect 3734 4528 3738 4532
rect 3750 4528 3754 4532
rect 3806 4528 3810 4532
rect 3934 4528 3938 4532
rect 4102 4528 4106 4532
rect 4182 4528 4186 4532
rect 4198 4528 4202 4532
rect 4238 4528 4242 4532
rect 4254 4528 4258 4532
rect 4470 4528 4474 4532
rect 4670 4528 4674 4532
rect 4758 4528 4762 4532
rect 4862 4528 4866 4532
rect 5094 4528 5098 4532
rect 5158 4528 5162 4532
rect 5278 4528 5282 4532
rect 62 4518 66 4522
rect 358 4518 362 4522
rect 390 4518 394 4522
rect 414 4518 418 4522
rect 494 4518 498 4522
rect 566 4518 570 4522
rect 598 4518 602 4522
rect 630 4518 634 4522
rect 694 4518 698 4522
rect 798 4518 802 4522
rect 830 4518 834 4522
rect 942 4518 946 4522
rect 966 4518 970 4522
rect 1094 4518 1098 4522
rect 1150 4518 1154 4522
rect 1158 4518 1162 4522
rect 1230 4518 1234 4522
rect 1254 4518 1258 4522
rect 1334 4518 1338 4522
rect 1718 4518 1722 4522
rect 1742 4518 1746 4522
rect 1766 4518 1770 4522
rect 1814 4518 1818 4522
rect 2318 4518 2322 4522
rect 2406 4518 2410 4522
rect 2638 4518 2642 4522
rect 2646 4518 2650 4522
rect 2750 4518 2754 4522
rect 2830 4518 2834 4522
rect 3006 4518 3010 4522
rect 3110 4518 3114 4522
rect 3118 4518 3122 4522
rect 3478 4518 3482 4522
rect 3718 4518 3722 4522
rect 3766 4518 3770 4522
rect 3902 4518 3906 4522
rect 4094 4518 4098 4522
rect 4134 4518 4138 4522
rect 4166 4518 4170 4522
rect 4294 4518 4298 4522
rect 4414 4518 4418 4522
rect 4510 4518 4514 4522
rect 4630 4518 4634 4522
rect 4638 4518 4642 4522
rect 4790 4518 4794 4522
rect 4870 4518 4874 4522
rect 4990 4518 4994 4522
rect 5102 4518 5106 4522
rect 5166 4518 5170 4522
rect 5198 4518 5202 4522
rect 5214 4518 5218 4522
rect 850 4503 854 4507
rect 857 4503 861 4507
rect 1874 4503 1878 4507
rect 1881 4503 1885 4507
rect 2890 4503 2894 4507
rect 2897 4503 2901 4507
rect 3922 4503 3926 4507
rect 3929 4503 3933 4507
rect 4938 4503 4942 4507
rect 4945 4503 4949 4507
rect 22 4488 26 4492
rect 94 4488 98 4492
rect 158 4488 162 4492
rect 214 4488 218 4492
rect 310 4488 314 4492
rect 382 4488 386 4492
rect 870 4488 874 4492
rect 982 4488 986 4492
rect 1166 4488 1170 4492
rect 1222 4488 1226 4492
rect 1310 4488 1314 4492
rect 1382 4488 1386 4492
rect 1582 4488 1586 4492
rect 1638 4488 1642 4492
rect 1686 4488 1690 4492
rect 1838 4488 1842 4492
rect 2382 4488 2386 4492
rect 2614 4488 2618 4492
rect 2806 4488 2810 4492
rect 2886 4488 2890 4492
rect 3038 4488 3042 4492
rect 3678 4488 3682 4492
rect 3742 4488 3746 4492
rect 4374 4488 4378 4492
rect 4534 4488 4538 4492
rect 4646 4488 4650 4492
rect 4822 4488 4826 4492
rect 4998 4488 5002 4492
rect 5134 4488 5138 4492
rect 62 4478 66 4482
rect 142 4478 146 4482
rect 6 4468 10 4472
rect 30 4468 34 4472
rect 126 4468 130 4472
rect 182 4478 186 4482
rect 206 4478 210 4482
rect 342 4478 346 4482
rect 390 4478 394 4482
rect 510 4478 514 4482
rect 590 4478 594 4482
rect 782 4478 786 4482
rect 934 4478 938 4482
rect 974 4478 978 4482
rect 166 4468 170 4472
rect 214 4468 218 4472
rect 270 4468 274 4472
rect 286 4468 290 4472
rect 358 4468 362 4472
rect 438 4468 442 4472
rect 454 4468 458 4472
rect 558 4468 562 4472
rect 574 4468 578 4472
rect 582 4468 586 4472
rect 638 4468 642 4472
rect 670 4468 674 4472
rect 726 4468 730 4472
rect 774 4468 778 4472
rect 806 4468 810 4472
rect 822 4468 826 4472
rect 886 4468 890 4472
rect 990 4468 994 4472
rect 1046 4468 1050 4472
rect 1070 4478 1074 4482
rect 1134 4478 1138 4482
rect 1246 4478 1250 4482
rect 1262 4478 1266 4482
rect 1278 4478 1282 4482
rect 1318 4478 1322 4482
rect 1326 4478 1330 4482
rect 1486 4478 1490 4482
rect 1806 4478 1810 4482
rect 2310 4478 2314 4482
rect 2374 4478 2378 4482
rect 2646 4478 2650 4482
rect 2702 4478 2706 4482
rect 2734 4478 2738 4482
rect 3062 4478 3066 4482
rect 3078 4478 3082 4482
rect 1086 4468 1090 4472
rect 1142 4468 1146 4472
rect 1150 4468 1154 4472
rect 1166 4468 1170 4472
rect 1182 4468 1186 4472
rect 1214 4468 1218 4472
rect 1238 4468 1242 4472
rect 1286 4468 1290 4472
rect 1390 4468 1394 4472
rect 1446 4468 1450 4472
rect 1526 4468 1530 4472
rect 1614 4468 1618 4472
rect 1630 4468 1634 4472
rect 1670 4468 1674 4472
rect 1774 4468 1778 4472
rect 1782 4468 1786 4472
rect 1846 4468 1850 4472
rect 1910 4468 1914 4472
rect 2022 4468 2026 4472
rect 2046 4468 2050 4472
rect 2070 4468 2074 4472
rect 2110 4468 2114 4472
rect 2198 4468 2202 4472
rect 2238 4468 2242 4472
rect 2334 4468 2338 4472
rect 2422 4468 2426 4472
rect 2470 4468 2474 4472
rect 2718 4468 2722 4472
rect 2734 4468 2738 4472
rect 2790 4466 2794 4470
rect 2798 4468 2802 4472
rect 2830 4468 2834 4472
rect 3102 4478 3106 4482
rect 3150 4478 3154 4482
rect 3582 4478 3586 4482
rect 3734 4478 3738 4482
rect 3862 4478 3866 4482
rect 3910 4478 3914 4482
rect 3094 4468 3098 4472
rect 3118 4468 3122 4472
rect 3158 4468 3162 4472
rect 3182 4468 3186 4472
rect 3214 4468 3218 4472
rect 3334 4468 3338 4472
rect 3374 4468 3378 4472
rect 3382 4468 3386 4472
rect 3406 4468 3410 4472
rect 3422 4468 3426 4472
rect 3534 4468 3538 4472
rect 3542 4468 3546 4472
rect 3558 4468 3562 4472
rect 3598 4468 3602 4472
rect 3718 4468 3722 4472
rect 3822 4468 3826 4472
rect 3846 4468 3850 4472
rect 3870 4468 3874 4472
rect 3886 4468 3890 4472
rect 4254 4478 4258 4482
rect 4446 4478 4450 4482
rect 4478 4478 4482 4482
rect 4726 4478 4730 4482
rect 4830 4478 4834 4482
rect 4958 4478 4962 4482
rect 4990 4478 4994 4482
rect 5142 4478 5146 4482
rect 3958 4468 3962 4472
rect 4054 4468 4058 4472
rect 4190 4468 4194 4472
rect 4302 4468 4306 4472
rect 4318 4468 4322 4472
rect 4398 4468 4402 4472
rect 4462 4468 4466 4472
rect 4502 4468 4506 4472
rect 4518 4468 4522 4472
rect 4590 4468 4594 4472
rect 4686 4468 4690 4472
rect 4750 4468 4754 4472
rect 4790 4468 4794 4472
rect 4862 4468 4866 4472
rect 4934 4468 4938 4472
rect 4974 4468 4978 4472
rect 5006 4468 5010 4472
rect 5102 4468 5106 4472
rect 5126 4468 5130 4472
rect 5190 4468 5194 4472
rect 5278 4468 5282 4472
rect 38 4458 42 4462
rect 62 4458 66 4462
rect 78 4458 82 4462
rect 94 4458 98 4462
rect 118 4458 122 4462
rect 174 4458 178 4462
rect 222 4458 226 4462
rect 278 4458 282 4462
rect 310 4458 314 4462
rect 334 4458 338 4462
rect 366 4458 370 4462
rect 374 4458 378 4462
rect 398 4458 402 4462
rect 414 4458 418 4462
rect 430 4458 434 4462
rect 478 4458 482 4462
rect 494 4458 498 4462
rect 526 4458 530 4462
rect 550 4458 554 4462
rect 582 4458 586 4462
rect 630 4458 634 4462
rect 646 4458 650 4462
rect 694 4458 698 4462
rect 718 4458 722 4462
rect 766 4458 770 4462
rect 790 4458 794 4462
rect 830 4458 834 4462
rect 870 4458 874 4462
rect 886 4458 890 4462
rect 918 4458 922 4462
rect 950 4458 954 4462
rect 998 4458 1002 4462
rect 1038 4458 1042 4462
rect 1094 4458 1098 4462
rect 1110 4458 1114 4462
rect 1158 4458 1162 4462
rect 1182 4458 1186 4462
rect 1206 4458 1210 4462
rect 1262 4458 1266 4462
rect 1294 4458 1298 4462
rect 1302 4458 1306 4462
rect 1350 4458 1354 4462
rect 1438 4458 1442 4462
rect 1470 4458 1474 4462
rect 1518 4459 1522 4463
rect 1598 4458 1602 4462
rect 1606 4458 1610 4462
rect 1622 4458 1626 4462
rect 1654 4458 1658 4462
rect 1702 4458 1706 4462
rect 1822 4458 1826 4462
rect 1854 4458 1858 4462
rect 1870 4458 1874 4462
rect 1910 4458 1914 4462
rect 1998 4458 2002 4462
rect 2062 4458 2066 4462
rect 2078 4458 2082 4462
rect 2086 4458 2090 4462
rect 2118 4458 2122 4462
rect 2134 4458 2138 4462
rect 2190 4458 2194 4462
rect 2302 4458 2306 4462
rect 2334 4458 2338 4462
rect 2358 4458 2362 4462
rect 2366 4458 2370 4462
rect 2390 4458 2394 4462
rect 2406 4458 2410 4462
rect 2462 4458 2466 4462
rect 2526 4458 2530 4462
rect 2550 4458 2554 4462
rect 2590 4458 2594 4462
rect 2598 4458 2602 4462
rect 2662 4458 2666 4462
rect 2686 4458 2690 4462
rect 2702 4458 2706 4462
rect 2750 4458 2754 4462
rect 2822 4458 2826 4462
rect 2838 4458 2842 4462
rect 2846 4458 2850 4462
rect 2870 4458 2874 4462
rect 2878 4458 2882 4462
rect 2958 4458 2962 4462
rect 2974 4458 2978 4462
rect 3022 4458 3026 4462
rect 3046 4458 3050 4462
rect 3054 4458 3058 4462
rect 3078 4458 3082 4462
rect 3126 4458 3130 4462
rect 3134 4458 3138 4462
rect 3150 4458 3154 4462
rect 3190 4458 3194 4462
rect 3206 4458 3210 4462
rect 3222 4458 3226 4462
rect 3238 4458 3242 4462
rect 3310 4458 3314 4462
rect 3350 4458 3354 4462
rect 3358 4458 3362 4462
rect 3366 4458 3370 4462
rect 3398 4458 3402 4462
rect 3502 4458 3506 4462
rect 3526 4458 3530 4462
rect 3566 4458 3570 4462
rect 3614 4459 3618 4463
rect 3702 4458 3706 4462
rect 3710 4458 3714 4462
rect 3798 4458 3802 4462
rect 3838 4458 3842 4462
rect 3878 4458 3882 4462
rect 3950 4458 3954 4462
rect 4030 4458 4034 4462
rect 4070 4458 4074 4462
rect 4094 4458 4098 4462
rect 4102 4458 4106 4462
rect 4150 4458 4154 4462
rect 4278 4458 4282 4462
rect 4326 4458 4330 4462
rect 4350 4458 4354 4462
rect 4358 4458 4362 4462
rect 4382 4458 4386 4462
rect 4390 4458 4394 4462
rect 4478 4458 4482 4462
rect 4494 4458 4498 4462
rect 4526 4458 4530 4462
rect 4574 4458 4578 4462
rect 4630 4458 4634 4462
rect 4654 4458 4658 4462
rect 4742 4458 4746 4462
rect 4798 4458 4802 4462
rect 4846 4458 4850 4462
rect 4854 4458 4858 4462
rect 4942 4458 4946 4462
rect 4982 4458 4986 4462
rect 5014 4458 5018 4462
rect 5078 4458 5082 4462
rect 5118 4458 5122 4462
rect 5150 4458 5154 4462
rect 5158 4458 5162 4462
rect 5182 4458 5186 4462
rect 5230 4458 5234 4462
rect 5254 4458 5258 4462
rect 22 4448 26 4452
rect 54 4448 58 4452
rect 86 4448 90 4452
rect 262 4448 266 4452
rect 318 4448 322 4452
rect 422 4448 426 4452
rect 462 4448 466 4452
rect 518 4448 522 4452
rect 558 4448 562 4452
rect 614 4448 618 4452
rect 646 4448 650 4452
rect 678 4448 682 4452
rect 702 4448 706 4452
rect 822 4448 826 4452
rect 878 4448 882 4452
rect 894 4448 898 4452
rect 942 4448 946 4452
rect 1102 4448 1106 4452
rect 1166 4448 1170 4452
rect 1190 4448 1194 4452
rect 1222 4448 1226 4452
rect 1254 4448 1258 4452
rect 1374 4448 1378 4452
rect 1462 4448 1466 4452
rect 1590 4448 1594 4452
rect 1782 4448 1786 4452
rect 1798 4448 1802 4452
rect 2014 4448 2018 4452
rect 2038 4448 2042 4452
rect 2446 4448 2450 4452
rect 2766 4448 2770 4452
rect 2806 4448 2810 4452
rect 3174 4448 3178 4452
rect 3190 4448 3194 4452
rect 3222 4448 3226 4452
rect 3382 4448 3386 4452
rect 3734 4448 3738 4452
rect 3894 4448 3898 4452
rect 4326 4448 4330 4452
rect 4342 4448 4346 4452
rect 4662 4448 4666 4452
rect 4814 4448 4818 4452
rect 4838 4448 4842 4452
rect 102 4438 106 4442
rect 302 4438 306 4442
rect 406 4438 410 4442
rect 534 4438 538 4442
rect 862 4438 866 4442
rect 958 4438 962 4442
rect 1110 4438 1114 4442
rect 1422 4438 1426 4442
rect 2158 4438 2162 4442
rect 3078 4438 3082 4442
rect 3094 4438 3098 4442
rect 3254 4438 3258 4442
rect 5022 4438 5026 4442
rect 2734 4428 2738 4432
rect 78 4418 82 4422
rect 526 4418 530 4422
rect 742 4418 746 4422
rect 950 4418 954 4422
rect 1110 4418 1114 4422
rect 1326 4418 1330 4422
rect 1718 4418 1722 4422
rect 1966 4418 1970 4422
rect 1998 4418 2002 4422
rect 2438 4418 2442 4422
rect 2478 4418 2482 4422
rect 2662 4418 2666 4422
rect 2686 4418 2690 4422
rect 2750 4418 2754 4422
rect 2774 4418 2778 4422
rect 3102 4418 3106 4422
rect 3166 4418 3170 4422
rect 3486 4418 3490 4422
rect 3694 4418 3698 4422
rect 3862 4418 3866 4422
rect 4022 4418 4026 4422
rect 4046 4418 4050 4422
rect 4086 4418 4090 4422
rect 4110 4418 4114 4422
rect 4206 4418 4210 4422
rect 4406 4418 4410 4422
rect 4646 4418 4650 4422
rect 4798 4418 4802 4422
rect 4878 4418 4882 4422
rect 5198 4418 5202 4422
rect 330 4403 334 4407
rect 337 4403 341 4407
rect 1354 4403 1358 4407
rect 1361 4403 1365 4407
rect 2386 4403 2390 4407
rect 2393 4403 2397 4407
rect 3402 4403 3406 4407
rect 3409 4403 3413 4407
rect 4426 4403 4430 4407
rect 4433 4403 4437 4407
rect 38 4388 42 4392
rect 110 4388 114 4392
rect 190 4388 194 4392
rect 246 4388 250 4392
rect 278 4388 282 4392
rect 430 4388 434 4392
rect 550 4388 554 4392
rect 686 4388 690 4392
rect 838 4388 842 4392
rect 862 4388 866 4392
rect 934 4388 938 4392
rect 1102 4388 1106 4392
rect 1910 4388 1914 4392
rect 2550 4388 2554 4392
rect 2854 4388 2858 4392
rect 3854 4388 3858 4392
rect 3950 4388 3954 4392
rect 4094 4388 4098 4392
rect 4158 4388 4162 4392
rect 4726 4388 4730 4392
rect 526 4378 530 4382
rect 22 4368 26 4372
rect 78 4368 82 4372
rect 254 4368 258 4372
rect 286 4368 290 4372
rect 806 4368 810 4372
rect 926 4368 930 4372
rect 966 4368 970 4372
rect 1110 4368 1114 4372
rect 1150 4368 1154 4372
rect 1174 4368 1178 4372
rect 2574 4378 2578 4382
rect 3134 4378 3138 4382
rect 1958 4368 1962 4372
rect 2958 4368 2962 4372
rect 3382 4368 3386 4372
rect 4198 4368 4202 4372
rect 6 4358 10 4362
rect 118 4358 122 4362
rect 198 4358 202 4362
rect 238 4358 242 4362
rect 270 4358 274 4362
rect 318 4358 322 4362
rect 382 4358 386 4362
rect 494 4358 498 4362
rect 566 4358 570 4362
rect 582 4358 586 4362
rect 614 4358 618 4362
rect 646 4358 650 4362
rect 750 4358 754 4362
rect 790 4358 794 4362
rect 942 4358 946 4362
rect 950 4358 954 4362
rect 1078 4358 1082 4362
rect 1134 4358 1138 4362
rect 1190 4358 1194 4362
rect 1222 4358 1226 4362
rect 1590 4358 1594 4362
rect 1622 4358 1626 4362
rect 1854 4358 1858 4362
rect 1926 4358 1930 4362
rect 1942 4358 1946 4362
rect 2158 4358 2162 4362
rect 2238 4358 2242 4362
rect 2462 4358 2466 4362
rect 2494 4358 2498 4362
rect 2670 4358 2674 4362
rect 2686 4358 2690 4362
rect 2702 4358 2706 4362
rect 2758 4358 2762 4362
rect 3166 4358 3170 4362
rect 3366 4358 3370 4362
rect 3414 4358 3418 4362
rect 3542 4358 3546 4362
rect 3558 4358 3562 4362
rect 3782 4358 3786 4362
rect 3798 4358 3802 4362
rect 3830 4358 3834 4362
rect 3886 4358 3890 4362
rect 3982 4358 3986 4362
rect 4038 4358 4042 4362
rect 4646 4358 4650 4362
rect 4766 4358 4770 4362
rect 5046 4358 5050 4362
rect 5174 4358 5178 4362
rect 94 4348 98 4352
rect 174 4348 178 4352
rect 206 4348 210 4352
rect 246 4348 250 4352
rect 278 4348 282 4352
rect 342 4348 346 4352
rect 358 4348 362 4352
rect 374 4348 378 4352
rect 398 4348 402 4352
rect 470 4348 474 4352
rect 518 4348 522 4352
rect 558 4348 562 4352
rect 598 4348 602 4352
rect 614 4348 618 4352
rect 638 4348 642 4352
rect 662 4348 666 4352
rect 702 4348 706 4352
rect 734 4348 738 4352
rect 782 4348 786 4352
rect 806 4348 810 4352
rect 886 4348 890 4352
rect 934 4348 938 4352
rect 958 4348 962 4352
rect 1006 4348 1010 4352
rect 1038 4348 1042 4352
rect 1118 4348 1122 4352
rect 1142 4348 1146 4352
rect 1182 4348 1186 4352
rect 1310 4348 1314 4352
rect 1326 4348 1330 4352
rect 1382 4348 1386 4352
rect 22 4338 26 4342
rect 30 4338 34 4342
rect 102 4338 106 4342
rect 126 4338 130 4342
rect 134 4340 138 4344
rect 1414 4348 1418 4352
rect 1470 4348 1474 4352
rect 1494 4348 1498 4352
rect 1534 4348 1538 4352
rect 1574 4348 1578 4352
rect 1606 4348 1610 4352
rect 1622 4348 1626 4352
rect 1654 4347 1658 4351
rect 1686 4348 1690 4352
rect 1726 4348 1730 4352
rect 1742 4348 1746 4352
rect 1782 4347 1786 4351
rect 1862 4348 1866 4352
rect 1870 4348 1874 4352
rect 1894 4348 1898 4352
rect 1926 4348 1930 4352
rect 1990 4347 1994 4351
rect 2094 4348 2098 4352
rect 2110 4348 2114 4352
rect 2174 4348 2178 4352
rect 2198 4348 2202 4352
rect 2222 4348 2226 4352
rect 2230 4348 2234 4352
rect 2286 4348 2290 4352
rect 2390 4348 2394 4352
rect 2414 4348 2418 4352
rect 2422 4348 2426 4352
rect 2454 4348 2458 4352
rect 2478 4348 2482 4352
rect 2510 4348 2514 4352
rect 2534 4348 2538 4352
rect 2558 4348 2562 4352
rect 2566 4348 2570 4352
rect 2606 4348 2610 4352
rect 2638 4347 2642 4351
rect 2702 4348 2706 4352
rect 2710 4348 2714 4352
rect 2718 4348 2722 4352
rect 2742 4348 2746 4352
rect 2774 4348 2778 4352
rect 2790 4348 2794 4352
rect 2806 4348 2810 4352
rect 2838 4348 2842 4352
rect 2934 4348 2938 4352
rect 3014 4348 3018 4352
rect 3030 4348 3034 4352
rect 3038 4348 3042 4352
rect 3070 4347 3074 4351
rect 3150 4348 3154 4352
rect 3238 4347 3242 4351
rect 3334 4347 3338 4351
rect 3382 4348 3386 4352
rect 3406 4348 3410 4352
rect 3430 4348 3434 4352
rect 3526 4348 3530 4352
rect 3542 4348 3546 4352
rect 3558 4348 3562 4352
rect 3614 4348 3618 4352
rect 3638 4348 3642 4352
rect 3710 4348 3714 4352
rect 3782 4348 3786 4352
rect 3814 4348 3818 4352
rect 3838 4348 3842 4352
rect 3894 4348 3898 4352
rect 3934 4348 3938 4352
rect 3942 4348 3946 4352
rect 3966 4348 3970 4352
rect 3998 4348 4002 4352
rect 4022 4348 4026 4352
rect 4030 4348 4034 4352
rect 4062 4348 4066 4352
rect 4070 4348 4074 4352
rect 4078 4348 4082 4352
rect 4102 4348 4106 4352
rect 4126 4348 4130 4352
rect 4134 4348 4138 4352
rect 4142 4348 4146 4352
rect 4174 4348 4178 4352
rect 4206 4348 4210 4352
rect 158 4338 162 4342
rect 214 4338 218 4342
rect 302 4338 306 4342
rect 334 4338 338 4342
rect 350 4338 354 4342
rect 366 4338 370 4342
rect 406 4338 410 4342
rect 414 4338 418 4342
rect 462 4338 466 4342
rect 470 4338 474 4342
rect 518 4338 522 4342
rect 534 4338 538 4342
rect 566 4338 570 4342
rect 590 4338 594 4342
rect 670 4338 674 4342
rect 678 4338 682 4342
rect 726 4338 730 4342
rect 814 4338 818 4342
rect 822 4338 826 4342
rect 838 4338 842 4342
rect 894 4338 898 4342
rect 1014 4338 1018 4342
rect 1030 4338 1034 4342
rect 1094 4338 1098 4342
rect 1246 4338 1250 4342
rect 1390 4338 1394 4342
rect 1406 4338 1410 4342
rect 1518 4338 1522 4342
rect 1542 4338 1546 4342
rect 1566 4338 1570 4342
rect 1582 4338 1586 4342
rect 1598 4338 1602 4342
rect 1750 4338 1754 4342
rect 1766 4338 1770 4342
rect 1814 4338 1818 4342
rect 1878 4338 1882 4342
rect 1934 4338 1938 4342
rect 2182 4338 2186 4342
rect 2190 4338 2194 4342
rect 2262 4338 2266 4342
rect 2374 4338 2378 4342
rect 2446 4338 2450 4342
rect 2486 4338 2490 4342
rect 2518 4338 2522 4342
rect 2694 4338 2698 4342
rect 2726 4338 2730 4342
rect 2734 4338 2738 4342
rect 2766 4338 2770 4342
rect 2782 4338 2786 4342
rect 2798 4338 2802 4342
rect 2814 4338 2818 4342
rect 2894 4338 2898 4342
rect 3054 4338 3058 4342
rect 3142 4338 3146 4342
rect 3214 4338 3218 4342
rect 3254 4338 3258 4342
rect 3302 4338 3306 4342
rect 3350 4338 3354 4342
rect 3390 4338 3394 4342
rect 3438 4338 3442 4342
rect 3446 4338 3450 4342
rect 3510 4338 3514 4342
rect 3518 4338 3522 4342
rect 4238 4348 4242 4352
rect 4286 4347 4290 4351
rect 4374 4348 4378 4352
rect 4390 4348 4394 4352
rect 4414 4348 4418 4352
rect 4486 4348 4490 4352
rect 4590 4347 4594 4351
rect 4630 4348 4634 4352
rect 4670 4348 4674 4352
rect 4702 4348 4706 4352
rect 4710 4348 4714 4352
rect 4750 4348 4754 4352
rect 4814 4348 4818 4352
rect 4870 4348 4874 4352
rect 4878 4348 4882 4352
rect 4902 4348 4906 4352
rect 4910 4348 4914 4352
rect 4926 4348 4930 4352
rect 5006 4348 5010 4352
rect 5062 4348 5066 4352
rect 5110 4348 5114 4352
rect 5118 4348 5122 4352
rect 5190 4348 5194 4352
rect 5238 4348 5242 4352
rect 3550 4338 3554 4342
rect 3774 4338 3778 4342
rect 3806 4338 3810 4342
rect 3822 4338 3826 4342
rect 3862 4338 3866 4342
rect 3870 4338 3874 4342
rect 4006 4338 4010 4342
rect 4014 4338 4018 4342
rect 4126 4338 4130 4342
rect 4182 4338 4186 4342
rect 4214 4338 4218 4342
rect 4230 4338 4234 4342
rect 4302 4338 4306 4342
rect 4398 4338 4402 4342
rect 4510 4338 4514 4342
rect 158 4328 162 4332
rect 230 4328 234 4332
rect 486 4328 490 4332
rect 542 4328 546 4332
rect 622 4328 626 4332
rect 686 4328 690 4332
rect 718 4328 722 4332
rect 886 4328 890 4332
rect 902 4328 906 4332
rect 958 4328 962 4332
rect 982 4328 986 4332
rect 1014 4328 1018 4332
rect 1038 4328 1042 4332
rect 1262 4328 1266 4332
rect 1558 4328 1562 4332
rect 1990 4328 1994 4332
rect 2238 4328 2242 4332
rect 2430 4328 2434 4332
rect 2638 4328 2642 4332
rect 2758 4328 2762 4332
rect 2830 4328 2834 4332
rect 2982 4328 2986 4332
rect 3646 4328 3650 4332
rect 3910 4328 3914 4332
rect 4046 4328 4050 4332
rect 4062 4328 4066 4332
rect 4622 4338 4626 4342
rect 4694 4338 4698 4342
rect 4734 4338 4738 4342
rect 4758 4338 4762 4342
rect 4854 4338 4858 4342
rect 5030 4338 5034 4342
rect 5070 4338 5074 4342
rect 5198 4338 5202 4342
rect 5246 4338 5250 4342
rect 4254 4328 4258 4332
rect 4358 4328 4362 4332
rect 4558 4328 4562 4332
rect 4590 4328 4594 4332
rect 4654 4328 4658 4332
rect 5278 4328 5282 4332
rect 382 4318 386 4322
rect 494 4318 498 4322
rect 550 4318 554 4322
rect 630 4318 634 4322
rect 646 4318 650 4322
rect 710 4318 714 4322
rect 750 4318 754 4322
rect 766 4318 770 4322
rect 990 4318 994 4322
rect 1086 4318 1090 4322
rect 1198 4318 1202 4322
rect 1358 4318 1362 4322
rect 1438 4318 1442 4322
rect 1550 4318 1554 4322
rect 1718 4318 1722 4322
rect 1846 4318 1850 4322
rect 2054 4318 2058 4322
rect 2150 4318 2154 4322
rect 2158 4318 2162 4322
rect 2438 4318 2442 4322
rect 2462 4318 2466 4322
rect 2494 4318 2498 4322
rect 2822 4318 2826 4322
rect 2974 4318 2978 4322
rect 3166 4318 3170 4322
rect 3174 4318 3178 4322
rect 3270 4318 3274 4322
rect 3582 4318 3586 4322
rect 3766 4318 3770 4322
rect 3878 4318 3882 4322
rect 3902 4318 3906 4322
rect 3982 4318 3986 4322
rect 4190 4318 4194 4322
rect 4350 4318 4354 4322
rect 4430 4318 4434 4322
rect 4526 4318 4530 4322
rect 4646 4318 4650 4322
rect 4686 4318 4690 4322
rect 4774 4318 4778 4322
rect 5046 4318 5050 4322
rect 5078 4318 5082 4322
rect 5174 4318 5178 4322
rect 850 4303 854 4307
rect 857 4303 861 4307
rect 1874 4303 1878 4307
rect 1881 4303 1885 4307
rect 2890 4303 2894 4307
rect 2897 4303 2901 4307
rect 3922 4303 3926 4307
rect 3929 4303 3933 4307
rect 4938 4303 4942 4307
rect 4945 4303 4949 4307
rect 6 4288 10 4292
rect 166 4288 170 4292
rect 278 4288 282 4292
rect 350 4288 354 4292
rect 510 4288 514 4292
rect 526 4288 530 4292
rect 598 4288 602 4292
rect 718 4288 722 4292
rect 774 4288 778 4292
rect 790 4288 794 4292
rect 878 4288 882 4292
rect 902 4288 906 4292
rect 958 4288 962 4292
rect 1030 4288 1034 4292
rect 1134 4288 1138 4292
rect 1174 4288 1178 4292
rect 1310 4288 1314 4292
rect 1606 4288 1610 4292
rect 1662 4288 1666 4292
rect 1758 4288 1762 4292
rect 1854 4288 1858 4292
rect 2022 4288 2026 4292
rect 2062 4288 2066 4292
rect 2086 4288 2090 4292
rect 2118 4288 2122 4292
rect 2318 4288 2322 4292
rect 2550 4288 2554 4292
rect 2766 4288 2770 4292
rect 2790 4288 2794 4292
rect 2934 4288 2938 4292
rect 3134 4288 3138 4292
rect 3254 4288 3258 4292
rect 3542 4288 3546 4292
rect 3966 4288 3970 4292
rect 4134 4288 4138 4292
rect 4606 4288 4610 4292
rect 4646 4288 4650 4292
rect 4766 4288 4770 4292
rect 4806 4288 4810 4292
rect 4862 4288 4866 4292
rect 5118 4288 5122 4292
rect 5190 4288 5194 4292
rect 5206 4288 5210 4292
rect 142 4278 146 4282
rect 206 4278 210 4282
rect 406 4278 410 4282
rect 422 4278 426 4282
rect 430 4278 434 4282
rect 518 4278 522 4282
rect 574 4278 578 4282
rect 590 4278 594 4282
rect 646 4278 650 4282
rect 926 4278 930 4282
rect 46 4268 50 4272
rect 86 4268 90 4272
rect 102 4268 106 4272
rect 150 4268 154 4272
rect 222 4268 226 4272
rect 254 4268 258 4272
rect 302 4268 306 4272
rect 310 4268 314 4272
rect 358 4268 362 4272
rect 374 4268 378 4272
rect 390 4268 394 4272
rect 454 4268 458 4272
rect 486 4268 490 4272
rect 534 4268 538 4272
rect 566 4268 570 4272
rect 606 4268 610 4272
rect 662 4268 666 4272
rect 686 4268 690 4272
rect 694 4268 698 4272
rect 702 4268 706 4272
rect 742 4268 746 4272
rect 750 4268 754 4272
rect 798 4268 802 4272
rect 854 4268 858 4272
rect 918 4268 922 4272
rect 1038 4278 1042 4282
rect 1054 4278 1058 4282
rect 1102 4278 1106 4282
rect 1182 4278 1186 4282
rect 1342 4278 1346 4282
rect 1414 4278 1418 4282
rect 1438 4278 1442 4282
rect 1670 4278 1674 4282
rect 1710 4278 1714 4282
rect 1902 4278 1906 4282
rect 2054 4278 2058 4282
rect 2094 4278 2098 4282
rect 2214 4278 2218 4282
rect 2798 4278 2802 4282
rect 2870 4278 2874 4282
rect 2974 4278 2978 4282
rect 3222 4278 3226 4282
rect 3302 4278 3306 4282
rect 3534 4278 3538 4282
rect 4062 4278 4066 4282
rect 4310 4278 4314 4282
rect 4334 4278 4338 4282
rect 4414 4278 4418 4282
rect 4526 4278 4530 4282
rect 982 4268 986 4272
rect 1030 4268 1034 4272
rect 1142 4268 1146 4272
rect 1150 4268 1154 4272
rect 1190 4268 1194 4272
rect 1302 4268 1306 4272
rect 1398 4268 1402 4272
rect 1422 4268 1426 4272
rect 1446 4268 1450 4272
rect 1510 4268 1514 4272
rect 1526 4268 1530 4272
rect 1614 4268 1618 4272
rect 1654 4268 1658 4272
rect 1702 4268 1706 4272
rect 1734 4268 1738 4272
rect 1766 4268 1770 4272
rect 1822 4268 1826 4272
rect 1830 4268 1834 4272
rect 1998 4268 2002 4272
rect 2222 4268 2226 4272
rect 2262 4268 2266 4272
rect 2326 4268 2330 4272
rect 2422 4268 2426 4272
rect 2454 4268 2458 4272
rect 2462 4268 2466 4272
rect 2494 4268 2498 4272
rect 2518 4268 2522 4272
rect 2542 4268 2546 4272
rect 2638 4268 2642 4272
rect 2774 4268 2778 4272
rect 2798 4268 2802 4272
rect 2870 4268 2874 4272
rect 2918 4268 2922 4272
rect 2982 4268 2986 4272
rect 62 4258 66 4262
rect 118 4258 122 4262
rect 222 4258 226 4262
rect 318 4258 322 4262
rect 366 4258 370 4262
rect 438 4258 442 4262
rect 462 4258 466 4262
rect 478 4258 482 4262
rect 494 4258 498 4262
rect 590 4258 594 4262
rect 614 4258 618 4262
rect 630 4258 634 4262
rect 670 4258 674 4262
rect 678 4258 682 4262
rect 710 4258 714 4262
rect 734 4258 738 4262
rect 750 4258 754 4262
rect 814 4258 818 4262
rect 838 4258 842 4262
rect 878 4258 882 4262
rect 950 4258 954 4262
rect 974 4258 978 4262
rect 1022 4258 1026 4262
rect 1070 4258 1074 4262
rect 1078 4258 1082 4262
rect 1102 4258 1106 4262
rect 1118 4258 1122 4262
rect 1158 4258 1162 4262
rect 1246 4258 1250 4262
rect 1254 4258 1258 4262
rect 1294 4258 1298 4262
rect 1326 4258 1330 4262
rect 1366 4258 1370 4262
rect 1414 4258 1418 4262
rect 1422 4258 1426 4262
rect 1454 4258 1458 4262
rect 1486 4258 1490 4262
rect 1502 4258 1506 4262
rect 1542 4259 1546 4263
rect 1622 4258 1626 4262
rect 1646 4258 1650 4262
rect 1710 4258 1714 4262
rect 1726 4258 1730 4262
rect 1742 4258 1746 4262
rect 1774 4258 1778 4262
rect 1814 4258 1818 4262
rect 1838 4258 1842 4262
rect 1918 4258 1922 4262
rect 1990 4258 1994 4262
rect 2014 4258 2018 4262
rect 2038 4258 2042 4262
rect 2046 4258 2050 4262
rect 2070 4258 2074 4262
rect 2102 4258 2106 4262
rect 2134 4258 2138 4262
rect 2142 4258 2146 4262
rect 2166 4258 2170 4262
rect 2174 4258 2178 4262
rect 2198 4258 2202 4262
rect 2254 4259 2258 4263
rect 2334 4258 2338 4262
rect 2366 4258 2370 4262
rect 3014 4268 3018 4272
rect 3054 4268 3058 4272
rect 3206 4268 3210 4272
rect 3262 4268 3266 4272
rect 3390 4268 3394 4272
rect 3502 4268 3506 4272
rect 3582 4268 3586 4272
rect 3622 4268 3626 4272
rect 3662 4268 3666 4272
rect 3694 4268 3698 4272
rect 3726 4268 3730 4272
rect 3758 4268 3762 4272
rect 3782 4268 3786 4272
rect 3790 4268 3794 4272
rect 3846 4268 3850 4272
rect 4046 4268 4050 4272
rect 4078 4268 4082 4272
rect 4158 4268 4162 4272
rect 4214 4268 4218 4272
rect 4246 4268 4250 4272
rect 4254 4268 4258 4272
rect 4286 4268 4290 4272
rect 4406 4268 4410 4272
rect 4518 4268 4522 4272
rect 4582 4268 4586 4272
rect 4598 4268 4602 4272
rect 4622 4278 4626 4282
rect 4790 4278 4794 4282
rect 4958 4278 4962 4282
rect 5078 4278 5082 4282
rect 5198 4278 5202 4282
rect 4726 4268 4730 4272
rect 4790 4268 4794 4272
rect 4830 4268 4834 4272
rect 4974 4268 4978 4272
rect 5014 4268 5018 4272
rect 5054 4268 5058 4272
rect 5126 4268 5130 4272
rect 5142 4268 5146 4272
rect 5182 4268 5186 4272
rect 2438 4258 2442 4262
rect 2470 4258 2474 4262
rect 2534 4258 2538 4262
rect 2566 4258 2570 4262
rect 2638 4258 2642 4262
rect 2710 4258 2714 4262
rect 2774 4258 2778 4262
rect 2814 4258 2818 4262
rect 2862 4258 2866 4262
rect 2910 4258 2914 4262
rect 2950 4258 2954 4262
rect 2990 4258 2994 4262
rect 3006 4258 3010 4262
rect 3022 4258 3026 4262
rect 3030 4258 3034 4262
rect 3070 4259 3074 4263
rect 3166 4258 3170 4262
rect 3182 4258 3186 4262
rect 3222 4258 3226 4262
rect 3238 4258 3242 4262
rect 3270 4258 3274 4262
rect 3310 4258 3314 4262
rect 3438 4258 3442 4262
rect 3446 4258 3450 4262
rect 3462 4258 3466 4262
rect 3486 4258 3490 4262
rect 3494 4258 3498 4262
rect 3526 4258 3530 4262
rect 3550 4258 3554 4262
rect 3558 4258 3562 4262
rect 3598 4258 3602 4262
rect 3614 4258 3618 4262
rect 3630 4258 3634 4262
rect 3654 4258 3658 4262
rect 3686 4258 3690 4262
rect 3702 4258 3706 4262
rect 3718 4258 3722 4262
rect 3726 4258 3730 4262
rect 3766 4258 3770 4262
rect 3790 4258 3794 4262
rect 3830 4258 3834 4262
rect 3838 4258 3842 4262
rect 3878 4259 3882 4263
rect 3910 4258 3914 4262
rect 4030 4259 4034 4263
rect 4110 4258 4114 4262
rect 4118 4258 4122 4262
rect 4150 4258 4154 4262
rect 4166 4258 4170 4262
rect 4206 4258 4210 4262
rect 4230 4258 4234 4262
rect 4246 4258 4250 4262
rect 4262 4258 4266 4262
rect 4278 4258 4282 4262
rect 4294 4258 4298 4262
rect 4318 4258 4322 4262
rect 4350 4258 4354 4262
rect 4366 4258 4370 4262
rect 4398 4258 4402 4262
rect 4446 4258 4450 4262
rect 4454 4258 4458 4262
rect 4542 4258 4546 4262
rect 4550 4258 4554 4262
rect 4574 4258 4578 4262
rect 4590 4258 4594 4262
rect 4638 4258 4642 4262
rect 4686 4258 4690 4262
rect 4742 4258 4746 4262
rect 4750 4258 4754 4262
rect 4782 4258 4786 4262
rect 4822 4258 4826 4262
rect 4830 4258 4834 4262
rect 4854 4258 4858 4262
rect 4894 4258 4898 4262
rect 4926 4259 4930 4263
rect 4990 4258 4994 4262
rect 5006 4258 5010 4262
rect 5022 4258 5026 4262
rect 5046 4258 5050 4262
rect 5062 4258 5066 4262
rect 5102 4258 5106 4262
rect 5134 4258 5138 4262
rect 5150 4258 5154 4262
rect 5174 4258 5178 4262
rect 5246 4258 5250 4262
rect 5270 4259 5274 4263
rect 102 4248 106 4252
rect 246 4248 250 4252
rect 382 4248 386 4252
rect 478 4248 482 4252
rect 550 4248 554 4252
rect 718 4248 722 4252
rect 774 4248 778 4252
rect 782 4248 786 4252
rect 870 4248 874 4252
rect 958 4248 962 4252
rect 1126 4248 1130 4252
rect 1470 4248 1474 4252
rect 1638 4248 1642 4252
rect 1678 4248 1682 4252
rect 1758 4248 1762 4252
rect 1774 4248 1778 4252
rect 1790 4248 1794 4252
rect 1798 4248 1802 4252
rect 1974 4248 1978 4252
rect 2206 4248 2210 4252
rect 2350 4248 2354 4252
rect 2382 4248 2386 4252
rect 2486 4248 2490 4252
rect 2510 4248 2514 4252
rect 2814 4248 2818 4252
rect 2838 4248 2842 4252
rect 2926 4248 2930 4252
rect 2934 4248 2938 4252
rect 3006 4248 3010 4252
rect 3038 4248 3042 4252
rect 3182 4248 3186 4252
rect 3614 4248 3618 4252
rect 3670 4248 3674 4252
rect 3718 4248 3722 4252
rect 3750 4248 3754 4252
rect 3782 4248 3786 4252
rect 3814 4248 3818 4252
rect 3822 4248 3826 4252
rect 4182 4248 4186 4252
rect 4190 4248 4194 4252
rect 4222 4248 4226 4252
rect 4382 4248 4386 4252
rect 4422 4248 4426 4252
rect 4558 4248 4562 4252
rect 4806 4248 4810 4252
rect 5030 4248 5034 4252
rect 5166 4248 5170 4252
rect 630 4238 634 4242
rect 878 4238 882 4242
rect 942 4238 946 4242
rect 1086 4238 1090 4242
rect 1286 4238 1290 4242
rect 1694 4238 1698 4242
rect 1862 4238 1866 4242
rect 1950 4238 1954 4242
rect 2190 4238 2194 4242
rect 2750 4238 2754 4242
rect 3630 4238 3634 4242
rect 3798 4238 3802 4242
rect 4294 4238 4298 4242
rect 4662 4238 4666 4242
rect 398 4228 402 4232
rect 1966 4228 1970 4232
rect 214 4218 218 4222
rect 238 4218 242 4222
rect 1078 4218 1082 4222
rect 1382 4218 1386 4222
rect 1502 4218 1506 4222
rect 1622 4218 1626 4222
rect 1726 4218 1730 4222
rect 1814 4218 1818 4222
rect 1990 4218 1994 4222
rect 2198 4218 2202 4222
rect 2406 4218 2410 4222
rect 2470 4218 2474 4222
rect 2582 4218 2586 4222
rect 3382 4218 3386 4222
rect 3470 4218 3474 4222
rect 3510 4218 3514 4222
rect 3574 4218 3578 4222
rect 3734 4218 3738 4222
rect 3942 4218 3946 4222
rect 4166 4218 4170 4222
rect 4206 4218 4210 4222
rect 4262 4218 4266 4222
rect 4350 4218 4354 4222
rect 4798 4218 4802 4222
rect 5046 4218 5050 4222
rect 5070 4218 5074 4222
rect 5150 4218 5154 4222
rect 330 4203 334 4207
rect 337 4203 341 4207
rect 1354 4203 1358 4207
rect 1361 4203 1365 4207
rect 2386 4203 2390 4207
rect 2393 4203 2397 4207
rect 3402 4203 3406 4207
rect 3409 4203 3413 4207
rect 4426 4203 4430 4207
rect 4433 4203 4437 4207
rect 14 4188 18 4192
rect 102 4188 106 4192
rect 222 4188 226 4192
rect 358 4188 362 4192
rect 470 4188 474 4192
rect 494 4188 498 4192
rect 534 4188 538 4192
rect 550 4188 554 4192
rect 566 4188 570 4192
rect 750 4188 754 4192
rect 814 4188 818 4192
rect 854 4188 858 4192
rect 1246 4188 1250 4192
rect 1510 4188 1514 4192
rect 1686 4188 1690 4192
rect 1814 4188 1818 4192
rect 2638 4188 2642 4192
rect 2942 4188 2946 4192
rect 3054 4188 3058 4192
rect 3798 4188 3802 4192
rect 4358 4188 4362 4192
rect 4374 4188 4378 4192
rect 4646 4188 4650 4192
rect 5198 4188 5202 4192
rect 5270 4188 5274 4192
rect 662 4178 666 4182
rect 2302 4178 2306 4182
rect 3022 4178 3026 4182
rect 4734 4178 4738 4182
rect 158 4168 162 4172
rect 222 4168 226 4172
rect 230 4168 234 4172
rect 526 4168 530 4172
rect 574 4168 578 4172
rect 606 4168 610 4172
rect 614 4168 618 4172
rect 654 4168 658 4172
rect 1166 4168 1170 4172
rect 1206 4168 1210 4172
rect 1886 4168 1890 4172
rect 2030 4168 2034 4172
rect 2198 4168 2202 4172
rect 2662 4168 2666 4172
rect 2750 4168 2754 4172
rect 2822 4168 2826 4172
rect 3622 4168 3626 4172
rect 4070 4168 4074 4172
rect 4390 4168 4394 4172
rect 4574 4168 4578 4172
rect 4918 4168 4922 4172
rect 22 4158 26 4162
rect 86 4158 90 4162
rect 214 4158 218 4162
rect 246 4158 250 4162
rect 374 4158 378 4162
rect 478 4158 482 4162
rect 510 4158 514 4162
rect 590 4158 594 4162
rect 622 4158 626 4162
rect 678 4158 682 4162
rect 734 4158 738 4162
rect 758 4158 762 4162
rect 886 4158 890 4162
rect 1182 4158 1186 4162
rect 158 4148 162 4152
rect 174 4148 178 4152
rect 222 4148 226 4152
rect 286 4148 290 4152
rect 294 4148 298 4152
rect 342 4148 346 4152
rect 414 4148 418 4152
rect 494 4148 498 4152
rect 518 4148 522 4152
rect 542 4148 546 4152
rect 582 4148 586 4152
rect 614 4148 618 4152
rect 662 4148 666 4152
rect 694 4148 698 4152
rect 790 4148 794 4152
rect 846 4148 850 4152
rect 1046 4147 1050 4151
rect 1110 4148 1114 4152
rect 1126 4148 1130 4152
rect 1182 4148 1186 4152
rect 1222 4148 1226 4152
rect 1246 4148 1250 4152
rect 1270 4158 1274 4162
rect 1454 4158 1458 4162
rect 1486 4158 1490 4162
rect 1286 4148 1290 4152
rect 1326 4147 1330 4151
rect 1438 4148 1442 4152
rect 1462 4148 1466 4152
rect 1470 4148 1474 4152
rect 1670 4158 1674 4162
rect 1830 4158 1834 4162
rect 1510 4148 1514 4152
rect 1550 4148 1554 4152
rect 1630 4148 1634 4152
rect 1686 4148 1690 4152
rect 1934 4158 1938 4162
rect 2078 4158 2082 4162
rect 2110 4158 2114 4162
rect 2598 4158 2602 4162
rect 1734 4148 1738 4152
rect 1758 4148 1762 4152
rect 1798 4148 1802 4152
rect 1846 4148 1850 4152
rect 1878 4148 1882 4152
rect 1902 4148 1906 4152
rect 1918 4148 1922 4152
rect 1934 4148 1938 4152
rect 1966 4147 1970 4151
rect 2054 4148 2058 4152
rect 2070 4148 2074 4152
rect 2086 4148 2090 4152
rect 2142 4148 2146 4152
rect 2150 4148 2154 4152
rect 2182 4148 2186 4152
rect 2190 4148 2194 4152
rect 2254 4148 2258 4152
rect 2318 4148 2322 4152
rect 2326 4148 2330 4152
rect 2334 4148 2338 4152
rect 2430 4147 2434 4151
rect 2462 4148 2466 4152
rect 2510 4148 2514 4152
rect 2558 4148 2562 4152
rect 2590 4148 2594 4152
rect 2614 4148 2618 4152
rect 2638 4148 2642 4152
rect 2678 4148 2682 4152
rect 2694 4148 2698 4152
rect 2734 4148 2738 4152
rect 2742 4148 2746 4152
rect 2750 4148 2754 4152
rect 2790 4158 2794 4162
rect 2806 4158 2810 4162
rect 2774 4148 2778 4152
rect 2806 4148 2810 4152
rect 2854 4148 2858 4152
rect 2878 4148 2882 4152
rect 2934 4148 2938 4152
rect 2966 4158 2970 4162
rect 3038 4158 3042 4162
rect 3086 4158 3090 4162
rect 3302 4158 3306 4162
rect 4062 4158 4066 4162
rect 4126 4158 4130 4162
rect 4342 4158 4346 4162
rect 4654 4158 4658 4162
rect 4718 4158 4722 4162
rect 4838 4158 4842 4162
rect 4902 4158 4906 4162
rect 5110 4158 5114 4162
rect 5286 4158 5290 4162
rect 2982 4148 2986 4152
rect 3022 4148 3026 4152
rect 3086 4148 3090 4152
rect 3102 4148 3106 4152
rect 3118 4148 3122 4152
rect 3126 4148 3130 4152
rect 3150 4148 3154 4152
rect 3214 4148 3218 4152
rect 3238 4148 3242 4152
rect 3278 4148 3282 4152
rect 3334 4148 3338 4152
rect 3374 4148 3378 4152
rect 6 4138 10 4142
rect 78 4138 82 4142
rect 110 4138 114 4142
rect 118 4138 122 4142
rect 134 4138 138 4142
rect 166 4138 170 4142
rect 182 4138 186 4142
rect 254 4138 258 4142
rect 278 4138 282 4142
rect 286 4138 290 4142
rect 310 4138 314 4142
rect 350 4138 354 4142
rect 390 4138 394 4142
rect 502 4138 506 4142
rect 710 4138 714 4142
rect 758 4138 762 4142
rect 870 4138 874 4142
rect 902 4138 906 4142
rect 926 4138 930 4142
rect 974 4138 978 4142
rect 1030 4138 1034 4142
rect 1174 4138 1178 4142
rect 1230 4138 1234 4142
rect 1238 4138 1242 4142
rect 1294 4138 1298 4142
rect 1310 4138 1314 4142
rect 1462 4138 1466 4142
rect 1518 4138 1522 4142
rect 1566 4138 1570 4142
rect 1654 4138 1658 4142
rect 1694 4138 1698 4142
rect 1854 4138 1858 4142
rect 1878 4138 1882 4142
rect 1910 4138 1914 4142
rect 1950 4138 1954 4142
rect 2054 4138 2058 4142
rect 2086 4138 2090 4142
rect 2118 4138 2122 4142
rect 2134 4138 2138 4142
rect 2230 4138 2234 4142
rect 2262 4138 2266 4142
rect 2366 4138 2370 4142
rect 2550 4138 2554 4142
rect 2622 4138 2626 4142
rect 2630 4138 2634 4142
rect 2686 4138 2690 4142
rect 2710 4140 2714 4144
rect 2718 4138 2722 4142
rect 2726 4138 2730 4142
rect 2782 4138 2786 4142
rect 2814 4138 2818 4142
rect 2918 4138 2922 4142
rect 2990 4138 2994 4142
rect 3078 4138 3082 4142
rect 3406 4147 3410 4151
rect 3470 4148 3474 4152
rect 3502 4148 3506 4152
rect 3110 4138 3114 4142
rect 3158 4138 3162 4142
rect 3278 4138 3282 4142
rect 3310 4138 3314 4142
rect 3446 4138 3450 4142
rect 3478 4138 3482 4142
rect 3494 4138 3498 4142
rect 3502 4138 3506 4142
rect 3558 4147 3562 4151
rect 3662 4148 3666 4152
rect 3774 4148 3778 4152
rect 3782 4148 3786 4152
rect 3790 4148 3794 4152
rect 3846 4148 3850 4152
rect 3870 4148 3874 4152
rect 3950 4147 3954 4151
rect 4038 4148 4042 4152
rect 4046 4148 4050 4152
rect 4094 4148 4098 4152
rect 4102 4148 4106 4152
rect 4150 4148 4154 4152
rect 4158 4148 4162 4152
rect 4182 4148 4186 4152
rect 4222 4148 4226 4152
rect 4302 4148 4306 4152
rect 4366 4148 4370 4152
rect 4430 4148 4434 4152
rect 4518 4148 4522 4152
rect 4598 4148 4602 4152
rect 4630 4148 4634 4152
rect 4678 4148 4682 4152
rect 4710 4148 4714 4152
rect 4734 4148 4738 4152
rect 4750 4148 4754 4152
rect 4766 4148 4770 4152
rect 4774 4148 4778 4152
rect 4798 4148 4802 4152
rect 4822 4148 4826 4152
rect 4846 4148 4850 4152
rect 4878 4148 4882 4152
rect 4974 4148 4978 4152
rect 4998 4148 5002 4152
rect 5070 4148 5074 4152
rect 5150 4148 5154 4152
rect 5182 4148 5186 4152
rect 5198 4148 5202 4152
rect 5214 4148 5218 4152
rect 5230 4148 5234 4152
rect 5270 4148 5274 4152
rect 3542 4138 3546 4142
rect 3638 4138 3642 4142
rect 3726 4138 3730 4142
rect 3742 4138 3746 4142
rect 4038 4138 4042 4142
rect 4086 4138 4090 4142
rect 4102 4138 4106 4142
rect 4182 4138 4186 4142
rect 4214 4138 4218 4142
rect 4326 4138 4330 4142
rect 4366 4138 4370 4142
rect 4454 4138 4458 4142
rect 4606 4138 4610 4142
rect 4622 4138 4626 4142
rect 4638 4138 4642 4142
rect 4654 4138 4658 4142
rect 4702 4138 4706 4142
rect 4742 4138 4746 4142
rect 4806 4138 4810 4142
rect 4830 4138 4834 4142
rect 4854 4138 4858 4142
rect 4870 4138 4874 4142
rect 4902 4138 4906 4142
rect 4918 4138 4922 4142
rect 5158 4138 5162 4142
rect 5174 4138 5178 4142
rect 5190 4138 5194 4142
rect 5222 4138 5226 4142
rect 5262 4138 5266 4142
rect 142 4128 146 4132
rect 198 4128 202 4132
rect 262 4128 266 4132
rect 326 4128 330 4132
rect 438 4128 442 4132
rect 558 4128 562 4132
rect 638 4128 642 4132
rect 814 4128 818 4132
rect 894 4128 898 4132
rect 1414 4128 1418 4132
rect 1526 4128 1530 4132
rect 2046 4128 2050 4132
rect 2118 4128 2122 4132
rect 2398 4128 2402 4132
rect 2534 4128 2538 4132
rect 2998 4128 3002 4132
rect 3358 4128 3362 4132
rect 3454 4128 3458 4132
rect 3526 4128 3530 4132
rect 3806 4128 3810 4132
rect 4134 4128 4138 4132
rect 4198 4128 4202 4132
rect 4750 4128 4754 4132
rect 4894 4128 4898 4132
rect 5006 4128 5010 4132
rect 5246 4128 5250 4132
rect 62 4118 66 4122
rect 134 4118 138 4122
rect 598 4118 602 4122
rect 678 4118 682 4122
rect 918 4118 922 4122
rect 942 4118 946 4122
rect 982 4118 986 4122
rect 1390 4118 1394 4122
rect 1534 4118 1538 4122
rect 1574 4118 1578 4122
rect 1830 4118 1834 4122
rect 2038 4118 2042 4122
rect 2126 4118 2130 4122
rect 2174 4118 2178 4122
rect 2494 4118 2498 4122
rect 2526 4118 2530 4122
rect 2574 4118 2578 4122
rect 2598 4118 2602 4122
rect 2758 4118 2762 4122
rect 3518 4118 3522 4122
rect 3814 4118 3818 4122
rect 4126 4118 4130 4122
rect 4142 4118 4146 4122
rect 4206 4118 4210 4122
rect 4374 4118 4378 4122
rect 4694 4118 4698 4122
rect 4782 4118 4786 4122
rect 850 4103 854 4107
rect 857 4103 861 4107
rect 1874 4103 1878 4107
rect 1881 4103 1885 4107
rect 2890 4103 2894 4107
rect 2897 4103 2901 4107
rect 3922 4103 3926 4107
rect 3929 4103 3933 4107
rect 4938 4103 4942 4107
rect 4945 4103 4949 4107
rect 6 4088 10 4092
rect 134 4088 138 4092
rect 166 4088 170 4092
rect 198 4088 202 4092
rect 270 4088 274 4092
rect 342 4088 346 4092
rect 382 4088 386 4092
rect 502 4088 506 4092
rect 518 4088 522 4092
rect 542 4088 546 4092
rect 590 4088 594 4092
rect 622 4088 626 4092
rect 686 4088 690 4092
rect 702 4088 706 4092
rect 718 4088 722 4092
rect 1046 4088 1050 4092
rect 1286 4088 1290 4092
rect 1310 4088 1314 4092
rect 1446 4088 1450 4092
rect 1534 4088 1538 4092
rect 1606 4088 1610 4092
rect 1710 4088 1714 4092
rect 1742 4088 1746 4092
rect 1902 4088 1906 4092
rect 2558 4088 2562 4092
rect 2638 4088 2642 4092
rect 2926 4088 2930 4092
rect 3326 4088 3330 4092
rect 3510 4088 3514 4092
rect 3886 4088 3890 4092
rect 3982 4088 3986 4092
rect 4070 4088 4074 4092
rect 4310 4088 4314 4092
rect 4390 4088 4394 4092
rect 4518 4088 4522 4092
rect 4534 4088 4538 4092
rect 4630 4088 4634 4092
rect 4726 4088 4730 4092
rect 198 4078 202 4082
rect 390 4078 394 4082
rect 398 4078 402 4082
rect 462 4078 466 4082
rect 510 4078 514 4082
rect 550 4078 554 4082
rect 558 4078 562 4082
rect 766 4078 770 4082
rect 878 4078 882 4082
rect 1190 4078 1194 4082
rect 1358 4078 1362 4082
rect 1566 4078 1570 4082
rect 1718 4078 1722 4082
rect 1750 4078 1754 4082
rect 1758 4078 1762 4082
rect 1886 4078 1890 4082
rect 2326 4078 2330 4082
rect 3270 4078 3274 4082
rect 3278 4078 3282 4082
rect 3518 4078 3522 4082
rect 4198 4078 4202 4082
rect 4326 4078 4330 4082
rect 4342 4078 4346 4082
rect 4382 4078 4386 4082
rect 5182 4078 5186 4082
rect 5254 4078 5258 4082
rect 86 4068 90 4072
rect 102 4068 106 4072
rect 150 4068 154 4072
rect 182 4068 186 4072
rect 198 4068 202 4072
rect 230 4068 234 4072
rect 286 4068 290 4072
rect 366 4068 370 4072
rect 414 4068 418 4072
rect 438 4068 442 4072
rect 478 4068 482 4072
rect 534 4068 538 4072
rect 550 4068 554 4072
rect 574 4068 578 4072
rect 606 4068 610 4072
rect 614 4068 618 4072
rect 670 4068 674 4072
rect 710 4068 714 4072
rect 726 4068 730 4072
rect 782 4068 786 4072
rect 910 4068 914 4072
rect 918 4068 922 4072
rect 62 4058 66 4062
rect 206 4058 210 4062
rect 310 4058 314 4062
rect 358 4058 362 4062
rect 374 4058 378 4062
rect 462 4058 466 4062
rect 486 4058 490 4062
rect 526 4058 530 4062
rect 646 4058 650 4062
rect 798 4059 802 4063
rect 1030 4068 1034 4072
rect 1126 4068 1130 4072
rect 1150 4068 1154 4072
rect 1230 4068 1234 4072
rect 1302 4068 1306 4072
rect 1366 4068 1370 4072
rect 1398 4068 1402 4072
rect 1430 4068 1434 4072
rect 1454 4068 1458 4072
rect 1510 4068 1514 4072
rect 1526 4068 1530 4072
rect 1582 4068 1586 4072
rect 1598 4068 1602 4072
rect 1654 4068 1658 4072
rect 1734 4068 1738 4072
rect 1782 4068 1786 4072
rect 1814 4068 1818 4072
rect 1854 4068 1858 4072
rect 1934 4068 1938 4072
rect 1950 4068 1954 4072
rect 2102 4068 2106 4072
rect 2118 4068 2122 4072
rect 2230 4068 2234 4072
rect 2350 4068 2354 4072
rect 2406 4068 2410 4072
rect 2462 4068 2466 4072
rect 2478 4068 2482 4072
rect 2566 4068 2570 4072
rect 2622 4068 2626 4072
rect 2686 4068 2690 4072
rect 2750 4068 2754 4072
rect 2766 4068 2770 4072
rect 2774 4068 2778 4072
rect 2830 4068 2834 4072
rect 2846 4068 2850 4072
rect 3014 4068 3018 4072
rect 3054 4068 3058 4072
rect 3102 4068 3106 4072
rect 3118 4068 3122 4072
rect 3222 4068 3226 4072
rect 3262 4068 3266 4072
rect 3286 4068 3290 4072
rect 3302 4068 3306 4072
rect 3350 4068 3354 4072
rect 3390 4068 3394 4072
rect 3502 4068 3506 4072
rect 3606 4068 3610 4072
rect 3622 4068 3626 4072
rect 3678 4068 3682 4072
rect 3710 4068 3714 4072
rect 3726 4068 3730 4072
rect 3774 4068 3778 4072
rect 3790 4068 3794 4072
rect 3894 4068 3898 4072
rect 3942 4068 3946 4072
rect 3958 4068 3962 4072
rect 3990 4068 3994 4072
rect 4046 4068 4050 4072
rect 4126 4068 4130 4072
rect 4142 4068 4146 4072
rect 4230 4068 4234 4072
rect 830 4058 834 4062
rect 902 4058 906 4062
rect 918 4058 922 4062
rect 942 4058 946 4062
rect 990 4058 994 4062
rect 998 4058 1002 4062
rect 1110 4059 1114 4063
rect 1142 4058 1146 4062
rect 1158 4058 1162 4062
rect 1174 4058 1178 4062
rect 1222 4059 1226 4063
rect 1254 4058 1258 4062
rect 1294 4058 1298 4062
rect 1326 4058 1330 4062
rect 1342 4058 1346 4062
rect 1382 4058 1386 4062
rect 1390 4058 1394 4062
rect 1462 4058 1466 4062
rect 1502 4058 1506 4062
rect 1550 4058 1554 4062
rect 1590 4058 1594 4062
rect 1662 4058 1666 4062
rect 1702 4058 1706 4062
rect 1726 4058 1730 4062
rect 1774 4058 1778 4062
rect 1790 4058 1794 4062
rect 1806 4058 1810 4062
rect 1822 4058 1826 4062
rect 1846 4058 1850 4062
rect 1854 4058 1858 4062
rect 1918 4058 1922 4062
rect 1942 4058 1946 4062
rect 1966 4058 1970 4062
rect 1990 4058 1994 4062
rect 1998 4058 2002 4062
rect 2086 4059 2090 4063
rect 2126 4058 2130 4062
rect 2134 4058 2138 4062
rect 2158 4058 2162 4062
rect 2182 4058 2186 4062
rect 2190 4058 2194 4062
rect 2238 4058 2242 4062
rect 2310 4058 2314 4062
rect 2318 4058 2322 4062
rect 2342 4058 2346 4062
rect 2366 4058 2370 4062
rect 2414 4058 2418 4062
rect 2438 4058 2442 4062
rect 2454 4058 2458 4062
rect 2502 4058 2506 4062
rect 2574 4058 2578 4062
rect 2582 4058 2586 4062
rect 2662 4058 2666 4062
rect 2694 4058 2698 4062
rect 2726 4058 2730 4062
rect 2734 4058 2738 4062
rect 2766 4058 2770 4062
rect 2782 4058 2786 4062
rect 2830 4058 2834 4062
rect 2862 4059 2866 4063
rect 2894 4058 2898 4062
rect 2942 4058 2946 4062
rect 3022 4058 3026 4062
rect 3094 4058 3098 4062
rect 3134 4059 3138 4063
rect 3222 4058 3226 4062
rect 3230 4058 3234 4062
rect 3238 4058 3242 4062
rect 3254 4058 3258 4062
rect 3294 4058 3298 4062
rect 3350 4058 3354 4062
rect 3358 4058 3362 4062
rect 3422 4059 3426 4063
rect 3454 4058 3458 4062
rect 3494 4058 3498 4062
rect 3590 4059 3594 4063
rect 4286 4068 4290 4072
rect 4350 4068 4354 4072
rect 4382 4068 4386 4072
rect 4398 4068 4402 4072
rect 4462 4068 4466 4072
rect 4622 4068 4626 4072
rect 4710 4068 4714 4072
rect 4734 4068 4738 4072
rect 4806 4068 4810 4072
rect 4918 4068 4922 4072
rect 5006 4068 5010 4072
rect 5046 4068 5050 4072
rect 5110 4068 5114 4072
rect 5166 4068 5170 4072
rect 3630 4058 3634 4062
rect 3670 4058 3674 4062
rect 3678 4058 3682 4062
rect 3702 4058 3706 4062
rect 3718 4058 3722 4062
rect 3734 4058 3738 4062
rect 3766 4058 3770 4062
rect 3814 4058 3818 4062
rect 3950 4058 3954 4062
rect 3966 4058 3970 4062
rect 4006 4058 4010 4062
rect 4030 4058 4034 4062
rect 4046 4058 4050 4062
rect 4054 4058 4058 4062
rect 4086 4058 4090 4062
rect 4110 4058 4114 4062
rect 4118 4058 4122 4062
rect 4158 4058 4162 4062
rect 4174 4058 4178 4062
rect 4182 4058 4186 4062
rect 4190 4058 4194 4062
rect 4214 4058 4218 4062
rect 4222 4058 4226 4062
rect 4262 4058 4266 4062
rect 4278 4058 4282 4062
rect 4294 4058 4298 4062
rect 4326 4058 4330 4062
rect 4358 4058 4362 4062
rect 4406 4058 4410 4062
rect 4454 4059 4458 4063
rect 4486 4058 4490 4062
rect 4550 4058 4554 4062
rect 4558 4058 4562 4062
rect 4694 4059 4698 4063
rect 4782 4058 4786 4062
rect 4894 4058 4898 4062
rect 5014 4059 5018 4063
rect 5054 4058 5058 4062
rect 5094 4058 5098 4062
rect 5150 4058 5154 4062
rect 5158 4058 5162 4062
rect 5230 4058 5234 4062
rect 158 4048 162 4052
rect 270 4048 274 4052
rect 318 4048 322 4052
rect 342 4048 346 4052
rect 422 4048 426 4052
rect 470 4048 474 4052
rect 590 4048 594 4052
rect 630 4048 634 4052
rect 638 4048 642 4052
rect 686 4048 690 4052
rect 838 4048 842 4052
rect 886 4048 890 4052
rect 902 4048 906 4052
rect 942 4048 946 4052
rect 1390 4048 1394 4052
rect 1422 4048 1426 4052
rect 1446 4048 1450 4052
rect 1478 4048 1482 4052
rect 1502 4048 1506 4052
rect 1574 4048 1578 4052
rect 1822 4048 1826 4052
rect 1926 4048 1930 4052
rect 2142 4048 2146 4052
rect 2294 4048 2298 4052
rect 2382 4048 2386 4052
rect 2430 4048 2434 4052
rect 2438 4048 2442 4052
rect 2598 4048 2602 4052
rect 2742 4048 2746 4052
rect 2798 4048 2802 4052
rect 2822 4048 2826 4052
rect 3070 4048 3074 4052
rect 3246 4048 3250 4052
rect 3310 4048 3314 4052
rect 3390 4048 3394 4052
rect 3542 4048 3546 4052
rect 3630 4048 3634 4052
rect 3654 4048 3658 4052
rect 3686 4048 3690 4052
rect 3750 4048 3754 4052
rect 3910 4048 3914 4052
rect 4070 4048 4074 4052
rect 4142 4048 4146 4052
rect 4174 4048 4178 4052
rect 4254 4048 4258 4052
rect 4262 4048 4266 4052
rect 4374 4048 4378 4052
rect 5054 4048 5058 4052
rect 5134 4048 5138 4052
rect 254 4038 258 4042
rect 302 4038 306 4042
rect 414 4038 418 4042
rect 454 4038 458 4042
rect 654 4038 658 4042
rect 950 4038 954 4042
rect 1622 4038 1626 4042
rect 1862 4038 1866 4042
rect 1982 4038 1986 4042
rect 3094 4038 3098 4042
rect 5078 4038 5082 4042
rect 310 4028 314 4032
rect 662 4028 666 4032
rect 4950 4028 4954 4032
rect 5190 4028 5194 4032
rect 702 4018 706 4022
rect 734 4018 738 4022
rect 854 4018 858 4022
rect 1286 4018 1290 4022
rect 1406 4018 1410 4022
rect 1774 4018 1778 4022
rect 1806 4018 1810 4022
rect 2006 4018 2010 4022
rect 2174 4018 2178 4022
rect 2366 4018 2370 4022
rect 2414 4018 2418 4022
rect 2638 4018 2642 4022
rect 2710 4018 2714 4022
rect 3038 4018 3042 4022
rect 3486 4018 3490 4022
rect 3526 4018 3530 4022
rect 4094 4018 4098 4022
rect 4134 4018 4138 4022
rect 4238 4018 4242 4022
rect 4518 4018 4522 4022
rect 4566 4018 4570 4022
rect 4822 4018 4826 4022
rect 5174 4018 5178 4022
rect 330 4003 334 4007
rect 337 4003 341 4007
rect 1354 4003 1358 4007
rect 1361 4003 1365 4007
rect 2386 4003 2390 4007
rect 2393 4003 2397 4007
rect 3402 4003 3406 4007
rect 3409 4003 3413 4007
rect 4426 4003 4430 4007
rect 4433 4003 4437 4007
rect 62 3988 66 3992
rect 102 3988 106 3992
rect 230 3988 234 3992
rect 270 3988 274 3992
rect 278 3988 282 3992
rect 294 3988 298 3992
rect 318 3988 322 3992
rect 430 3988 434 3992
rect 510 3988 514 3992
rect 542 3988 546 3992
rect 574 3988 578 3992
rect 606 3988 610 3992
rect 694 3988 698 3992
rect 1030 3988 1034 3992
rect 1270 3988 1274 3992
rect 1454 3988 1458 3992
rect 1518 3988 1522 3992
rect 1950 3988 1954 3992
rect 2102 3988 2106 3992
rect 2694 3988 2698 3992
rect 2894 3988 2898 3992
rect 3118 3988 3122 3992
rect 3206 3988 3210 3992
rect 3390 3988 3394 3992
rect 3470 3988 3474 3992
rect 3566 3988 3570 3992
rect 3646 3988 3650 3992
rect 4006 3988 4010 3992
rect 4038 3988 4042 3992
rect 4062 3988 4066 3992
rect 4358 3988 4362 3992
rect 4670 3988 4674 3992
rect 5190 3988 5194 3992
rect 5222 3988 5226 3992
rect 206 3978 210 3982
rect 366 3978 370 3982
rect 1350 3978 1354 3982
rect 3094 3978 3098 3982
rect 3222 3978 3226 3982
rect 3438 3978 3442 3982
rect 198 3968 202 3972
rect 222 3968 226 3972
rect 286 3968 290 3972
rect 358 3968 362 3972
rect 422 3968 426 3972
rect 454 3968 458 3972
rect 566 3968 570 3972
rect 598 3968 602 3972
rect 934 3968 938 3972
rect 1062 3968 1066 3972
rect 1286 3968 1290 3972
rect 1654 3968 1658 3972
rect 2230 3968 2234 3972
rect 2334 3968 2338 3972
rect 2942 3968 2946 3972
rect 3046 3968 3050 3972
rect 3326 3968 3330 3972
rect 3918 3968 3922 3972
rect 4374 3968 4378 3972
rect 4766 3968 4770 3972
rect 4782 3968 4786 3972
rect 4822 3968 4826 3972
rect 5014 3968 5018 3972
rect 5110 3968 5114 3972
rect 6 3958 10 3962
rect 142 3958 146 3962
rect 22 3948 26 3952
rect 38 3948 42 3952
rect 86 3948 90 3952
rect 62 3938 66 3942
rect 78 3938 82 3942
rect 86 3938 90 3942
rect 126 3948 130 3952
rect 238 3958 242 3962
rect 302 3958 306 3962
rect 310 3958 314 3962
rect 374 3958 378 3962
rect 406 3958 410 3962
rect 438 3958 442 3962
rect 470 3958 474 3962
rect 502 3958 506 3962
rect 582 3958 586 3962
rect 622 3958 626 3962
rect 678 3958 682 3962
rect 158 3948 162 3952
rect 166 3948 170 3952
rect 230 3948 234 3952
rect 254 3948 258 3952
rect 294 3948 298 3952
rect 366 3948 370 3952
rect 390 3948 394 3952
rect 406 3948 410 3952
rect 430 3948 434 3952
rect 454 3948 458 3952
rect 486 3948 490 3952
rect 510 3948 514 3952
rect 526 3948 530 3952
rect 574 3948 578 3952
rect 606 3948 610 3952
rect 630 3948 634 3952
rect 638 3948 642 3952
rect 686 3948 690 3952
rect 702 3948 706 3952
rect 734 3948 738 3952
rect 758 3948 762 3952
rect 174 3938 178 3942
rect 326 3938 330 3942
rect 382 3938 386 3942
rect 446 3938 450 3942
rect 478 3938 482 3942
rect 646 3938 650 3942
rect 702 3938 706 3942
rect 742 3938 746 3942
rect 790 3948 794 3952
rect 838 3948 842 3952
rect 894 3948 898 3952
rect 966 3948 970 3952
rect 974 3948 978 3952
rect 990 3958 994 3962
rect 1046 3958 1050 3962
rect 1078 3958 1082 3962
rect 1006 3948 1010 3952
rect 1030 3948 1034 3952
rect 1062 3948 1066 3952
rect 1118 3948 1122 3952
rect 1134 3948 1138 3952
rect 1222 3948 1226 3952
rect 1230 3948 1234 3952
rect 1286 3948 1290 3952
rect 1310 3958 1314 3962
rect 1414 3958 1418 3962
rect 1326 3948 1330 3952
rect 1374 3948 1378 3952
rect 1382 3948 1386 3952
rect 1534 3958 1538 3962
rect 1470 3948 1474 3952
rect 1502 3948 1506 3952
rect 1518 3948 1522 3952
rect 1542 3948 1546 3952
rect 1558 3948 1562 3952
rect 1598 3948 1602 3952
rect 1622 3948 1626 3952
rect 1670 3948 1674 3952
rect 1694 3958 1698 3962
rect 1750 3948 1754 3952
rect 1766 3948 1770 3952
rect 1790 3958 1794 3962
rect 2006 3958 2010 3962
rect 2022 3958 2026 3962
rect 2038 3958 2042 3962
rect 2166 3958 2170 3962
rect 2222 3958 2226 3962
rect 1806 3948 1810 3952
rect 1878 3948 1882 3952
rect 1950 3948 1954 3952
rect 1958 3948 1962 3952
rect 2006 3948 2010 3952
rect 2038 3948 2042 3952
rect 2054 3948 2058 3952
rect 2086 3948 2090 3952
rect 2094 3948 2098 3952
rect 2118 3948 2122 3952
rect 2126 3948 2130 3952
rect 2190 3948 2194 3952
rect 2198 3948 2202 3952
rect 2262 3948 2266 3952
rect 798 3938 802 3942
rect 958 3938 962 3942
rect 1014 3938 1018 3942
rect 1022 3938 1026 3942
rect 1054 3938 1058 3942
rect 1278 3938 1282 3942
rect 1334 3938 1338 3942
rect 1390 3938 1394 3942
rect 1446 3938 1450 3942
rect 1486 3938 1490 3942
rect 1510 3938 1514 3942
rect 1558 3938 1562 3942
rect 1662 3938 1666 3942
rect 1678 3938 1682 3942
rect 1718 3938 1722 3942
rect 2294 3947 2298 3951
rect 2334 3948 2338 3952
rect 2358 3958 2362 3962
rect 2534 3958 2538 3962
rect 2822 3958 2826 3962
rect 2854 3958 2858 3962
rect 3070 3958 3074 3962
rect 2374 3948 2378 3952
rect 2430 3948 2434 3952
rect 2502 3947 2506 3951
rect 2534 3948 2538 3952
rect 2550 3948 2554 3952
rect 2566 3948 2570 3952
rect 2622 3948 2626 3952
rect 2646 3948 2650 3952
rect 1758 3938 1762 3942
rect 1782 3938 1786 3942
rect 1814 3938 1818 3942
rect 1854 3938 1858 3942
rect 1902 3938 1906 3942
rect 1966 3938 1970 3942
rect 2014 3938 2018 3942
rect 2046 3938 2050 3942
rect 2062 3938 2066 3942
rect 2158 3938 2162 3942
rect 2190 3938 2194 3942
rect 2206 3938 2210 3942
rect 2310 3938 2314 3942
rect 2326 3938 2330 3942
rect 2382 3938 2386 3942
rect 2422 3938 2426 3942
rect 2766 3947 2770 3951
rect 2814 3948 2818 3952
rect 2846 3948 2850 3952
rect 2878 3948 2882 3952
rect 2926 3948 2930 3952
rect 3006 3948 3010 3952
rect 3094 3948 3098 3952
rect 3134 3948 3138 3952
rect 3150 3948 3154 3952
rect 3166 3948 3170 3952
rect 3182 3948 3186 3952
rect 3198 3948 3202 3952
rect 3286 3947 3290 3951
rect 3326 3948 3330 3952
rect 3350 3958 3354 3962
rect 3422 3958 3426 3962
rect 3510 3958 3514 3962
rect 3622 3958 3626 3962
rect 3638 3958 3642 3962
rect 3694 3958 3698 3962
rect 3366 3948 3370 3952
rect 3430 3948 3434 3952
rect 3470 3948 3474 3952
rect 3478 3948 3482 3952
rect 3510 3948 3514 3952
rect 3526 3948 3530 3952
rect 3606 3948 3610 3952
rect 3622 3948 3626 3952
rect 3646 3948 3650 3952
rect 3670 3948 3674 3952
rect 3718 3958 3722 3962
rect 4014 3958 4018 3962
rect 4222 3958 4226 3962
rect 4262 3958 4266 3962
rect 4494 3958 4498 3962
rect 4798 3958 4802 3962
rect 3718 3948 3722 3952
rect 3782 3948 3786 3952
rect 3862 3948 3866 3952
rect 3942 3948 3946 3952
rect 3974 3948 3978 3952
rect 4022 3948 4026 3952
rect 4054 3948 4058 3952
rect 4078 3948 4082 3952
rect 4086 3948 4090 3952
rect 4110 3948 4114 3952
rect 4118 3948 4122 3952
rect 2558 3938 2562 3942
rect 2598 3938 2602 3942
rect 2750 3938 2754 3942
rect 2838 3938 2842 3942
rect 2870 3938 2874 3942
rect 2918 3938 2922 3942
rect 2966 3938 2970 3942
rect 3054 3938 3058 3942
rect 3142 3938 3146 3942
rect 3158 3938 3162 3942
rect 3190 3938 3194 3942
rect 3262 3938 3266 3942
rect 3302 3938 3306 3942
rect 3318 3938 3322 3942
rect 3374 3938 3378 3942
rect 3382 3938 3386 3942
rect 3470 3938 3474 3942
rect 3486 3938 3490 3942
rect 3534 3938 3538 3942
rect 3542 3938 3546 3942
rect 3598 3938 3602 3942
rect 3614 3938 3618 3942
rect 3670 3938 3674 3942
rect 3726 3938 3730 3942
rect 3790 3938 3794 3942
rect 3950 3938 3954 3942
rect 3998 3938 4002 3942
rect 4150 3947 4154 3951
rect 4246 3948 4250 3952
rect 4270 3948 4274 3952
rect 4294 3948 4298 3952
rect 4302 3948 4306 3952
rect 4310 3948 4314 3952
rect 4334 3948 4338 3952
rect 4358 3948 4362 3952
rect 4166 3938 4170 3942
rect 4446 3947 4450 3951
rect 4510 3948 4514 3952
rect 4558 3948 4562 3952
rect 4622 3948 4626 3952
rect 4646 3948 4650 3952
rect 4654 3948 4658 3952
rect 4678 3948 4682 3952
rect 4726 3948 4730 3952
rect 4750 3948 4754 3952
rect 4798 3948 4802 3952
rect 4902 3958 4906 3962
rect 4982 3958 4986 3962
rect 4998 3958 5002 3962
rect 5118 3958 5122 3962
rect 5150 3958 5154 3962
rect 5206 3958 5210 3962
rect 4838 3948 4842 3952
rect 4870 3948 4874 3952
rect 4886 3948 4890 3952
rect 4966 3948 4970 3952
rect 4982 3948 4986 3952
rect 4998 3948 5002 3952
rect 5046 3947 5050 3951
rect 5070 3948 5074 3952
rect 5134 3948 5138 3952
rect 5166 3948 5170 3952
rect 5190 3948 5194 3952
rect 4350 3938 4354 3942
rect 4462 3938 4466 3942
rect 4518 3938 4522 3942
rect 4566 3938 4570 3942
rect 4686 3938 4690 3942
rect 4790 3938 4794 3942
rect 4846 3938 4850 3942
rect 4894 3938 4898 3942
rect 4910 3938 4914 3942
rect 4918 3940 4922 3944
rect 4958 3938 4962 3942
rect 4990 3938 4994 3942
rect 5142 3938 5146 3942
rect 5174 3938 5178 3942
rect 5182 3938 5186 3942
rect 5278 3938 5282 3942
rect 54 3928 58 3932
rect 62 3928 66 3932
rect 110 3928 114 3932
rect 182 3928 186 3932
rect 198 3928 202 3932
rect 526 3928 530 3932
rect 550 3928 554 3932
rect 686 3928 690 3932
rect 726 3928 730 3932
rect 766 3928 770 3932
rect 806 3928 810 3932
rect 822 3928 826 3932
rect 886 3928 890 3932
rect 1542 3928 1546 3932
rect 1934 3928 1938 3932
rect 1982 3928 1986 3932
rect 2078 3928 2082 3932
rect 2222 3928 2226 3932
rect 2246 3928 2250 3932
rect 2398 3928 2402 3932
rect 2502 3928 2506 3932
rect 2582 3928 2586 3932
rect 2798 3928 2802 3932
rect 2982 3928 2986 3932
rect 3110 3928 3114 3932
rect 3126 3928 3130 3932
rect 3214 3928 3218 3932
rect 3446 3928 3450 3932
rect 3582 3928 3586 3932
rect 3662 3928 3666 3932
rect 3958 3928 3962 3932
rect 3990 3928 3994 3932
rect 4070 3928 4074 3932
rect 4446 3928 4450 3932
rect 4598 3928 4602 3932
rect 4638 3928 4642 3932
rect 4854 3928 4858 3932
rect 5150 3928 5154 3932
rect 6 3918 10 3922
rect 502 3918 506 3922
rect 718 3918 722 3922
rect 950 3918 954 3922
rect 1174 3918 1178 3922
rect 1430 3918 1434 3922
rect 1454 3918 1458 3922
rect 1734 3918 1738 3922
rect 1822 3918 1826 3922
rect 2070 3918 2074 3922
rect 2150 3918 2154 3922
rect 2414 3918 2418 3922
rect 2438 3918 2442 3922
rect 2574 3918 2578 3922
rect 2702 3918 2706 3922
rect 2854 3918 2858 3922
rect 3182 3918 3186 3922
rect 3438 3918 3442 3922
rect 3590 3918 3594 3922
rect 3734 3918 3738 3922
rect 4278 3918 4282 3922
rect 4318 3918 4322 3922
rect 4382 3918 4386 3922
rect 4494 3918 4498 3922
rect 4630 3918 4634 3922
rect 4934 3918 4938 3922
rect 5110 3918 5114 3922
rect 5118 3918 5122 3922
rect 850 3903 854 3907
rect 857 3903 861 3907
rect 1874 3903 1878 3907
rect 1881 3903 1885 3907
rect 2890 3903 2894 3907
rect 2897 3903 2901 3907
rect 3922 3903 3926 3907
rect 3929 3903 3933 3907
rect 4938 3903 4942 3907
rect 4945 3903 4949 3907
rect 46 3888 50 3892
rect 94 3888 98 3892
rect 182 3888 186 3892
rect 222 3888 226 3892
rect 254 3888 258 3892
rect 278 3888 282 3892
rect 430 3888 434 3892
rect 470 3888 474 3892
rect 510 3888 514 3892
rect 526 3888 530 3892
rect 582 3888 586 3892
rect 822 3888 826 3892
rect 926 3888 930 3892
rect 1118 3888 1122 3892
rect 1486 3888 1490 3892
rect 1598 3888 1602 3892
rect 1670 3888 1674 3892
rect 1702 3888 1706 3892
rect 1790 3888 1794 3892
rect 1838 3888 1842 3892
rect 2158 3888 2162 3892
rect 2326 3888 2330 3892
rect 2486 3888 2490 3892
rect 2694 3888 2698 3892
rect 2726 3888 2730 3892
rect 2742 3888 2746 3892
rect 2926 3888 2930 3892
rect 3286 3888 3290 3892
rect 3318 3888 3322 3892
rect 3398 3888 3402 3892
rect 3590 3888 3594 3892
rect 3614 3888 3618 3892
rect 3638 3888 3642 3892
rect 3942 3888 3946 3892
rect 3974 3888 3978 3892
rect 4398 3888 4402 3892
rect 4478 3888 4482 3892
rect 4566 3888 4570 3892
rect 4894 3888 4898 3892
rect 54 3878 58 3882
rect 190 3878 194 3882
rect 358 3878 362 3882
rect 518 3878 522 3882
rect 590 3878 594 3882
rect 630 3878 634 3882
rect 950 3878 954 3882
rect 62 3868 66 3872
rect 70 3868 74 3872
rect 126 3868 130 3872
rect 158 3868 162 3872
rect 174 3868 178 3872
rect 198 3868 202 3872
rect 230 3868 234 3872
rect 262 3868 266 3872
rect 318 3868 322 3872
rect 382 3868 386 3872
rect 422 3868 426 3872
rect 438 3868 442 3872
rect 486 3868 490 3872
rect 566 3868 570 3872
rect 574 3868 578 3872
rect 694 3868 698 3872
rect 710 3868 714 3872
rect 758 3868 762 3872
rect 782 3868 786 3872
rect 846 3868 850 3872
rect 886 3868 890 3872
rect 942 3868 946 3872
rect 966 3878 970 3882
rect 1078 3878 1082 3882
rect 1150 3878 1154 3882
rect 1174 3878 1178 3882
rect 1206 3878 1210 3882
rect 1222 3878 1226 3882
rect 1462 3878 1466 3882
rect 1622 3878 1626 3882
rect 1006 3868 1010 3872
rect 1054 3868 1058 3872
rect 1078 3868 1082 3872
rect 1094 3868 1098 3872
rect 1110 3868 1114 3872
rect 1182 3868 1186 3872
rect 1214 3868 1218 3872
rect 1238 3868 1242 3872
rect 1334 3868 1338 3872
rect 1366 3868 1370 3872
rect 1382 3868 1386 3872
rect 1422 3868 1426 3872
rect 1454 3868 1458 3872
rect 1550 3868 1554 3872
rect 1774 3878 1778 3882
rect 2134 3878 2138 3882
rect 2270 3878 2274 3882
rect 1646 3868 1650 3872
rect 1662 3868 1666 3872
rect 1686 3868 1690 3872
rect 1814 3868 1818 3872
rect 1886 3868 1890 3872
rect 1902 3868 1906 3872
rect 1934 3868 1938 3872
rect 1966 3868 1970 3872
rect 1998 3868 2002 3872
rect 2030 3868 2034 3872
rect 2038 3868 2042 3872
rect 2086 3868 2090 3872
rect 2102 3868 2106 3872
rect 2254 3868 2258 3872
rect 2262 3868 2266 3872
rect 2286 3878 2290 3882
rect 2646 3878 2650 3882
rect 2734 3878 2738 3882
rect 3110 3878 3114 3882
rect 3494 3878 3498 3882
rect 3662 3878 3666 3882
rect 4230 3878 4234 3882
rect 4334 3878 4338 3882
rect 4430 3878 4434 3882
rect 4598 3878 4602 3882
rect 4606 3878 4610 3882
rect 4886 3878 4890 3882
rect 4934 3878 4938 3882
rect 5038 3878 5042 3882
rect 2342 3868 2346 3872
rect 2510 3868 2514 3872
rect 2638 3868 2642 3872
rect 2670 3868 2674 3872
rect 2702 3868 2706 3872
rect 2822 3868 2826 3872
rect 2838 3868 2842 3872
rect 2846 3868 2850 3872
rect 2878 3868 2882 3872
rect 2902 3868 2906 3872
rect 2974 3868 2978 3872
rect 3046 3868 3050 3872
rect 3150 3868 3154 3872
rect 3262 3868 3266 3872
rect 3278 3868 3282 3872
rect 3342 3868 3346 3872
rect 3574 3868 3578 3872
rect 3702 3868 3706 3872
rect 3742 3868 3746 3872
rect 3870 3868 3874 3872
rect 3910 3868 3914 3872
rect 3950 3868 3954 3872
rect 4062 3868 4066 3872
rect 4094 3868 4098 3872
rect 4118 3868 4122 3872
rect 4142 3868 4146 3872
rect 4318 3868 4322 3872
rect 4342 3868 4346 3872
rect 4390 3868 4394 3872
rect 4422 3868 4426 3872
rect 4486 3868 4490 3872
rect 4502 3868 4506 3872
rect 4534 3868 4538 3872
rect 4638 3868 4642 3872
rect 4686 3868 4690 3872
rect 4726 3868 4730 3872
rect 4750 3868 4754 3872
rect 4766 3868 4770 3872
rect 4854 3868 4858 3872
rect 4918 3868 4922 3872
rect 4958 3868 4962 3872
rect 4990 3868 4994 3872
rect 5134 3868 5138 3872
rect 5174 3868 5178 3872
rect 5254 3868 5258 3872
rect 46 3858 50 3862
rect 78 3858 82 3862
rect 118 3858 122 3862
rect 158 3858 162 3862
rect 166 3858 170 3862
rect 206 3858 210 3862
rect 238 3858 242 3862
rect 310 3858 314 3862
rect 318 3858 322 3862
rect 366 3858 370 3862
rect 374 3858 378 3862
rect 390 3858 394 3862
rect 462 3858 466 3862
rect 494 3858 498 3862
rect 534 3858 538 3862
rect 630 3858 634 3862
rect 654 3858 658 3862
rect 702 3858 706 3862
rect 750 3859 754 3863
rect 870 3858 874 3862
rect 934 3858 938 3862
rect 982 3858 986 3862
rect 1038 3858 1042 3862
rect 1062 3858 1066 3862
rect 1086 3858 1090 3862
rect 1094 3858 1098 3862
rect 1102 3858 1106 3862
rect 1134 3858 1138 3862
rect 1150 3858 1154 3862
rect 1174 3858 1178 3862
rect 1190 3858 1194 3862
rect 1206 3858 1210 3862
rect 1246 3858 1250 3862
rect 1318 3859 1322 3863
rect 1374 3858 1378 3862
rect 1414 3858 1418 3862
rect 1446 3858 1450 3862
rect 1502 3858 1506 3862
rect 1542 3858 1546 3862
rect 1606 3858 1610 3862
rect 1622 3858 1626 3862
rect 1654 3858 1658 3862
rect 1678 3858 1682 3862
rect 1710 3858 1714 3862
rect 1718 3858 1722 3862
rect 1750 3858 1754 3862
rect 1758 3858 1762 3862
rect 1814 3858 1818 3862
rect 1822 3858 1826 3862
rect 1910 3858 1914 3862
rect 1942 3858 1946 3862
rect 1990 3858 1994 3862
rect 2006 3858 2010 3862
rect 2046 3858 2050 3862
rect 2078 3858 2082 3862
rect 2094 3858 2098 3862
rect 2110 3858 2114 3862
rect 2150 3858 2154 3862
rect 2190 3858 2194 3862
rect 2222 3859 2226 3863
rect 2254 3858 2258 3862
rect 2302 3858 2306 3862
rect 2310 3858 2314 3862
rect 2350 3858 2354 3862
rect 2374 3858 2378 3862
rect 2414 3859 2418 3863
rect 2446 3858 2450 3862
rect 2502 3858 2506 3862
rect 2550 3858 2554 3862
rect 2574 3858 2578 3862
rect 2638 3858 2642 3862
rect 2662 3858 2666 3862
rect 2678 3858 2682 3862
rect 2710 3858 2714 3862
rect 2806 3859 2810 3863
rect 2862 3858 2866 3862
rect 2870 3858 2874 3862
rect 2902 3858 2906 3862
rect 2910 3858 2914 3862
rect 2966 3858 2970 3862
rect 3078 3858 3082 3862
rect 3086 3858 3090 3862
rect 3094 3858 3098 3862
rect 3118 3858 3122 3862
rect 3126 3858 3130 3862
rect 3230 3858 3234 3862
rect 3302 3858 3306 3862
rect 3334 3858 3338 3862
rect 3382 3858 3386 3862
rect 3494 3859 3498 3863
rect 3526 3858 3530 3862
rect 3534 3858 3538 3862
rect 3558 3858 3562 3862
rect 3598 3858 3602 3862
rect 3654 3858 3658 3862
rect 3678 3858 3682 3862
rect 3710 3858 3714 3862
rect 3718 3858 3722 3862
rect 3782 3858 3786 3862
rect 3814 3859 3818 3863
rect 3862 3858 3866 3862
rect 3878 3858 3882 3862
rect 3902 3858 3906 3862
rect 3918 3858 3922 3862
rect 4054 3858 4058 3862
rect 4102 3858 4106 3862
rect 4222 3858 4226 3862
rect 4270 3858 4274 3862
rect 4294 3858 4298 3862
rect 4302 3858 4306 3862
rect 4310 3858 4314 3862
rect 4350 3858 4354 3862
rect 4414 3858 4418 3862
rect 4462 3858 4466 3862
rect 4494 3858 4498 3862
rect 4510 3858 4514 3862
rect 4526 3858 4530 3862
rect 4542 3858 4546 3862
rect 4550 3858 4554 3862
rect 4606 3858 4610 3862
rect 4622 3858 4626 3862
rect 4686 3858 4690 3862
rect 4734 3858 4738 3862
rect 4782 3859 4786 3863
rect 4862 3858 4866 3862
rect 4902 3858 4906 3862
rect 4910 3858 4914 3862
rect 4998 3858 5002 3862
rect 5022 3858 5026 3862
rect 5118 3859 5122 3863
rect 5158 3858 5162 3862
rect 5166 3858 5170 3862
rect 5182 3858 5186 3862
rect 5262 3858 5266 3862
rect 102 3848 106 3852
rect 134 3848 138 3852
rect 150 3848 154 3852
rect 262 3848 266 3852
rect 278 3848 282 3852
rect 286 3848 290 3852
rect 302 3848 306 3852
rect 406 3848 410 3852
rect 454 3848 458 3852
rect 718 3848 722 3852
rect 990 3848 994 3852
rect 1046 3848 1050 3852
rect 1398 3848 1402 3852
rect 1430 3848 1434 3852
rect 1702 3848 1706 3852
rect 1838 3848 1842 3852
rect 1926 3848 1930 3852
rect 1958 3848 1962 3852
rect 2062 3848 2066 3852
rect 2126 3848 2130 3852
rect 2366 3848 2370 3852
rect 2486 3848 2490 3852
rect 2630 3848 2634 3852
rect 2646 3848 2650 3852
rect 2854 3848 2858 3852
rect 2926 3848 2930 3852
rect 3294 3848 3298 3852
rect 3366 3848 3370 3852
rect 3590 3848 3594 3852
rect 3846 3848 3850 3852
rect 3862 3848 3866 3852
rect 3878 3848 3882 3852
rect 3974 3848 3978 3852
rect 4126 3848 4130 3852
rect 4374 3848 4378 3852
rect 4398 3848 4402 3852
rect 4750 3848 4754 3852
rect 4846 3848 4850 3852
rect 4878 3848 4882 3852
rect 4982 3848 4986 3852
rect 5014 3848 5018 3852
rect 5150 3848 5154 3852
rect 118 3838 122 3842
rect 470 3838 474 3842
rect 1006 3838 1010 3842
rect 1254 3838 1258 3842
rect 1870 3838 1874 3842
rect 2478 3838 2482 3842
rect 3542 3838 3546 3842
rect 5070 3838 5074 3842
rect 5222 3838 5226 3842
rect 3038 3828 3042 3832
rect 4150 3828 4154 3832
rect 4862 3828 4866 3832
rect 478 3818 482 3822
rect 598 3818 602 3822
rect 1022 3818 1026 3822
rect 1222 3818 1226 3822
rect 1446 3818 1450 3822
rect 1470 3818 1474 3822
rect 1726 3818 1730 3822
rect 1766 3818 1770 3822
rect 1790 3818 1794 3822
rect 1910 3818 1914 3822
rect 1990 3818 1994 3822
rect 2110 3818 2114 3822
rect 2142 3818 2146 3822
rect 2606 3818 2610 3822
rect 2694 3818 2698 3822
rect 3102 3818 3106 3822
rect 3166 3818 3170 3822
rect 3358 3818 3362 3822
rect 3686 3818 3690 3822
rect 3750 3818 3754 3822
rect 3982 3818 3986 3822
rect 4278 3818 4282 3822
rect 4334 3818 4338 3822
rect 4350 3818 4354 3822
rect 4510 3818 4514 3822
rect 4614 3818 4618 3822
rect 4966 3818 4970 3822
rect 4998 3818 5002 3822
rect 5054 3818 5058 3822
rect 5190 3818 5194 3822
rect 5206 3818 5210 3822
rect 330 3803 334 3807
rect 337 3803 341 3807
rect 1354 3803 1358 3807
rect 1361 3803 1365 3807
rect 2386 3803 2390 3807
rect 2393 3803 2397 3807
rect 3402 3803 3406 3807
rect 3409 3803 3413 3807
rect 4426 3803 4430 3807
rect 4433 3803 4437 3807
rect 14 3788 18 3792
rect 46 3788 50 3792
rect 142 3788 146 3792
rect 230 3788 234 3792
rect 254 3788 258 3792
rect 278 3788 282 3792
rect 326 3788 330 3792
rect 358 3788 362 3792
rect 1054 3788 1058 3792
rect 1582 3788 1586 3792
rect 1694 3788 1698 3792
rect 2622 3788 2626 3792
rect 3158 3788 3162 3792
rect 3622 3788 3626 3792
rect 4054 3788 4058 3792
rect 4198 3788 4202 3792
rect 4318 3788 4322 3792
rect 4686 3788 4690 3792
rect 4782 3788 4786 3792
rect 5110 3788 5114 3792
rect 78 3778 82 3782
rect 2150 3778 2154 3782
rect 3270 3778 3274 3782
rect 3886 3778 3890 3782
rect 4174 3778 4178 3782
rect 54 3768 58 3772
rect 86 3768 90 3772
rect 110 3768 114 3772
rect 246 3768 250 3772
rect 630 3768 634 3772
rect 646 3768 650 3772
rect 1150 3768 1154 3772
rect 1454 3768 1458 3772
rect 1478 3768 1482 3772
rect 1750 3768 1754 3772
rect 1854 3768 1858 3772
rect 2798 3768 2802 3772
rect 3030 3768 3034 3772
rect 3054 3768 3058 3772
rect 3926 3768 3930 3772
rect 4406 3768 4410 3772
rect 4822 3768 4826 3772
rect 4998 3768 5002 3772
rect 30 3758 34 3762
rect 38 3758 42 3762
rect 78 3758 82 3762
rect 126 3758 130 3762
rect 254 3758 258 3762
rect 294 3758 298 3762
rect 390 3758 394 3762
rect 398 3758 402 3762
rect 414 3758 418 3762
rect 478 3758 482 3762
rect 942 3758 946 3762
rect 1158 3758 1162 3762
rect 1190 3758 1194 3762
rect 14 3748 18 3752
rect 46 3748 50 3752
rect 78 3748 82 3752
rect 110 3748 114 3752
rect 254 3748 258 3752
rect 278 3748 282 3752
rect 366 3748 370 3752
rect 422 3748 426 3752
rect 462 3748 466 3752
rect 470 3748 474 3752
rect 590 3748 594 3752
rect 678 3747 682 3751
rect 790 3748 794 3752
rect 854 3748 858 3752
rect 878 3748 882 3752
rect 910 3748 914 3752
rect 918 3748 922 3752
rect 934 3748 938 3752
rect 974 3747 978 3751
rect 1094 3748 1098 3752
rect 1174 3748 1178 3752
rect 1198 3748 1202 3752
rect 1206 3748 1210 3752
rect 1238 3748 1242 3752
rect 1310 3748 1314 3752
rect 1374 3748 1378 3752
rect 1398 3758 1402 3762
rect 1414 3748 1418 3752
rect 1614 3758 1618 3762
rect 1478 3748 1482 3752
rect 1518 3747 1522 3751
rect 1598 3748 1602 3752
rect 1646 3748 1650 3752
rect 1678 3748 1682 3752
rect 1718 3748 1722 3752
rect 1814 3747 1818 3751
rect 1854 3748 1858 3752
rect 1878 3758 1882 3762
rect 1950 3758 1954 3762
rect 1982 3758 1986 3762
rect 2246 3758 2250 3762
rect 2502 3758 2506 3762
rect 2566 3758 2570 3762
rect 2742 3758 2746 3762
rect 2758 3758 2762 3762
rect 2814 3758 2818 3762
rect 2822 3758 2826 3762
rect 3174 3758 3178 3762
rect 3230 3758 3234 3762
rect 3470 3758 3474 3762
rect 3790 3758 3794 3762
rect 1934 3748 1938 3752
rect 1958 3748 1962 3752
rect 1966 3748 1970 3752
rect 2030 3748 2034 3752
rect 2038 3748 2042 3752
rect 2094 3748 2098 3752
rect 2110 3748 2114 3752
rect 2126 3748 2130 3752
rect 2182 3748 2186 3752
rect 2206 3748 2210 3752
rect 2246 3748 2250 3752
rect 2270 3748 2274 3752
rect 2318 3748 2322 3752
rect 2326 3748 2330 3752
rect 2358 3748 2362 3752
rect 2430 3748 2434 3752
rect 2446 3748 2450 3752
rect 2470 3748 2474 3752
rect 2478 3748 2482 3752
rect 2510 3748 2514 3752
rect 2558 3748 2562 3752
rect 2574 3748 2578 3752
rect 2582 3748 2586 3752
rect 2630 3748 2634 3752
rect 2670 3748 2674 3752
rect 2702 3748 2706 3752
rect 2734 3748 2738 3752
rect 2766 3748 2770 3752
rect 2782 3748 2786 3752
rect 2798 3748 2802 3752
rect 2822 3748 2826 3752
rect 2838 3748 2842 3752
rect 2926 3748 2930 3752
rect 2998 3748 3002 3752
rect 3022 3748 3026 3752
rect 3086 3748 3090 3752
rect 3110 3748 3114 3752
rect 3158 3748 3162 3752
rect 3182 3748 3186 3752
rect 3214 3748 3218 3752
rect 3238 3748 3242 3752
rect 6 3738 10 3742
rect 102 3738 106 3742
rect 198 3738 202 3742
rect 206 3738 210 3742
rect 214 3740 218 3744
rect 270 3738 274 3742
rect 310 3738 314 3742
rect 374 3738 378 3742
rect 398 3738 402 3742
rect 486 3738 490 3742
rect 550 3738 554 3742
rect 566 3738 570 3742
rect 662 3738 666 3742
rect 758 3738 762 3742
rect 870 3738 874 3742
rect 918 3738 922 3742
rect 958 3738 962 3742
rect 1070 3738 1074 3742
rect 1118 3738 1122 3742
rect 1158 3738 1162 3742
rect 1182 3738 1186 3742
rect 1214 3738 1218 3742
rect 1222 3738 1226 3742
rect 1246 3738 1250 3742
rect 1302 3738 1306 3742
rect 1358 3738 1362 3742
rect 1366 3738 1370 3742
rect 1382 3738 1386 3742
rect 1422 3738 1426 3742
rect 1430 3738 1434 3742
rect 1486 3738 1490 3742
rect 1502 3738 1506 3742
rect 1638 3738 1642 3742
rect 1670 3738 1674 3742
rect 1718 3738 1722 3742
rect 1782 3738 1786 3742
rect 1830 3738 1834 3742
rect 1846 3738 1850 3742
rect 1918 3738 1922 3742
rect 1958 3738 1962 3742
rect 1982 3738 1986 3742
rect 2086 3738 2090 3742
rect 2118 3738 2122 3742
rect 2126 3738 2130 3742
rect 3334 3747 3338 3751
rect 3366 3748 3370 3752
rect 3382 3748 3386 3752
rect 3414 3748 3418 3752
rect 3470 3748 3474 3752
rect 3478 3748 3482 3752
rect 3494 3748 3498 3752
rect 3502 3748 3506 3752
rect 3526 3748 3530 3752
rect 3614 3748 3618 3752
rect 3654 3748 3658 3752
rect 3686 3747 3690 3751
rect 3718 3748 3722 3752
rect 3750 3748 3754 3752
rect 3830 3748 3834 3752
rect 3902 3748 3906 3752
rect 3910 3748 3914 3752
rect 4390 3758 4394 3762
rect 4630 3758 4634 3762
rect 4798 3758 4802 3762
rect 3958 3748 3962 3752
rect 3990 3748 3994 3752
rect 4022 3748 4026 3752
rect 4030 3748 4034 3752
rect 4038 3748 4042 3752
rect 4070 3748 4074 3752
rect 4118 3748 4122 3752
rect 4214 3748 4218 3752
rect 4270 3748 4274 3752
rect 4342 3748 4346 3752
rect 4358 3748 4362 3752
rect 4374 3748 4378 3752
rect 4398 3748 4402 3752
rect 4446 3748 4450 3752
rect 4470 3748 4474 3752
rect 4542 3748 4546 3752
rect 4558 3748 4562 3752
rect 4614 3748 4618 3752
rect 4654 3748 4658 3752
rect 4662 3748 4666 3752
rect 4726 3748 4730 3752
rect 4750 3748 4754 3752
rect 4790 3748 4794 3752
rect 4942 3758 4946 3762
rect 4838 3748 4842 3752
rect 4862 3748 4866 3752
rect 4910 3748 4914 3752
rect 4926 3748 4930 3752
rect 5094 3758 5098 3762
rect 5150 3758 5154 3762
rect 5158 3758 5162 3762
rect 4982 3748 4986 3752
rect 5038 3748 5042 3752
rect 5110 3748 5114 3752
rect 5134 3748 5138 3752
rect 5174 3748 5178 3752
rect 5222 3748 5226 3752
rect 2262 3738 2266 3742
rect 2278 3738 2282 3742
rect 2334 3738 2338 3742
rect 2366 3738 2370 3742
rect 2486 3738 2490 3742
rect 2502 3738 2506 3742
rect 2590 3738 2594 3742
rect 2598 3738 2602 3742
rect 2694 3738 2698 3742
rect 2710 3738 2714 3742
rect 2726 3738 2730 3742
rect 2742 3738 2746 3742
rect 2790 3738 2794 3742
rect 2846 3738 2850 3742
rect 2950 3738 2954 3742
rect 2982 3738 2986 3742
rect 3046 3738 3050 3742
rect 3150 3738 3154 3742
rect 3182 3738 3186 3742
rect 3206 3738 3210 3742
rect 3318 3738 3322 3742
rect 3374 3738 3378 3742
rect 3454 3738 3458 3742
rect 3494 3738 3498 3742
rect 3550 3738 3554 3742
rect 3630 3738 3634 3742
rect 3702 3738 3706 3742
rect 3726 3738 3730 3742
rect 3774 3738 3778 3742
rect 3806 3738 3810 3742
rect 3894 3738 3898 3742
rect 3966 3738 3970 3742
rect 4014 3738 4018 3742
rect 4110 3738 4114 3742
rect 4230 3738 4234 3742
rect 4334 3738 4338 3742
rect 4366 3738 4370 3742
rect 4494 3738 4498 3742
rect 4606 3738 4610 3742
rect 4622 3738 4626 3742
rect 5254 3747 5258 3751
rect 5286 3748 5290 3752
rect 4790 3738 4794 3742
rect 4846 3738 4850 3742
rect 4854 3738 4858 3742
rect 4902 3738 4906 3742
rect 4918 3738 4922 3742
rect 4974 3738 4978 3742
rect 4990 3738 4994 3742
rect 5062 3738 5066 3742
rect 5118 3738 5122 3742
rect 5126 3738 5130 3742
rect 5142 3738 5146 3742
rect 5182 3738 5186 3742
rect 302 3728 306 3732
rect 350 3728 354 3732
rect 446 3728 450 3732
rect 894 3728 898 3732
rect 1006 3728 1010 3732
rect 1630 3728 1634 3732
rect 1654 3728 1658 3732
rect 1726 3728 1730 3732
rect 1742 3728 1746 3732
rect 1766 3728 1770 3732
rect 2142 3728 2146 3732
rect 2214 3728 2218 3732
rect 2302 3728 2306 3732
rect 2350 3728 2354 3732
rect 2406 3728 2410 3732
rect 2542 3728 2546 3732
rect 2782 3728 2786 3732
rect 2966 3728 2970 3732
rect 3198 3728 3202 3732
rect 3262 3728 3266 3732
rect 3390 3728 3394 3732
rect 3398 3728 3402 3732
rect 3446 3728 3450 3732
rect 3518 3728 3522 3732
rect 3526 3728 3530 3732
rect 3542 3728 3546 3732
rect 3766 3728 3770 3732
rect 3974 3728 3978 3732
rect 3998 3728 4002 3732
rect 4182 3728 4186 3732
rect 4326 3728 4330 3732
rect 4358 3728 4362 3732
rect 4638 3728 4642 3732
rect 4654 3728 4658 3732
rect 4686 3728 4690 3732
rect 4886 3728 4890 3732
rect 5222 3728 5226 3732
rect 5302 3728 5306 3732
rect 742 3718 746 3722
rect 838 3718 842 3722
rect 1254 3718 1258 3722
rect 1662 3718 1666 3722
rect 1990 3718 1994 3722
rect 2110 3718 2114 3722
rect 2286 3718 2290 3722
rect 2342 3718 2346 3722
rect 2374 3718 2378 3722
rect 2494 3718 2498 3722
rect 2526 3718 2530 3722
rect 2654 3718 2658 3722
rect 2710 3718 2714 3722
rect 2870 3718 2874 3722
rect 2974 3718 2978 3722
rect 3030 3718 3034 3722
rect 3254 3718 3258 3722
rect 3510 3718 3514 3722
rect 3734 3718 3738 3722
rect 3782 3718 3786 3722
rect 3982 3718 3986 3722
rect 4006 3718 4010 3722
rect 4166 3718 4170 3722
rect 4310 3718 4314 3722
rect 4318 3718 4322 3722
rect 4398 3718 4402 3722
rect 4510 3718 4514 3722
rect 4878 3718 4882 3722
rect 4894 3718 4898 3722
rect 5158 3718 5162 3722
rect 5294 3718 5298 3722
rect 850 3703 854 3707
rect 857 3703 861 3707
rect 1874 3703 1878 3707
rect 1881 3703 1885 3707
rect 2890 3703 2894 3707
rect 2897 3703 2901 3707
rect 3922 3703 3926 3707
rect 3929 3703 3933 3707
rect 4938 3703 4942 3707
rect 4945 3703 4949 3707
rect 22 3688 26 3692
rect 70 3688 74 3692
rect 94 3688 98 3692
rect 190 3688 194 3692
rect 222 3688 226 3692
rect 406 3688 410 3692
rect 430 3688 434 3692
rect 470 3688 474 3692
rect 646 3688 650 3692
rect 878 3688 882 3692
rect 1110 3688 1114 3692
rect 1142 3688 1146 3692
rect 1190 3688 1194 3692
rect 1262 3688 1266 3692
rect 1310 3688 1314 3692
rect 1550 3688 1554 3692
rect 1670 3688 1674 3692
rect 1958 3688 1962 3692
rect 2014 3688 2018 3692
rect 2038 3688 2042 3692
rect 2278 3688 2282 3692
rect 2374 3688 2378 3692
rect 2406 3688 2410 3692
rect 2422 3688 2426 3692
rect 2662 3688 2666 3692
rect 2798 3688 2802 3692
rect 3094 3688 3098 3692
rect 3286 3688 3290 3692
rect 3526 3688 3530 3692
rect 3758 3688 3762 3692
rect 3782 3688 3786 3692
rect 3950 3688 3954 3692
rect 4118 3688 4122 3692
rect 4214 3688 4218 3692
rect 4382 3688 4386 3692
rect 4542 3688 4546 3692
rect 4558 3688 4562 3692
rect 4702 3688 4706 3692
rect 4718 3688 4722 3692
rect 4862 3688 4866 3692
rect 5254 3688 5258 3692
rect 30 3678 34 3682
rect 62 3678 66 3682
rect 142 3678 146 3682
rect 198 3678 202 3682
rect 14 3668 18 3672
rect 38 3668 42 3672
rect 102 3668 106 3672
rect 110 3668 114 3672
rect 126 3668 130 3672
rect 150 3668 154 3672
rect 182 3668 186 3672
rect 214 3668 218 3672
rect 462 3678 466 3682
rect 566 3678 570 3682
rect 678 3678 682 3682
rect 750 3678 754 3682
rect 318 3668 322 3672
rect 326 3668 330 3672
rect 398 3668 402 3672
rect 422 3668 426 3672
rect 582 3668 586 3672
rect 590 3668 594 3672
rect 638 3668 642 3672
rect 1238 3678 1242 3682
rect 1270 3678 1274 3682
rect 1766 3678 1770 3682
rect 1838 3678 1842 3682
rect 1918 3678 1922 3682
rect 1998 3678 2002 3682
rect 774 3668 778 3672
rect 798 3668 802 3672
rect 846 3668 850 3672
rect 942 3668 946 3672
rect 958 3668 962 3672
rect 974 3668 978 3672
rect 1014 3668 1018 3672
rect 1030 3668 1034 3672
rect 1070 3668 1074 3672
rect 1118 3668 1122 3672
rect 1150 3668 1154 3672
rect 1254 3668 1258 3672
rect 1278 3668 1282 3672
rect 1294 3668 1298 3672
rect 1358 3668 1362 3672
rect 1406 3668 1410 3672
rect 1478 3668 1482 3672
rect 1510 3668 1514 3672
rect 1566 3668 1570 3672
rect 1574 3668 1578 3672
rect 1630 3668 1634 3672
rect 1662 3668 1666 3672
rect 1750 3668 1754 3672
rect 1814 3668 1818 3672
rect 1910 3668 1914 3672
rect 1950 3668 1954 3672
rect 2078 3678 2082 3682
rect 2214 3678 2218 3682
rect 2246 3678 2250 3682
rect 2494 3678 2498 3682
rect 2654 3678 2658 3682
rect 2726 3678 2730 3682
rect 2830 3678 2834 3682
rect 2974 3678 2978 3682
rect 2982 3678 2986 3682
rect 3342 3678 3346 3682
rect 2022 3668 2026 3672
rect 2094 3668 2098 3672
rect 2110 3668 2114 3672
rect 2134 3668 2138 3672
rect 2150 3668 2154 3672
rect 2294 3668 2298 3672
rect 2414 3668 2418 3672
rect 2446 3668 2450 3672
rect 2454 3668 2458 3672
rect 2518 3668 2522 3672
rect 2550 3668 2554 3672
rect 2582 3668 2586 3672
rect 2590 3668 2594 3672
rect 2686 3668 2690 3672
rect 2694 3668 2698 3672
rect 2782 3668 2786 3672
rect 2790 3668 2794 3672
rect 6 3658 10 3662
rect 54 3658 58 3662
rect 78 3658 82 3662
rect 118 3658 122 3662
rect 174 3658 178 3662
rect 206 3658 210 3662
rect 262 3658 266 3662
rect 398 3658 402 3662
rect 414 3658 418 3662
rect 446 3658 450 3662
rect 502 3658 506 3662
rect 526 3658 530 3662
rect 590 3658 594 3662
rect 614 3658 618 3662
rect 622 3658 626 3662
rect 630 3658 634 3662
rect 662 3658 666 3662
rect 686 3658 690 3662
rect 702 3658 706 3662
rect 718 3658 722 3662
rect 726 3658 730 3662
rect 734 3658 738 3662
rect 766 3658 770 3662
rect 782 3658 786 3662
rect 814 3659 818 3663
rect 926 3658 930 3662
rect 950 3658 954 3662
rect 966 3658 970 3662
rect 998 3658 1002 3662
rect 1046 3659 1050 3663
rect 1126 3658 1130 3662
rect 1158 3658 1162 3662
rect 1190 3658 1194 3662
rect 1206 3658 1210 3662
rect 1222 3658 1226 3662
rect 1246 3658 1250 3662
rect 1286 3658 1290 3662
rect 1374 3659 1378 3663
rect 1430 3658 1434 3662
rect 1438 3658 1442 3662
rect 1470 3658 1474 3662
rect 1502 3658 1506 3662
rect 1542 3658 1546 3662
rect 1582 3658 1586 3662
rect 1622 3658 1626 3662
rect 1654 3658 1658 3662
rect 1726 3658 1730 3662
rect 1790 3658 1794 3662
rect 1870 3658 1874 3662
rect 1902 3658 1906 3662
rect 1934 3658 1938 3662
rect 1974 3658 1978 3662
rect 1982 3658 1986 3662
rect 2030 3658 2034 3662
rect 2054 3658 2058 3662
rect 2086 3658 2090 3662
rect 2118 3658 2122 3662
rect 2126 3658 2130 3662
rect 2142 3658 2146 3662
rect 2182 3658 2186 3662
rect 2222 3658 2226 3662
rect 2318 3658 2322 3662
rect 2438 3658 2442 3662
rect 2462 3658 2466 3662
rect 2494 3658 2498 3662
rect 2542 3658 2546 3662
rect 2574 3658 2578 3662
rect 2598 3658 2602 3662
rect 2622 3658 2626 3662
rect 2630 3658 2634 3662
rect 2638 3658 2642 3662
rect 2678 3658 2682 3662
rect 2702 3658 2706 3662
rect 2718 3658 2722 3662
rect 2742 3658 2746 3662
rect 2766 3658 2770 3662
rect 2774 3658 2778 3662
rect 2814 3658 2818 3662
rect 2838 3658 2842 3662
rect 2854 3658 2858 3662
rect 2870 3668 2874 3672
rect 2918 3668 2922 3672
rect 2958 3668 2962 3672
rect 2974 3668 2978 3672
rect 2982 3668 2986 3672
rect 3038 3668 3042 3672
rect 3086 3668 3090 3672
rect 3190 3668 3194 3672
rect 3206 3668 3210 3672
rect 3238 3668 3242 3672
rect 3334 3668 3338 3672
rect 3462 3668 3466 3672
rect 3518 3668 3522 3672
rect 3566 3668 3570 3672
rect 3598 3668 3602 3672
rect 3790 3678 3794 3682
rect 3830 3678 3834 3682
rect 4206 3678 4210 3682
rect 4398 3678 4402 3682
rect 4406 3678 4410 3682
rect 4414 3678 4418 3682
rect 4446 3678 4450 3682
rect 4550 3678 4554 3682
rect 4590 3678 4594 3682
rect 4614 3678 4618 3682
rect 4662 3678 4666 3682
rect 4678 3678 4682 3682
rect 4814 3678 4818 3682
rect 5246 3678 5250 3682
rect 5278 3678 5282 3682
rect 3622 3668 3626 3672
rect 2870 3658 2874 3662
rect 2878 3658 2882 3662
rect 2926 3658 2930 3662
rect 2950 3658 2954 3662
rect 3006 3658 3010 3662
rect 3030 3658 3034 3662
rect 3046 3658 3050 3662
rect 3054 3658 3058 3662
rect 3142 3658 3146 3662
rect 3166 3658 3170 3662
rect 3214 3658 3218 3662
rect 3230 3658 3234 3662
rect 3270 3658 3274 3662
rect 3302 3658 3306 3662
rect 3326 3658 3330 3662
rect 3390 3658 3394 3662
rect 3422 3659 3426 3663
rect 3662 3668 3666 3672
rect 3694 3668 3698 3672
rect 3702 3668 3706 3672
rect 3774 3668 3778 3672
rect 3822 3668 3826 3672
rect 3854 3668 3858 3672
rect 3894 3668 3898 3672
rect 3974 3668 3978 3672
rect 4006 3668 4010 3672
rect 4038 3668 4042 3672
rect 4086 3668 4090 3672
rect 4166 3668 4170 3672
rect 4198 3668 4202 3672
rect 4222 3668 4226 3672
rect 4262 3668 4266 3672
rect 4318 3668 4322 3672
rect 4334 3668 4338 3672
rect 4366 3668 4370 3672
rect 4462 3668 4466 3672
rect 4566 3668 4570 3672
rect 4630 3668 4634 3672
rect 4766 3668 4770 3672
rect 4838 3668 4842 3672
rect 4878 3668 4882 3672
rect 5022 3668 5026 3672
rect 5078 3668 5082 3672
rect 5142 3668 5146 3672
rect 5262 3668 5266 3672
rect 3478 3658 3482 3662
rect 3502 3658 3506 3662
rect 3510 3658 3514 3662
rect 3558 3658 3562 3662
rect 3574 3658 3578 3662
rect 3614 3658 3618 3662
rect 3630 3658 3634 3662
rect 3638 3658 3642 3662
rect 3654 3658 3658 3662
rect 3710 3658 3714 3662
rect 3766 3658 3770 3662
rect 3822 3658 3826 3662
rect 3846 3658 3850 3662
rect 3910 3658 3914 3662
rect 3966 3658 3970 3662
rect 4014 3658 4018 3662
rect 4062 3658 4066 3662
rect 4094 3658 4098 3662
rect 4102 3658 4106 3662
rect 4134 3658 4138 3662
rect 4158 3658 4162 3662
rect 4190 3658 4194 3662
rect 4230 3658 4234 3662
rect 4238 3658 4242 3662
rect 4254 3658 4258 3662
rect 4270 3658 4274 3662
rect 4278 3658 4282 3662
rect 4302 3658 4306 3662
rect 4358 3658 4362 3662
rect 4366 3658 4370 3662
rect 4398 3658 4402 3662
rect 4414 3658 4418 3662
rect 4478 3659 4482 3663
rect 4574 3658 4578 3662
rect 4606 3658 4610 3662
rect 4638 3658 4642 3662
rect 4646 3658 4650 3662
rect 4686 3658 4690 3662
rect 4774 3658 4778 3662
rect 4838 3658 4842 3662
rect 4846 3658 4850 3662
rect 4886 3658 4890 3662
rect 4958 3658 4962 3662
rect 4990 3659 4994 3663
rect 5030 3658 5034 3662
rect 5038 3658 5042 3662
rect 5078 3658 5082 3662
rect 5134 3658 5138 3662
rect 5182 3658 5186 3662
rect 5206 3658 5210 3662
rect 5278 3658 5282 3662
rect 5294 3658 5298 3662
rect 54 3648 58 3652
rect 86 3648 90 3652
rect 134 3648 138 3652
rect 934 3648 938 3652
rect 1142 3648 1146 3652
rect 1174 3648 1178 3652
rect 1302 3648 1306 3652
rect 1454 3648 1458 3652
rect 1550 3648 1554 3652
rect 1582 3648 1586 3652
rect 1598 3648 1602 3652
rect 1606 3648 1610 3652
rect 1622 3648 1626 3652
rect 1638 3648 1642 3652
rect 1830 3648 1834 3652
rect 1886 3648 1890 3652
rect 1918 3648 1922 3652
rect 2038 3648 2042 3652
rect 2390 3648 2394 3652
rect 2422 3648 2426 3652
rect 2478 3648 2482 3652
rect 2526 3648 2530 3652
rect 2646 3648 2650 3652
rect 2662 3648 2666 3652
rect 2702 3648 2706 3652
rect 2718 3648 2722 3652
rect 2750 3648 2754 3652
rect 2838 3648 2842 3652
rect 2894 3648 2898 3652
rect 2926 3648 2930 3652
rect 2942 3648 2946 3652
rect 3014 3648 3018 3652
rect 3310 3648 3314 3652
rect 3534 3648 3538 3652
rect 3638 3648 3642 3652
rect 3798 3648 3802 3652
rect 3830 3648 3834 3652
rect 3998 3648 4002 3652
rect 4014 3648 4018 3652
rect 4038 3648 4042 3652
rect 4054 3648 4058 3652
rect 4142 3648 4146 3652
rect 4174 3648 4178 3652
rect 4238 3648 4242 3652
rect 4318 3648 4322 3652
rect 4902 3648 4906 3652
rect 5054 3648 5058 3652
rect 5134 3648 5138 3652
rect 910 3638 914 3642
rect 1486 3638 1490 3642
rect 1654 3638 1658 3642
rect 3590 3638 3594 3642
rect 4158 3638 4162 3642
rect 5110 3638 5114 3642
rect 5150 3638 5154 3642
rect 3982 3628 3986 3632
rect 4046 3628 4050 3632
rect 246 3618 250 3622
rect 294 3618 298 3622
rect 894 3618 898 3622
rect 990 3618 994 3622
rect 1502 3618 1506 3622
rect 1790 3618 1794 3622
rect 1838 3618 1842 3622
rect 2110 3618 2114 3622
rect 2558 3618 2562 3622
rect 2766 3618 2770 3622
rect 2878 3618 2882 3622
rect 3214 3618 3218 3622
rect 3254 3618 3258 3622
rect 3326 3618 3330 3622
rect 3542 3618 3546 3622
rect 3814 3618 3818 3622
rect 4078 3618 4082 3622
rect 4190 3618 4194 3622
rect 4358 3618 4362 3622
rect 4614 3618 4618 3622
rect 4646 3618 4650 3622
rect 4670 3618 4674 3622
rect 4702 3618 4706 3622
rect 4814 3618 4818 3622
rect 4886 3618 4890 3622
rect 4926 3618 4930 3622
rect 5286 3618 5290 3622
rect 330 3603 334 3607
rect 337 3603 341 3607
rect 1354 3603 1358 3607
rect 1361 3603 1365 3607
rect 2386 3603 2390 3607
rect 2393 3603 2397 3607
rect 3402 3603 3406 3607
rect 3409 3603 3413 3607
rect 4426 3603 4430 3607
rect 4433 3603 4437 3607
rect 950 3588 954 3592
rect 1054 3588 1058 3592
rect 1150 3588 1154 3592
rect 1166 3588 1170 3592
rect 1334 3588 1338 3592
rect 1462 3588 1466 3592
rect 2534 3588 2538 3592
rect 2678 3588 2682 3592
rect 2974 3588 2978 3592
rect 3022 3588 3026 3592
rect 3062 3588 3066 3592
rect 3246 3588 3250 3592
rect 3478 3588 3482 3592
rect 4446 3588 4450 3592
rect 4662 3588 4666 3592
rect 5150 3588 5154 3592
rect 5166 3588 5170 3592
rect 2510 3578 2514 3582
rect 3990 3578 3994 3582
rect 486 3568 490 3572
rect 758 3568 762 3572
rect 790 3568 794 3572
rect 1022 3568 1026 3572
rect 1190 3568 1194 3572
rect 1214 3568 1218 3572
rect 1750 3568 1754 3572
rect 1766 3568 1770 3572
rect 2686 3568 2690 3572
rect 2830 3568 2834 3572
rect 2958 3568 2962 3572
rect 3174 3568 3178 3572
rect 3670 3568 3674 3572
rect 3950 3568 3954 3572
rect 4558 3568 4562 3572
rect 102 3558 106 3562
rect 390 3558 394 3562
rect 550 3558 554 3562
rect 566 3558 570 3562
rect 70 3547 74 3551
rect 126 3548 130 3552
rect 150 3548 154 3552
rect 158 3548 162 3552
rect 206 3548 210 3552
rect 262 3548 266 3552
rect 86 3538 90 3542
rect 118 3538 122 3542
rect 174 3538 178 3542
rect 198 3538 202 3542
rect 286 3538 290 3542
rect 326 3548 330 3552
rect 342 3548 346 3552
rect 430 3548 434 3552
rect 494 3548 498 3552
rect 510 3548 514 3552
rect 526 3548 530 3552
rect 566 3548 570 3552
rect 590 3548 594 3552
rect 614 3548 618 3552
rect 622 3548 626 3552
rect 702 3548 706 3552
rect 774 3548 778 3552
rect 990 3558 994 3562
rect 1158 3558 1162 3562
rect 814 3548 818 3552
rect 830 3548 834 3552
rect 886 3548 890 3552
rect 918 3548 922 3552
rect 974 3548 978 3552
rect 1006 3548 1010 3552
rect 1038 3548 1042 3552
rect 1054 3548 1058 3552
rect 1102 3548 1106 3552
rect 1190 3548 1194 3552
rect 1230 3548 1234 3552
rect 1286 3548 1290 3552
rect 1342 3548 1346 3552
rect 1390 3558 1394 3562
rect 1446 3558 1450 3562
rect 1454 3558 1458 3562
rect 1526 3558 1530 3562
rect 1582 3558 1586 3562
rect 1654 3558 1658 3562
rect 1782 3558 1786 3562
rect 2110 3558 2114 3562
rect 2174 3558 2178 3562
rect 2246 3558 2250 3562
rect 2278 3558 2282 3562
rect 1422 3548 1426 3552
rect 1430 3548 1434 3552
rect 1478 3548 1482 3552
rect 1510 3548 1514 3552
rect 1558 3548 1562 3552
rect 1566 3548 1570 3552
rect 1598 3548 1602 3552
rect 1606 3548 1610 3552
rect 1622 3548 1626 3552
rect 1638 3548 1642 3552
rect 1694 3548 1698 3552
rect 1766 3548 1770 3552
rect 1806 3548 1810 3552
rect 1846 3548 1850 3552
rect 1902 3548 1906 3552
rect 1982 3548 1986 3552
rect 2006 3548 2010 3552
rect 2014 3548 2018 3552
rect 2022 3548 2026 3552
rect 2054 3548 2058 3552
rect 2086 3548 2090 3552
rect 2126 3548 2130 3552
rect 2142 3548 2146 3552
rect 2174 3548 2178 3552
rect 2190 3548 2194 3552
rect 2214 3548 2218 3552
rect 2230 3548 2234 3552
rect 2246 3548 2250 3552
rect 2262 3548 2266 3552
rect 2294 3548 2298 3552
rect 2302 3548 2306 3552
rect 2342 3548 2346 3552
rect 2350 3548 2354 3552
rect 2374 3548 2378 3552
rect 2438 3548 2442 3552
rect 2518 3548 2522 3552
rect 2590 3558 2594 3562
rect 2606 3558 2610 3562
rect 2638 3558 2642 3562
rect 2566 3548 2570 3552
rect 2590 3548 2594 3552
rect 2622 3548 2626 3552
rect 2814 3558 2818 3562
rect 2846 3558 2850 3562
rect 2990 3558 2994 3562
rect 3054 3558 3058 3562
rect 3158 3558 3162 3562
rect 3190 3558 3194 3562
rect 3462 3558 3466 3562
rect 3550 3558 3554 3562
rect 3702 3558 3706 3562
rect 3758 3558 3762 3562
rect 3974 3558 3978 3562
rect 4006 3558 4010 3562
rect 4022 3558 4026 3562
rect 4038 3558 4042 3562
rect 4350 3558 4354 3562
rect 4486 3558 4490 3562
rect 4502 3558 4506 3562
rect 4518 3558 4522 3562
rect 4534 3558 4538 3562
rect 4542 3558 4546 3562
rect 4574 3558 4578 3562
rect 4694 3558 4698 3562
rect 4910 3558 4914 3562
rect 5006 3558 5010 3562
rect 5134 3558 5138 3562
rect 2654 3548 2658 3552
rect 2662 3548 2666 3552
rect 2750 3548 2754 3552
rect 2798 3548 2802 3552
rect 2814 3548 2818 3552
rect 2830 3548 2834 3552
rect 302 3538 306 3542
rect 366 3538 370 3542
rect 406 3538 410 3542
rect 502 3538 506 3542
rect 582 3538 586 3542
rect 662 3538 666 3542
rect 678 3538 682 3542
rect 766 3538 770 3542
rect 798 3538 802 3542
rect 822 3538 826 3542
rect 862 3538 866 3542
rect 910 3538 914 3542
rect 926 3538 930 3542
rect 966 3538 970 3542
rect 1030 3538 1034 3542
rect 1070 3538 1074 3542
rect 1174 3538 1178 3542
rect 1182 3538 1186 3542
rect 1238 3538 1242 3542
rect 1278 3538 1282 3542
rect 1342 3538 1346 3542
rect 1414 3538 1418 3542
rect 1422 3538 1426 3542
rect 1470 3538 1474 3542
rect 1478 3538 1482 3542
rect 1494 3538 1498 3542
rect 1534 3538 1538 3542
rect 1550 3538 1554 3542
rect 1590 3538 1594 3542
rect 1622 3538 1626 3542
rect 1630 3538 1634 3542
rect 1670 3538 1674 3542
rect 1758 3538 1762 3542
rect 1814 3538 1818 3542
rect 1830 3538 1834 3542
rect 1894 3538 1898 3542
rect 1974 3538 1978 3542
rect 2030 3538 2034 3542
rect 2054 3538 2058 3542
rect 2062 3538 2066 3542
rect 2134 3538 2138 3542
rect 2150 3538 2154 3542
rect 2198 3538 2202 3542
rect 2206 3538 2210 3542
rect 2238 3538 2242 3542
rect 2302 3538 2306 3542
rect 2326 3540 2330 3544
rect 2334 3538 2338 3542
rect 2398 3538 2402 3542
rect 2446 3538 2450 3542
rect 2550 3538 2554 3542
rect 2574 3538 2578 3542
rect 2582 3538 2586 3542
rect 2614 3538 2618 3542
rect 2670 3538 2674 3542
rect 2774 3538 2778 3542
rect 2790 3538 2794 3542
rect 2894 3547 2898 3551
rect 2926 3548 2930 3552
rect 2974 3548 2978 3552
rect 2998 3548 3002 3552
rect 3030 3548 3034 3552
rect 3054 3548 3058 3552
rect 3126 3547 3130 3551
rect 3174 3548 3178 3552
rect 3190 3548 3194 3552
rect 3206 3548 3210 3552
rect 3238 3548 3242 3552
rect 3326 3547 3330 3551
rect 3366 3548 3370 3552
rect 3390 3548 3394 3552
rect 3398 3548 3402 3552
rect 3422 3548 3426 3552
rect 3454 3548 3458 3552
rect 3478 3548 3482 3552
rect 3494 3548 3498 3552
rect 3502 3548 3506 3552
rect 3526 3548 3530 3552
rect 3606 3548 3610 3552
rect 3686 3548 3690 3552
rect 3726 3548 3730 3552
rect 3734 3548 3738 3552
rect 3806 3548 3810 3552
rect 3886 3547 3890 3551
rect 3990 3548 3994 3552
rect 4030 3548 4034 3552
rect 4054 3548 4058 3552
rect 4070 3548 4074 3552
rect 4086 3548 4090 3552
rect 4102 3548 4106 3552
rect 4118 3548 4122 3552
rect 4158 3548 4162 3552
rect 4166 3548 4170 3552
rect 4182 3548 4186 3552
rect 4198 3548 4202 3552
rect 4214 3548 4218 3552
rect 4262 3548 4266 3552
rect 4326 3548 4330 3552
rect 4366 3548 4370 3552
rect 4406 3548 4410 3552
rect 4414 3548 4418 3552
rect 4462 3548 4466 3552
rect 4470 3548 4474 3552
rect 4486 3548 4490 3552
rect 4518 3548 4522 3552
rect 4558 3548 4562 3552
rect 4598 3548 4602 3552
rect 4630 3548 4634 3552
rect 4638 3548 4642 3552
rect 4646 3548 4650 3552
rect 4670 3548 4674 3552
rect 4734 3548 4738 3552
rect 4742 3548 4746 3552
rect 4758 3548 4762 3552
rect 4870 3548 4874 3552
rect 4926 3548 4930 3552
rect 4982 3548 4986 3552
rect 5030 3548 5034 3552
rect 5094 3548 5098 3552
rect 5158 3548 5162 3552
rect 5246 3547 5250 3551
rect 5278 3548 5282 3552
rect 2822 3538 2826 3542
rect 2854 3538 2858 3542
rect 2966 3538 2970 3542
rect 3006 3538 3010 3542
rect 3030 3538 3034 3542
rect 3102 3538 3106 3542
rect 3142 3538 3146 3542
rect 3182 3538 3186 3542
rect 3214 3538 3218 3542
rect 3318 3538 3322 3542
rect 3358 3538 3362 3542
rect 3430 3538 3434 3542
rect 3446 3538 3450 3542
rect 3486 3538 3490 3542
rect 3534 3538 3538 3542
rect 3638 3538 3642 3542
rect 3654 3538 3658 3542
rect 3678 3538 3682 3542
rect 3710 3538 3714 3542
rect 3774 3538 3778 3542
rect 3894 3538 3898 3542
rect 3998 3538 4002 3542
rect 4030 3538 4034 3542
rect 4046 3538 4050 3542
rect 4062 3538 4066 3542
rect 4094 3538 4098 3542
rect 4126 3538 4130 3542
rect 4190 3538 4194 3542
rect 4222 3538 4226 3542
rect 4270 3538 4274 3542
rect 4374 3538 4378 3542
rect 4398 3538 4402 3542
rect 4478 3538 4482 3542
rect 4510 3538 4514 3542
rect 4566 3538 4570 3542
rect 4590 3538 4594 3542
rect 4606 3538 4610 3542
rect 4622 3538 4626 3542
rect 4790 3538 4794 3542
rect 4894 3538 4898 3542
rect 4918 3538 4922 3542
rect 4934 3538 4938 3542
rect 4974 3538 4978 3542
rect 4990 3538 4994 3542
rect 5094 3538 5098 3542
rect 5158 3538 5162 3542
rect 5286 3538 5290 3542
rect 70 3528 74 3532
rect 102 3528 106 3532
rect 310 3528 314 3532
rect 342 3528 346 3532
rect 390 3528 394 3532
rect 542 3528 546 3532
rect 846 3528 850 3532
rect 870 3528 874 3532
rect 902 3528 906 3532
rect 1038 3528 1042 3532
rect 1494 3528 1498 3532
rect 1534 3528 1538 3532
rect 1790 3528 1794 3532
rect 1990 3528 1994 3532
rect 2046 3528 2050 3532
rect 2102 3528 2106 3532
rect 3022 3528 3026 3532
rect 3222 3528 3226 3532
rect 3326 3528 3330 3532
rect 3710 3528 3714 3532
rect 4086 3528 4090 3532
rect 4166 3528 4170 3532
rect 4342 3528 4346 3532
rect 4382 3528 4386 3532
rect 4574 3528 4578 3532
rect 4606 3528 4610 3532
rect 4694 3528 4698 3532
rect 4950 3528 4954 3532
rect 5014 3528 5018 3532
rect 5246 3528 5250 3532
rect 5302 3528 5306 3532
rect 6 3518 10 3522
rect 254 3518 258 3522
rect 606 3518 610 3522
rect 654 3518 658 3522
rect 934 3518 938 3522
rect 1366 3518 1370 3522
rect 1446 3518 1450 3522
rect 1542 3518 1546 3522
rect 1582 3518 1586 3522
rect 1654 3518 1658 3522
rect 2070 3518 2074 3522
rect 2110 3518 2114 3522
rect 2214 3518 2218 3522
rect 3230 3518 3234 3522
rect 3438 3518 3442 3522
rect 3662 3518 3666 3522
rect 3758 3518 3762 3522
rect 3854 3518 3858 3522
rect 4118 3518 4122 3522
rect 4142 3518 4146 3522
rect 4214 3518 4218 3522
rect 4318 3518 4322 3522
rect 4334 3518 4338 3522
rect 4350 3518 4354 3522
rect 4390 3518 4394 3522
rect 4726 3518 4730 3522
rect 4814 3518 4818 3522
rect 5038 3518 5042 3522
rect 5182 3518 5186 3522
rect 5294 3518 5298 3522
rect 850 3503 854 3507
rect 857 3503 861 3507
rect 1874 3503 1878 3507
rect 1881 3503 1885 3507
rect 2890 3503 2894 3507
rect 2897 3503 2901 3507
rect 3922 3503 3926 3507
rect 3929 3503 3933 3507
rect 4938 3503 4942 3507
rect 4945 3503 4949 3507
rect 94 3488 98 3492
rect 158 3488 162 3492
rect 438 3488 442 3492
rect 478 3488 482 3492
rect 582 3488 586 3492
rect 814 3488 818 3492
rect 830 3488 834 3492
rect 878 3488 882 3492
rect 902 3488 906 3492
rect 1070 3488 1074 3492
rect 1094 3488 1098 3492
rect 1294 3488 1298 3492
rect 1390 3488 1394 3492
rect 1502 3488 1506 3492
rect 1542 3488 1546 3492
rect 1606 3488 1610 3492
rect 1710 3488 1714 3492
rect 1758 3488 1762 3492
rect 2014 3488 2018 3492
rect 2038 3488 2042 3492
rect 2134 3488 2138 3492
rect 2150 3488 2154 3492
rect 2334 3488 2338 3492
rect 2358 3488 2362 3492
rect 2374 3488 2378 3492
rect 2838 3488 2842 3492
rect 3006 3488 3010 3492
rect 3158 3488 3162 3492
rect 3182 3488 3186 3492
rect 3526 3488 3530 3492
rect 3590 3488 3594 3492
rect 3766 3488 3770 3492
rect 3806 3488 3810 3492
rect 3958 3488 3962 3492
rect 3990 3488 3994 3492
rect 4022 3488 4026 3492
rect 4198 3488 4202 3492
rect 4262 3488 4266 3492
rect 4310 3488 4314 3492
rect 4342 3488 4346 3492
rect 4670 3488 4674 3492
rect 4718 3488 4722 3492
rect 198 3478 202 3482
rect 574 3478 578 3482
rect 822 3478 826 3482
rect 894 3478 898 3482
rect 1598 3478 1602 3482
rect 126 3468 130 3472
rect 270 3468 274 3472
rect 294 3468 298 3472
rect 342 3468 346 3472
rect 446 3468 450 3472
rect 502 3468 506 3472
rect 510 3468 514 3472
rect 526 3468 530 3472
rect 566 3468 570 3472
rect 678 3468 682 3472
rect 6 3458 10 3462
rect 166 3458 170 3462
rect 206 3458 210 3462
rect 286 3458 290 3462
rect 302 3458 306 3462
rect 318 3458 322 3462
rect 382 3458 386 3462
rect 406 3458 410 3462
rect 454 3458 458 3462
rect 494 3458 498 3462
rect 518 3458 522 3462
rect 558 3458 562 3462
rect 590 3458 594 3462
rect 662 3459 666 3463
rect 718 3468 722 3472
rect 918 3468 922 3472
rect 974 3468 978 3472
rect 1118 3468 1122 3472
rect 1206 3468 1210 3472
rect 1238 3468 1242 3472
rect 1262 3468 1266 3472
rect 1270 3468 1274 3472
rect 1310 3468 1314 3472
rect 1446 3468 1450 3472
rect 1510 3468 1514 3472
rect 1558 3468 1562 3472
rect 1590 3468 1594 3472
rect 1630 3468 1634 3472
rect 1670 3468 1674 3472
rect 1750 3468 1754 3472
rect 1774 3468 1778 3472
rect 1790 3468 1794 3472
rect 1862 3468 1866 3472
rect 1902 3478 1906 3482
rect 2214 3478 2218 3482
rect 2502 3478 2506 3482
rect 2518 3478 2522 3482
rect 2630 3478 2634 3482
rect 2982 3478 2986 3482
rect 3406 3478 3410 3482
rect 3550 3478 3554 3482
rect 3566 3478 3570 3482
rect 3846 3478 3850 3482
rect 3862 3478 3866 3482
rect 3894 3478 3898 3482
rect 3998 3478 4002 3482
rect 4294 3478 4298 3482
rect 4350 3478 4354 3482
rect 4926 3478 4930 3482
rect 4974 3478 4978 3482
rect 1934 3468 1938 3472
rect 1966 3468 1970 3472
rect 2158 3468 2162 3472
rect 2310 3468 2314 3472
rect 2326 3468 2330 3472
rect 2350 3468 2354 3472
rect 2534 3468 2538 3472
rect 2638 3468 2642 3472
rect 2686 3468 2690 3472
rect 2726 3468 2730 3472
rect 2814 3468 2818 3472
rect 2870 3468 2874 3472
rect 2878 3468 2882 3472
rect 2950 3468 2954 3472
rect 3102 3468 3106 3472
rect 3166 3468 3170 3472
rect 3206 3468 3210 3472
rect 3238 3468 3242 3472
rect 3278 3468 3282 3472
rect 3326 3468 3330 3472
rect 3518 3468 3522 3472
rect 3542 3468 3546 3472
rect 3574 3468 3578 3472
rect 3606 3468 3610 3472
rect 3622 3468 3626 3472
rect 3782 3468 3786 3472
rect 4046 3468 4050 3472
rect 4062 3468 4066 3472
rect 4174 3468 4178 3472
rect 4190 3468 4194 3472
rect 4238 3468 4242 3472
rect 4254 3468 4258 3472
rect 4302 3468 4306 3472
rect 4334 3468 4338 3472
rect 4366 3468 4370 3472
rect 4470 3468 4474 3472
rect 4486 3468 4490 3472
rect 4582 3468 4586 3472
rect 4606 3468 4610 3472
rect 4622 3468 4626 3472
rect 4662 3468 4666 3472
rect 4710 3468 4714 3472
rect 4766 3468 4770 3472
rect 4798 3468 4802 3472
rect 4982 3468 4986 3472
rect 5006 3468 5010 3472
rect 5038 3468 5042 3472
rect 5094 3468 5098 3472
rect 5126 3468 5130 3472
rect 5174 3468 5178 3472
rect 5246 3468 5250 3472
rect 694 3458 698 3462
rect 710 3458 714 3462
rect 766 3458 770 3462
rect 774 3458 778 3462
rect 838 3458 842 3462
rect 862 3458 866 3462
rect 910 3458 914 3462
rect 926 3458 930 3462
rect 958 3458 962 3462
rect 966 3458 970 3462
rect 1006 3459 1010 3463
rect 1038 3458 1042 3462
rect 1078 3458 1082 3462
rect 1142 3458 1146 3462
rect 1214 3458 1218 3462
rect 1254 3458 1258 3462
rect 1278 3458 1282 3462
rect 1334 3458 1338 3462
rect 1454 3458 1458 3462
rect 1510 3458 1514 3462
rect 1582 3458 1586 3462
rect 1614 3458 1618 3462
rect 1646 3459 1650 3463
rect 1726 3458 1730 3462
rect 1782 3458 1786 3462
rect 1814 3458 1818 3462
rect 1838 3458 1842 3462
rect 1846 3458 1850 3462
rect 1854 3458 1858 3462
rect 1894 3458 1898 3462
rect 1918 3458 1922 3462
rect 1950 3459 1954 3463
rect 2038 3458 2042 3462
rect 2070 3459 2074 3463
rect 2102 3458 2106 3462
rect 2166 3458 2170 3462
rect 2198 3458 2202 3462
rect 2206 3458 2210 3462
rect 2286 3458 2290 3462
rect 2438 3458 2442 3462
rect 2462 3458 2466 3462
rect 2502 3458 2506 3462
rect 2558 3458 2562 3462
rect 2582 3458 2586 3462
rect 2670 3458 2674 3462
rect 2678 3458 2682 3462
rect 2694 3458 2698 3462
rect 2750 3458 2754 3462
rect 2822 3458 2826 3462
rect 2862 3458 2866 3462
rect 2950 3458 2954 3462
rect 2966 3458 2970 3462
rect 2990 3458 2994 3462
rect 2998 3458 3002 3462
rect 3078 3458 3082 3462
rect 3142 3458 3146 3462
rect 3198 3458 3202 3462
rect 3214 3458 3218 3462
rect 3230 3458 3234 3462
rect 3246 3458 3250 3462
rect 3254 3458 3258 3462
rect 3286 3458 3290 3462
rect 3318 3459 3322 3463
rect 3350 3458 3354 3462
rect 3430 3458 3434 3462
rect 3454 3458 3458 3462
rect 3566 3458 3570 3462
rect 3590 3458 3594 3462
rect 3630 3458 3634 3462
rect 3694 3458 3698 3462
rect 3710 3458 3714 3462
rect 3750 3458 3754 3462
rect 3822 3458 3826 3462
rect 3894 3459 3898 3463
rect 3926 3458 3930 3462
rect 3982 3458 3986 3462
rect 3998 3458 4002 3462
rect 4030 3458 4034 3462
rect 4070 3458 4074 3462
rect 4150 3458 4154 3462
rect 4230 3458 4234 3462
rect 4238 3458 4242 3462
rect 4278 3458 4282 3462
rect 4326 3458 4330 3462
rect 4382 3459 4386 3463
rect 4566 3459 4570 3463
rect 4614 3458 4618 3462
rect 4654 3458 4658 3462
rect 4702 3458 4706 3462
rect 4774 3458 4778 3462
rect 4846 3458 4850 3462
rect 4870 3458 4874 3462
rect 4910 3458 4914 3462
rect 4950 3458 4954 3462
rect 4990 3458 4994 3462
rect 5030 3458 5034 3462
rect 5038 3458 5042 3462
rect 5086 3458 5090 3462
rect 5142 3458 5146 3462
rect 5150 3458 5154 3462
rect 5174 3458 5178 3462
rect 5230 3458 5234 3462
rect 110 3448 114 3452
rect 270 3448 274 3452
rect 302 3448 306 3452
rect 470 3448 474 3452
rect 478 3448 482 3452
rect 542 3448 546 3452
rect 694 3448 698 3452
rect 942 3448 946 3452
rect 1230 3448 1234 3452
rect 1294 3448 1298 3452
rect 1534 3448 1538 3452
rect 1542 3448 1546 3452
rect 1566 3448 1570 3452
rect 1582 3448 1586 3452
rect 1750 3448 1754 3452
rect 1766 3448 1770 3452
rect 1798 3448 1802 3452
rect 2038 3448 2042 3452
rect 2142 3448 2146 3452
rect 2342 3448 2346 3452
rect 2366 3448 2370 3452
rect 2710 3448 2714 3452
rect 2846 3448 2850 3452
rect 2902 3448 2906 3452
rect 3150 3448 3154 3452
rect 3446 3448 3450 3452
rect 3526 3448 3530 3452
rect 3590 3448 3594 3452
rect 3798 3448 3802 3452
rect 4214 3448 4218 3452
rect 4494 3448 4498 3452
rect 4598 3448 4602 3452
rect 4678 3448 4682 3452
rect 4686 3448 4690 3452
rect 5014 3448 5018 3452
rect 246 3438 250 3442
rect 262 3438 266 3442
rect 1198 3438 1202 3442
rect 1518 3438 1522 3442
rect 1694 3438 1698 3442
rect 2190 3438 2194 3442
rect 2246 3438 2250 3442
rect 2806 3438 2810 3442
rect 3038 3438 3042 3442
rect 3766 3438 3770 3442
rect 4110 3438 4114 3442
rect 5062 3438 5066 3442
rect 3182 3428 3186 3432
rect 22 3418 26 3422
rect 118 3418 122 3422
rect 158 3418 162 3422
rect 454 3418 458 3422
rect 598 3418 602 3422
rect 1094 3418 1098 3422
rect 1502 3418 1506 3422
rect 1822 3418 1826 3422
rect 2694 3418 2698 3422
rect 2942 3418 2946 3422
rect 3126 3418 3130 3422
rect 3214 3418 3218 3422
rect 3430 3418 3434 3422
rect 3654 3418 3658 3422
rect 3854 3418 3858 3422
rect 3958 3418 3962 3422
rect 4022 3418 4026 3422
rect 4094 3418 4098 3422
rect 4310 3418 4314 3422
rect 4446 3418 4450 3422
rect 4502 3418 4506 3422
rect 4638 3418 4642 3422
rect 4702 3418 4706 3422
rect 4814 3418 4818 3422
rect 4942 3418 4946 3422
rect 5190 3418 5194 3422
rect 330 3403 334 3407
rect 337 3403 341 3407
rect 1354 3403 1358 3407
rect 1361 3403 1365 3407
rect 2386 3403 2390 3407
rect 2393 3403 2397 3407
rect 3402 3403 3406 3407
rect 3409 3403 3413 3407
rect 4426 3403 4430 3407
rect 4433 3403 4437 3407
rect 166 3388 170 3392
rect 942 3388 946 3392
rect 1550 3388 1554 3392
rect 1790 3388 1794 3392
rect 2086 3388 2090 3392
rect 3230 3388 3234 3392
rect 3294 3388 3298 3392
rect 3318 3388 3322 3392
rect 3710 3388 3714 3392
rect 3814 3388 3818 3392
rect 3886 3388 3890 3392
rect 3982 3388 3986 3392
rect 4126 3388 4130 3392
rect 4470 3388 4474 3392
rect 4566 3388 4570 3392
rect 4686 3388 4690 3392
rect 4766 3388 4770 3392
rect 5246 3388 5250 3392
rect 494 3378 498 3382
rect 734 3378 738 3382
rect 1518 3378 1522 3382
rect 318 3368 322 3372
rect 350 3368 354 3372
rect 1254 3368 1258 3372
rect 1294 3368 1298 3372
rect 1446 3368 1450 3372
rect 1462 3368 1466 3372
rect 1534 3368 1538 3372
rect 1606 3368 1610 3372
rect 1646 3368 1650 3372
rect 1774 3368 1778 3372
rect 1950 3368 1954 3372
rect 2118 3368 2122 3372
rect 2862 3368 2866 3372
rect 3006 3368 3010 3372
rect 3478 3368 3482 3372
rect 4406 3368 4410 3372
rect 4438 3368 4442 3372
rect 4518 3368 4522 3372
rect 4606 3368 4610 3372
rect 4902 3368 4906 3372
rect 78 3358 82 3362
rect 206 3358 210 3362
rect 94 3348 98 3352
rect 262 3348 266 3352
rect 334 3348 338 3352
rect 374 3358 378 3362
rect 558 3358 562 3362
rect 614 3358 618 3362
rect 750 3358 754 3362
rect 1006 3358 1010 3362
rect 1022 3358 1026 3362
rect 1126 3358 1130 3362
rect 1270 3358 1274 3362
rect 390 3348 394 3352
rect 438 3348 442 3352
rect 502 3348 506 3352
rect 550 3348 554 3352
rect 574 3348 578 3352
rect 598 3348 602 3352
rect 622 3348 626 3352
rect 638 3348 642 3352
rect 670 3347 674 3351
rect 742 3348 746 3352
rect 798 3348 802 3352
rect 862 3348 866 3352
rect 926 3348 930 3352
rect 958 3348 962 3352
rect 974 3348 978 3352
rect 990 3348 994 3352
rect 1006 3348 1010 3352
rect 1062 3348 1066 3352
rect 1198 3348 1202 3352
rect 1270 3348 1274 3352
rect 1494 3358 1498 3362
rect 1318 3348 1322 3352
rect 1406 3348 1410 3352
rect 1478 3348 1482 3352
rect 1502 3348 1506 3352
rect 1518 3348 1522 3352
rect 1550 3348 1554 3352
rect 1582 3348 1586 3352
rect 1590 3348 1594 3352
rect 1670 3358 1674 3362
rect 1806 3358 1810 3362
rect 2030 3358 2034 3362
rect 2070 3358 2074 3362
rect 2134 3358 2138 3362
rect 2142 3358 2146 3362
rect 2678 3358 2682 3362
rect 2734 3358 2738 3362
rect 3070 3358 3074 3362
rect 3270 3358 3274 3362
rect 3342 3358 3346 3362
rect 3358 3358 3362 3362
rect 3574 3358 3578 3362
rect 3590 3358 3594 3362
rect 3726 3358 3730 3362
rect 3782 3358 3786 3362
rect 3862 3358 3866 3362
rect 1670 3348 1674 3352
rect 6 3338 10 3342
rect 86 3338 90 3342
rect 102 3338 106 3342
rect 110 3338 114 3342
rect 182 3338 186 3342
rect 222 3338 226 3342
rect 254 3338 258 3342
rect 286 3338 290 3342
rect 342 3338 346 3342
rect 398 3338 402 3342
rect 414 3338 418 3342
rect 510 3338 514 3342
rect 582 3338 586 3342
rect 590 3338 594 3342
rect 678 3338 682 3342
rect 774 3338 778 3342
rect 886 3338 890 3342
rect 966 3338 970 3342
rect 998 3338 1002 3342
rect 1038 3338 1042 3342
rect 1142 3338 1146 3342
rect 1150 3338 1154 3342
rect 1174 3338 1178 3342
rect 1262 3338 1266 3342
rect 1318 3338 1322 3342
rect 1326 3338 1330 3342
rect 1334 3340 1338 3344
rect 1382 3338 1386 3342
rect 1470 3338 1474 3342
rect 1486 3338 1490 3342
rect 1526 3338 1530 3342
rect 1558 3338 1562 3342
rect 1710 3347 1714 3351
rect 1790 3348 1794 3352
rect 1814 3348 1818 3352
rect 1830 3348 1834 3352
rect 1894 3348 1898 3352
rect 1918 3348 1922 3352
rect 1958 3348 1962 3352
rect 1990 3348 1994 3352
rect 2014 3348 2018 3352
rect 2054 3348 2058 3352
rect 2078 3348 2082 3352
rect 2102 3348 2106 3352
rect 2126 3348 2130 3352
rect 2166 3348 2170 3352
rect 1622 3338 1626 3342
rect 1678 3338 1682 3342
rect 1694 3338 1698 3342
rect 1782 3338 1786 3342
rect 1822 3338 1826 3342
rect 1854 3338 1858 3342
rect 1966 3338 1970 3342
rect 2046 3338 2050 3342
rect 2262 3347 2266 3351
rect 2310 3348 2314 3352
rect 2342 3348 2346 3352
rect 2398 3348 2402 3352
rect 2422 3348 2426 3352
rect 2478 3348 2482 3352
rect 2486 3348 2490 3352
rect 2518 3348 2522 3352
rect 2558 3348 2562 3352
rect 2582 3348 2586 3352
rect 2622 3348 2626 3352
rect 2654 3348 2658 3352
rect 2694 3348 2698 3352
rect 2710 3348 2714 3352
rect 2718 3348 2722 3352
rect 2750 3348 2754 3352
rect 2766 3348 2770 3352
rect 2798 3347 2802 3351
rect 2886 3348 2890 3352
rect 2942 3347 2946 3351
rect 2974 3348 2978 3352
rect 3030 3348 3034 3352
rect 3046 3348 3050 3352
rect 3054 3348 3058 3352
rect 3078 3348 3082 3352
rect 3142 3348 3146 3352
rect 3166 3348 3170 3352
rect 3254 3348 3258 3352
rect 3278 3348 3282 3352
rect 3334 3348 3338 3352
rect 3358 3348 3362 3352
rect 3422 3348 3426 3352
rect 3446 3348 3450 3352
rect 3534 3348 3538 3352
rect 3542 3348 3546 3352
rect 3550 3348 3554 3352
rect 3590 3348 3594 3352
rect 3598 3348 3602 3352
rect 3622 3348 3626 3352
rect 3662 3348 3666 3352
rect 3678 3348 3682 3352
rect 3694 3348 3698 3352
rect 3710 3348 3714 3352
rect 3758 3348 3762 3352
rect 3766 3348 3770 3352
rect 3790 3348 3794 3352
rect 3798 3348 3802 3352
rect 3830 3348 3834 3352
rect 3846 3348 3850 3352
rect 3902 3358 3906 3362
rect 3950 3358 3954 3362
rect 4078 3358 4082 3362
rect 4094 3358 4098 3362
rect 4390 3358 4394 3362
rect 4486 3358 4490 3362
rect 3886 3348 3890 3352
rect 3902 3348 3906 3352
rect 3918 3348 3922 3352
rect 3966 3348 3970 3352
rect 4038 3348 4042 3352
rect 4102 3348 4106 3352
rect 4134 3348 4138 3352
rect 4142 3348 4146 3352
rect 4246 3348 4250 3352
rect 4358 3348 4362 3352
rect 4382 3348 4386 3352
rect 4406 3348 4410 3352
rect 4502 3348 4506 3352
rect 4534 3358 4538 3362
rect 4550 3358 4554 3362
rect 4550 3348 4554 3352
rect 4566 3348 4570 3352
rect 4590 3348 4594 3352
rect 4670 3358 4674 3362
rect 4630 3348 4634 3352
rect 4654 3348 4658 3352
rect 4686 3348 4690 3352
rect 4702 3348 4706 3352
rect 4718 3348 4722 3352
rect 4734 3348 4738 3352
rect 4750 3348 4754 3352
rect 4806 3348 4810 3352
rect 4830 3348 4834 3352
rect 4878 3348 4882 3352
rect 4934 3348 4938 3352
rect 5054 3348 5058 3352
rect 5094 3348 5098 3352
rect 5102 3348 5106 3352
rect 5118 3348 5122 3352
rect 5126 3348 5130 3352
rect 5198 3348 5202 3352
rect 2158 3338 2162 3342
rect 2246 3338 2250 3342
rect 2318 3338 2322 3342
rect 2334 3338 2338 3342
rect 2462 3338 2466 3342
rect 2630 3338 2634 3342
rect 2686 3338 2690 3342
rect 2702 3338 2706 3342
rect 2782 3338 2786 3342
rect 2894 3338 2898 3342
rect 3038 3338 3042 3342
rect 3086 3338 3090 3342
rect 3206 3338 3210 3342
rect 3246 3338 3250 3342
rect 3374 3338 3378 3342
rect 3598 3338 3602 3342
rect 3750 3338 3754 3342
rect 3838 3338 3842 3342
rect 3894 3338 3898 3342
rect 3942 3338 3946 3342
rect 3974 3338 3978 3342
rect 4014 3338 4018 3342
rect 4062 3338 4066 3342
rect 4094 3338 4098 3342
rect 4110 3338 4114 3342
rect 4174 3338 4178 3342
rect 4278 3338 4282 3342
rect 4294 3338 4298 3342
rect 4358 3338 4362 3342
rect 4366 3338 4370 3342
rect 4398 3338 4402 3342
rect 4478 3338 4482 3342
rect 4494 3338 4498 3342
rect 4542 3338 4546 3342
rect 4574 3338 4578 3342
rect 4582 3338 4586 3342
rect 4638 3338 4642 3342
rect 4646 3338 4650 3342
rect 4718 3338 4722 3342
rect 4806 3338 4810 3342
rect 4870 3338 4874 3342
rect 4966 3338 4970 3342
rect 5062 3338 5066 3342
rect 5222 3338 5226 3342
rect 5238 3338 5242 3342
rect 5302 3338 5306 3342
rect 534 3328 538 3332
rect 550 3328 554 3332
rect 622 3328 626 3332
rect 702 3328 706 3332
rect 758 3328 762 3332
rect 894 3328 898 3332
rect 910 3328 914 3332
rect 990 3328 994 3332
rect 1150 3328 1154 3332
rect 1566 3328 1570 3332
rect 1582 3328 1586 3332
rect 1838 3328 1842 3332
rect 2006 3328 2010 3332
rect 2294 3328 2298 3332
rect 2390 3328 2394 3332
rect 2494 3328 2498 3332
rect 2638 3328 2642 3332
rect 2670 3328 2674 3332
rect 2766 3328 2770 3332
rect 3566 3328 3570 3332
rect 3622 3328 3626 3332
rect 3662 3328 3666 3332
rect 3950 3328 3954 3332
rect 4126 3328 4130 3332
rect 4190 3328 4194 3332
rect 4718 3328 4722 3332
rect 4734 3328 4738 3332
rect 4806 3328 4810 3332
rect 4822 3328 4826 3332
rect 4846 3328 4850 3332
rect 62 3318 66 3322
rect 198 3318 202 3322
rect 214 3318 218 3322
rect 518 3318 522 3322
rect 630 3318 634 3322
rect 854 3318 858 3322
rect 1118 3318 1122 3322
rect 1126 3318 1130 3322
rect 1366 3318 1370 3322
rect 1974 3318 1978 3322
rect 2118 3318 2122 3322
rect 2142 3318 2146 3322
rect 2182 3318 2186 3322
rect 2198 3318 2202 3322
rect 2614 3318 2618 3322
rect 2870 3318 2874 3322
rect 3014 3318 3018 3322
rect 3270 3318 3274 3322
rect 3294 3318 3298 3322
rect 3318 3318 3322 3322
rect 3518 3318 3522 3322
rect 3558 3318 3562 3322
rect 3638 3318 3642 3322
rect 3782 3318 3786 3322
rect 4614 3318 4618 3322
rect 4862 3318 4866 3322
rect 4886 3318 4890 3322
rect 4998 3318 5002 3322
rect 5142 3318 5146 3322
rect 850 3303 854 3307
rect 857 3303 861 3307
rect 1874 3303 1878 3307
rect 1881 3303 1885 3307
rect 2890 3303 2894 3307
rect 2897 3303 2901 3307
rect 3922 3303 3926 3307
rect 3929 3303 3933 3307
rect 4938 3303 4942 3307
rect 4945 3303 4949 3307
rect 6 3288 10 3292
rect 110 3288 114 3292
rect 438 3288 442 3292
rect 454 3288 458 3292
rect 598 3288 602 3292
rect 654 3288 658 3292
rect 1486 3288 1490 3292
rect 2134 3288 2138 3292
rect 2230 3288 2234 3292
rect 2286 3288 2290 3292
rect 2462 3288 2466 3292
rect 2510 3288 2514 3292
rect 2582 3288 2586 3292
rect 2654 3288 2658 3292
rect 2710 3288 2714 3292
rect 2942 3288 2946 3292
rect 3086 3288 3090 3292
rect 3102 3288 3106 3292
rect 3286 3288 3290 3292
rect 3566 3288 3570 3292
rect 3830 3288 3834 3292
rect 4174 3288 4178 3292
rect 4270 3288 4274 3292
rect 4366 3288 4370 3292
rect 4486 3288 4490 3292
rect 4534 3288 4538 3292
rect 4790 3288 4794 3292
rect 5206 3288 5210 3292
rect 70 3278 74 3282
rect 102 3278 106 3282
rect 446 3278 450 3282
rect 558 3278 562 3282
rect 774 3278 778 3282
rect 854 3278 858 3282
rect 982 3278 986 3282
rect 1206 3278 1210 3282
rect 1382 3278 1386 3282
rect 1638 3278 1642 3282
rect 2030 3278 2034 3282
rect 2390 3278 2394 3282
rect 2494 3278 2498 3282
rect 2646 3278 2650 3282
rect 2694 3278 2698 3282
rect 2726 3278 2730 3282
rect 3222 3278 3226 3282
rect 3350 3278 3354 3282
rect 3398 3278 3402 3282
rect 3438 3278 3442 3282
rect 3470 3278 3474 3282
rect 3758 3278 3762 3282
rect 3990 3278 3994 3282
rect 4198 3278 4202 3282
rect 4622 3278 4626 3282
rect 4830 3278 4834 3282
rect 4942 3278 4946 3282
rect 4982 3278 4986 3282
rect 5102 3278 5106 3282
rect 5182 3278 5186 3282
rect 5270 3278 5274 3282
rect 118 3268 122 3272
rect 286 3268 290 3272
rect 406 3268 410 3272
rect 646 3268 650 3272
rect 678 3268 682 3272
rect 686 3268 690 3272
rect 742 3268 746 3272
rect 1150 3268 1154 3272
rect 1334 3268 1338 3272
rect 1478 3268 1482 3272
rect 1510 3268 1514 3272
rect 1542 3268 1546 3272
rect 1550 3268 1554 3272
rect 1582 3268 1586 3272
rect 1590 3268 1594 3272
rect 1710 3268 1714 3272
rect 1726 3268 1730 3272
rect 1774 3268 1778 3272
rect 1830 3268 1834 3272
rect 1870 3268 1874 3272
rect 1894 3268 1898 3272
rect 1910 3268 1914 3272
rect 1934 3268 1938 3272
rect 2038 3268 2042 3272
rect 2094 3268 2098 3272
rect 2102 3268 2106 3272
rect 2214 3268 2218 3272
rect 2254 3268 2258 3272
rect 2262 3268 2266 3272
rect 2294 3268 2298 3272
rect 2334 3268 2338 3272
rect 2406 3268 2410 3272
rect 2438 3268 2442 3272
rect 2470 3268 2474 3272
rect 2566 3268 2570 3272
rect 2638 3268 2642 3272
rect 2662 3268 2666 3272
rect 2694 3268 2698 3272
rect 2742 3268 2746 3272
rect 2806 3268 2810 3272
rect 2838 3268 2842 3272
rect 2870 3268 2874 3272
rect 2966 3268 2970 3272
rect 2990 3268 2994 3272
rect 3062 3268 3066 3272
rect 3126 3268 3130 3272
rect 3142 3268 3146 3272
rect 3238 3268 3242 3272
rect 3454 3268 3458 3272
rect 3470 3268 3474 3272
rect 3486 3268 3490 3272
rect 3582 3268 3586 3272
rect 3670 3268 3674 3272
rect 3686 3268 3690 3272
rect 3726 3268 3730 3272
rect 3742 3268 3746 3272
rect 3878 3268 3882 3272
rect 4022 3268 4026 3272
rect 4046 3268 4050 3272
rect 4078 3268 4082 3272
rect 4118 3268 4122 3272
rect 4222 3268 4226 3272
rect 4294 3268 4298 3272
rect 4302 3268 4306 3272
rect 4326 3268 4330 3272
rect 4358 3268 4362 3272
rect 4446 3268 4450 3272
rect 4478 3268 4482 3272
rect 4510 3268 4514 3272
rect 4518 3268 4522 3272
rect 4542 3268 4546 3272
rect 4598 3268 4602 3272
rect 4798 3268 4802 3272
rect 4878 3268 4882 3272
rect 4886 3268 4890 3272
rect 4902 3268 4906 3272
rect 4918 3268 4922 3272
rect 4950 3268 4954 3272
rect 5062 3268 5066 3272
rect 5126 3268 5130 3272
rect 5142 3268 5146 3272
rect 70 3259 74 3263
rect 198 3258 202 3262
rect 206 3258 210 3262
rect 294 3258 298 3262
rect 382 3258 386 3262
rect 470 3258 474 3262
rect 558 3259 562 3263
rect 614 3258 618 3262
rect 638 3258 642 3262
rect 670 3258 674 3262
rect 694 3258 698 3262
rect 734 3258 738 3262
rect 774 3259 778 3263
rect 886 3258 890 3262
rect 910 3258 914 3262
rect 918 3258 922 3262
rect 950 3258 954 3262
rect 990 3258 994 3262
rect 1078 3258 1082 3262
rect 1094 3258 1098 3262
rect 1102 3258 1106 3262
rect 1134 3258 1138 3262
rect 1142 3258 1146 3262
rect 1158 3258 1162 3262
rect 1166 3258 1170 3262
rect 1206 3259 1210 3263
rect 1278 3258 1282 3262
rect 1302 3258 1306 3262
rect 1326 3258 1330 3262
rect 1390 3258 1394 3262
rect 1478 3258 1482 3262
rect 1502 3258 1506 3262
rect 1534 3258 1538 3262
rect 1558 3258 1562 3262
rect 1582 3258 1586 3262
rect 1606 3258 1610 3262
rect 1646 3258 1650 3262
rect 1734 3258 1738 3262
rect 1758 3258 1762 3262
rect 1766 3258 1770 3262
rect 1782 3258 1786 3262
rect 1806 3258 1810 3262
rect 1822 3258 1826 3262
rect 1846 3258 1850 3262
rect 1902 3258 1906 3262
rect 1958 3258 1962 3262
rect 2046 3258 2050 3262
rect 2110 3258 2114 3262
rect 2198 3259 2202 3263
rect 2246 3258 2250 3262
rect 2270 3258 2274 3262
rect 2302 3258 2306 3262
rect 2382 3258 2386 3262
rect 2446 3258 2450 3262
rect 2478 3258 2482 3262
rect 2662 3258 2666 3262
rect 2670 3258 2674 3262
rect 2750 3258 2754 3262
rect 2758 3258 2762 3262
rect 2766 3258 2770 3262
rect 2790 3258 2794 3262
rect 2814 3258 2818 3262
rect 2830 3258 2834 3262
rect 2846 3258 2850 3262
rect 2870 3258 2874 3262
rect 2894 3258 2898 3262
rect 2902 3258 2906 3262
rect 2926 3258 2930 3262
rect 2958 3258 2962 3262
rect 3070 3258 3074 3262
rect 3118 3258 3122 3262
rect 3166 3258 3170 3262
rect 3230 3258 3234 3262
rect 3262 3258 3266 3262
rect 3326 3258 3330 3262
rect 3382 3258 3386 3262
rect 3414 3258 3418 3262
rect 3446 3258 3450 3262
rect 3502 3259 3506 3263
rect 3534 3258 3538 3262
rect 3614 3258 3618 3262
rect 3630 3258 3634 3262
rect 3678 3258 3682 3262
rect 3718 3258 3722 3262
rect 3734 3258 3738 3262
rect 3774 3258 3778 3262
rect 3798 3258 3802 3262
rect 3806 3258 3810 3262
rect 3814 3258 3818 3262
rect 3846 3258 3850 3262
rect 3886 3258 3890 3262
rect 3918 3258 3922 3262
rect 3990 3259 3994 3263
rect 4038 3258 4042 3262
rect 4062 3258 4066 3262
rect 4070 3258 4074 3262
rect 4126 3258 4130 3262
rect 4182 3258 4186 3262
rect 4198 3258 4202 3262
rect 4254 3258 4258 3262
rect 4262 3258 4266 3262
rect 4286 3258 4290 3262
rect 4310 3258 4314 3262
rect 4334 3258 4338 3262
rect 4342 3258 4346 3262
rect 4350 3258 4354 3262
rect 4422 3258 4426 3262
rect 4486 3258 4490 3262
rect 4502 3258 4506 3262
rect 4550 3258 4554 3262
rect 4590 3258 4594 3262
rect 4638 3258 4642 3262
rect 4662 3258 4666 3262
rect 4726 3259 4730 3263
rect 4846 3258 4850 3262
rect 4870 3258 4874 3262
rect 4878 3258 4882 3262
rect 4910 3258 4914 3262
rect 4926 3258 4930 3262
rect 4942 3258 4946 3262
rect 4966 3258 4970 3262
rect 5062 3258 5066 3262
rect 5118 3258 5122 3262
rect 5150 3258 5154 3262
rect 5158 3258 5162 3262
rect 5198 3258 5202 3262
rect 5270 3259 5274 3263
rect 190 3248 194 3252
rect 622 3248 626 3252
rect 638 3248 642 3252
rect 654 3248 658 3252
rect 710 3248 714 3252
rect 1094 3248 1098 3252
rect 1174 3248 1178 3252
rect 1294 3248 1298 3252
rect 1310 3248 1314 3252
rect 1454 3248 1458 3252
rect 1486 3248 1490 3252
rect 1518 3248 1522 3252
rect 1574 3248 1578 3252
rect 1606 3248 1610 3252
rect 1806 3248 1810 3252
rect 1918 3248 1922 3252
rect 2230 3248 2234 3252
rect 2286 3248 2290 3252
rect 2302 3248 2306 3252
rect 2462 3248 2466 3252
rect 2494 3248 2498 3252
rect 2702 3248 2706 3252
rect 2718 3248 2722 3252
rect 2830 3248 2834 3252
rect 2942 3248 2946 3252
rect 2974 3248 2978 3252
rect 2990 3248 2994 3252
rect 3102 3248 3106 3252
rect 3254 3248 3258 3252
rect 3902 3248 3906 3252
rect 4022 3248 4026 3252
rect 4054 3248 4058 3252
rect 4270 3248 4274 3252
rect 4334 3248 4338 3252
rect 4534 3248 4538 3252
rect 4590 3248 4594 3252
rect 4814 3248 4818 3252
rect 4854 3248 4858 3252
rect 4870 3248 4874 3252
rect 734 3238 738 3242
rect 838 3238 842 3242
rect 1470 3238 1474 3242
rect 1534 3238 1538 3242
rect 2046 3238 2050 3242
rect 2070 3238 2074 3242
rect 3662 3238 3666 3242
rect 3702 3238 3706 3242
rect 4566 3238 4570 3242
rect 4606 3238 4610 3242
rect 5158 3238 5162 3242
rect 1822 3228 1826 3232
rect 2110 3228 2114 3232
rect 110 3218 114 3222
rect 174 3218 178 3222
rect 222 3218 226 3222
rect 494 3218 498 3222
rect 870 3218 874 3222
rect 902 3218 906 3222
rect 934 3218 938 3222
rect 1062 3218 1066 3222
rect 1126 3218 1130 3222
rect 1270 3218 1274 3222
rect 1862 3218 1866 3222
rect 2014 3218 2018 3222
rect 2022 3218 2026 3222
rect 2726 3218 2730 3222
rect 2782 3218 2786 3222
rect 2862 3218 2866 3222
rect 2918 3218 2922 3222
rect 3006 3218 3010 3222
rect 3222 3218 3226 3222
rect 3390 3218 3394 3222
rect 3430 3218 3434 3222
rect 3758 3218 3762 3222
rect 3790 3218 3794 3222
rect 3862 3218 3866 3222
rect 4806 3218 4810 3222
rect 4830 3218 4834 3222
rect 4990 3218 4994 3222
rect 5190 3218 5194 3222
rect 330 3203 334 3207
rect 337 3203 341 3207
rect 1354 3203 1358 3207
rect 1361 3203 1365 3207
rect 2386 3203 2390 3207
rect 2393 3203 2397 3207
rect 3402 3203 3406 3207
rect 3409 3203 3413 3207
rect 4426 3203 4430 3207
rect 4433 3203 4437 3207
rect 278 3188 282 3192
rect 1134 3188 1138 3192
rect 1158 3188 1162 3192
rect 1182 3188 1186 3192
rect 1670 3188 1674 3192
rect 1694 3188 1698 3192
rect 2014 3188 2018 3192
rect 2030 3188 2034 3192
rect 2470 3188 2474 3192
rect 2606 3188 2610 3192
rect 2870 3188 2874 3192
rect 3742 3188 3746 3192
rect 4126 3188 4130 3192
rect 4318 3188 4322 3192
rect 4686 3188 4690 3192
rect 4710 3188 4714 3192
rect 4782 3188 4786 3192
rect 5030 3188 5034 3192
rect 5102 3188 5106 3192
rect 1350 3178 1354 3182
rect 1934 3178 1938 3182
rect 4590 3178 4594 3182
rect 5166 3178 5170 3182
rect 558 3168 562 3172
rect 622 3168 626 3172
rect 1222 3168 1226 3172
rect 1382 3168 1386 3172
rect 2790 3168 2794 3172
rect 3014 3168 3018 3172
rect 3126 3168 3130 3172
rect 4534 3168 4538 3172
rect 4550 3168 4554 3172
rect 4894 3168 4898 3172
rect 102 3147 106 3151
rect 198 3147 202 3151
rect 294 3148 298 3152
rect 342 3147 346 3151
rect 414 3148 418 3152
rect 446 3148 450 3152
rect 502 3148 506 3152
rect 582 3148 586 3152
rect 598 3148 602 3152
rect 702 3158 706 3162
rect 750 3158 754 3162
rect 766 3158 770 3162
rect 782 3158 786 3162
rect 886 3158 890 3162
rect 918 3158 922 3162
rect 1150 3158 1154 3162
rect 1190 3158 1194 3162
rect 638 3148 642 3152
rect 678 3148 682 3152
rect 686 3148 690 3152
rect 718 3148 722 3152
rect 774 3148 778 3152
rect 782 3148 786 3152
rect 798 3148 802 3152
rect 838 3148 842 3152
rect 870 3148 874 3152
rect 878 3148 882 3152
rect 902 3148 906 3152
rect 918 3148 922 3152
rect 950 3147 954 3151
rect 1022 3148 1026 3152
rect 1054 3148 1058 3152
rect 1078 3148 1082 3152
rect 1206 3148 1210 3152
rect 1398 3158 1402 3162
rect 1414 3158 1418 3162
rect 1430 3158 1434 3162
rect 1494 3158 1498 3162
rect 1590 3158 1594 3162
rect 1238 3148 1242 3152
rect 1246 3148 1250 3152
rect 1286 3147 1290 3151
rect 1374 3148 1378 3152
rect 1414 3148 1418 3152
rect 1438 3148 1442 3152
rect 1454 3148 1458 3152
rect 1478 3148 1482 3152
rect 1502 3148 1506 3152
rect 1558 3148 1562 3152
rect 1574 3148 1578 3152
rect 1654 3158 1658 3162
rect 1686 3158 1690 3162
rect 2078 3158 2082 3162
rect 2342 3158 2346 3162
rect 2358 3158 2362 3162
rect 2478 3158 2482 3162
rect 2510 3158 2514 3162
rect 2542 3158 2546 3162
rect 2622 3158 2626 3162
rect 2654 3158 2658 3162
rect 2670 3158 2674 3162
rect 2686 3158 2690 3162
rect 2822 3158 2826 3162
rect 2838 3158 2842 3162
rect 2878 3158 2882 3162
rect 3238 3158 3242 3162
rect 3358 3158 3362 3162
rect 3446 3158 3450 3162
rect 3686 3158 3690 3162
rect 3854 3158 3858 3162
rect 3966 3158 3970 3162
rect 4110 3158 4114 3162
rect 4350 3158 4354 3162
rect 4358 3158 4362 3162
rect 4430 3158 4434 3162
rect 4494 3158 4498 3162
rect 4558 3158 4562 3162
rect 4734 3158 4738 3162
rect 4822 3158 4826 3162
rect 4854 3158 4858 3162
rect 1622 3148 1626 3152
rect 1638 3148 1642 3152
rect 1670 3148 1674 3152
rect 1750 3148 1754 3152
rect 1806 3148 1810 3152
rect 1846 3148 1850 3152
rect 1974 3148 1978 3152
rect 1982 3148 1986 3152
rect 1990 3148 1994 3152
rect 2046 3148 2050 3152
rect 2062 3148 2066 3152
rect 2086 3148 2090 3152
rect 2102 3148 2106 3152
rect 2142 3148 2146 3152
rect 2166 3148 2170 3152
rect 2230 3148 2234 3152
rect 2254 3148 2258 3152
rect 2262 3148 2266 3152
rect 2270 3148 2274 3152
rect 2302 3148 2306 3152
rect 2334 3148 2338 3152
rect 2422 3148 2426 3152
rect 2478 3148 2482 3152
rect 2494 3148 2498 3152
rect 2518 3148 2522 3152
rect 2534 3148 2538 3152
rect 2574 3148 2578 3152
rect 2638 3148 2642 3152
rect 2654 3148 2658 3152
rect 2726 3148 2730 3152
rect 2798 3148 2802 3152
rect 2846 3148 2850 3152
rect 2894 3148 2898 3152
rect 2926 3148 2930 3152
rect 2974 3148 2978 3152
rect 2990 3148 2994 3152
rect 3006 3148 3010 3152
rect 3046 3148 3050 3152
rect 3054 3148 3058 3152
rect 3142 3148 3146 3152
rect 3166 3148 3170 3152
rect 3174 3148 3178 3152
rect 3198 3148 3202 3152
rect 3206 3148 3210 3152
rect 3222 3148 3226 3152
rect 3254 3148 3258 3152
rect 6 3138 10 3142
rect 70 3138 74 3142
rect 86 3138 90 3142
rect 182 3138 186 3142
rect 230 3138 234 3142
rect 326 3138 330 3142
rect 374 3138 378 3142
rect 422 3138 426 3142
rect 478 3138 482 3142
rect 590 3138 594 3142
rect 606 3138 610 3142
rect 646 3138 650 3142
rect 742 3138 746 3142
rect 774 3138 778 3142
rect 814 3138 818 3142
rect 822 3138 826 3142
rect 846 3138 850 3142
rect 894 3138 898 3142
rect 958 3138 962 3142
rect 1030 3138 1034 3142
rect 1078 3138 1082 3142
rect 1150 3138 1154 3142
rect 1174 3138 1178 3142
rect 1198 3138 1202 3142
rect 1254 3138 1258 3142
rect 1270 3138 1274 3142
rect 1374 3138 1378 3142
rect 1406 3138 1410 3142
rect 1446 3138 1450 3142
rect 1470 3138 1474 3142
rect 1550 3138 1554 3142
rect 1566 3138 1570 3142
rect 1606 3138 1610 3142
rect 1622 3138 1626 3142
rect 1630 3138 1634 3142
rect 1662 3138 1666 3142
rect 1774 3138 1778 3142
rect 1854 3138 1858 3142
rect 1942 3138 1946 3142
rect 1998 3138 2002 3142
rect 2054 3138 2058 3142
rect 3286 3147 3290 3151
rect 3374 3148 3378 3152
rect 3446 3148 3450 3152
rect 3470 3148 3474 3152
rect 3502 3148 3506 3152
rect 3510 3148 3514 3152
rect 3558 3148 3562 3152
rect 3590 3147 3594 3151
rect 3710 3148 3714 3152
rect 3734 3148 3738 3152
rect 3814 3148 3818 3152
rect 3854 3148 3858 3152
rect 3902 3148 3906 3152
rect 3910 3148 3914 3152
rect 4014 3147 4018 3151
rect 4094 3148 4098 3152
rect 4102 3148 4106 3152
rect 4126 3148 4130 3152
rect 4142 3148 4146 3152
rect 4150 3148 4154 3152
rect 4174 3148 4178 3152
rect 4262 3148 4266 3152
rect 4302 3148 4306 3152
rect 4374 3148 4378 3152
rect 4414 3148 4418 3152
rect 4438 3148 4442 3152
rect 4462 3148 4466 3152
rect 4510 3148 4514 3152
rect 4534 3148 4538 3152
rect 4574 3148 4578 3152
rect 4646 3148 4650 3152
rect 4726 3148 4730 3152
rect 4750 3148 4754 3152
rect 4766 3148 4770 3152
rect 4806 3148 4810 3152
rect 4838 3148 4842 3152
rect 5054 3158 5058 3162
rect 5086 3158 5090 3162
rect 5142 3158 5146 3162
rect 4870 3148 4874 3152
rect 4878 3148 4882 3152
rect 4942 3148 4946 3152
rect 5006 3148 5010 3152
rect 5014 3148 5018 3152
rect 5038 3148 5042 3152
rect 5086 3148 5090 3152
rect 5102 3148 5106 3152
rect 5118 3148 5122 3152
rect 5126 3148 5130 3152
rect 5174 3148 5178 3152
rect 5238 3147 5242 3151
rect 2222 3138 2226 3142
rect 2278 3138 2282 3142
rect 2310 3138 2314 3142
rect 2334 3138 2338 3142
rect 2390 3138 2394 3142
rect 2406 3138 2410 3142
rect 2502 3138 2506 3142
rect 2534 3138 2538 3142
rect 2558 3138 2562 3142
rect 2566 3138 2570 3142
rect 2598 3138 2602 3142
rect 2630 3138 2634 3142
rect 2662 3138 2666 3142
rect 2790 3138 2794 3142
rect 2838 3138 2842 3142
rect 2854 3138 2858 3142
rect 2902 3138 2906 3142
rect 2918 3138 2922 3142
rect 2998 3138 3002 3142
rect 3110 3138 3114 3142
rect 3134 3138 3138 3142
rect 3422 3138 3426 3142
rect 3478 3138 3482 3142
rect 3526 3138 3530 3142
rect 3534 3138 3538 3142
rect 3550 3138 3554 3142
rect 3558 3138 3562 3142
rect 3662 3138 3666 3142
rect 3838 3138 3842 3142
rect 3886 3138 3890 3142
rect 3902 3138 3906 3142
rect 4030 3138 4034 3142
rect 4070 3138 4074 3142
rect 4134 3138 4138 3142
rect 4182 3138 4186 3142
rect 4286 3138 4290 3142
rect 4334 3138 4338 3142
rect 4366 3138 4370 3142
rect 4382 3138 4386 3142
rect 4406 3138 4410 3142
rect 4470 3138 4474 3142
rect 4518 3138 4522 3142
rect 4526 3138 4530 3142
rect 4566 3138 4570 3142
rect 4582 3138 4586 3142
rect 4670 3138 4674 3142
rect 4758 3138 4762 3142
rect 4798 3138 4802 3142
rect 4830 3138 4834 3142
rect 4886 3138 4890 3142
rect 4974 3138 4978 3142
rect 5078 3138 5082 3142
rect 5110 3138 5114 3142
rect 5190 3138 5194 3142
rect 430 3128 434 3132
rect 462 3128 466 3132
rect 566 3128 570 3132
rect 1070 3128 1074 3132
rect 1094 3128 1098 3132
rect 1102 3128 1106 3132
rect 1462 3128 1466 3132
rect 1494 3128 1498 3132
rect 1534 3128 1538 3132
rect 1654 3128 1658 3132
rect 1790 3128 1794 3132
rect 1806 3128 1810 3132
rect 2014 3128 2018 3132
rect 2086 3128 2090 3132
rect 2294 3128 2298 3132
rect 2326 3128 2330 3132
rect 2654 3128 2658 3132
rect 2718 3128 2722 3132
rect 2950 3128 2954 3132
rect 2958 3128 2962 3132
rect 3286 3128 3290 3132
rect 3398 3128 3402 3132
rect 3454 3128 3458 3132
rect 3534 3128 3538 3132
rect 3718 3128 3722 3132
rect 3886 3128 3890 3132
rect 4046 3128 4050 3132
rect 4390 3128 4394 3132
rect 4422 3128 4426 3132
rect 4694 3128 4698 3132
rect 5174 3128 5178 3132
rect 5206 3128 5210 3132
rect 5238 3128 5242 3132
rect 166 3118 170 3122
rect 262 3118 266 3122
rect 278 3118 282 3122
rect 406 3118 410 3122
rect 574 3118 578 3122
rect 662 3118 666 3122
rect 1014 3118 1018 3122
rect 1038 3118 1042 3122
rect 1518 3118 1522 3122
rect 1542 3118 1546 3122
rect 1798 3118 1802 3122
rect 2030 3118 2034 3122
rect 2094 3118 2098 3122
rect 2286 3118 2290 3122
rect 2318 3118 2322 3122
rect 2542 3118 2546 3122
rect 2814 3118 2818 3122
rect 2942 3118 2946 3122
rect 3118 3118 3122 3122
rect 3158 3118 3162 3122
rect 3182 3118 3186 3122
rect 3446 3118 3450 3122
rect 3518 3118 3522 3122
rect 3654 3118 3658 3122
rect 4342 3118 4346 3122
rect 4398 3118 4402 3122
rect 4478 3118 4482 3122
rect 4734 3118 4738 3122
rect 4822 3118 4826 3122
rect 5054 3118 5058 3122
rect 5198 3118 5202 3122
rect 5302 3118 5306 3122
rect 850 3103 854 3107
rect 857 3103 861 3107
rect 1874 3103 1878 3107
rect 1881 3103 1885 3107
rect 2890 3103 2894 3107
rect 2897 3103 2901 3107
rect 3922 3103 3926 3107
rect 3929 3103 3933 3107
rect 4938 3103 4942 3107
rect 4945 3103 4949 3107
rect 94 3088 98 3092
rect 182 3088 186 3092
rect 310 3088 314 3092
rect 454 3088 458 3092
rect 590 3088 594 3092
rect 758 3088 762 3092
rect 1022 3088 1026 3092
rect 1374 3088 1378 3092
rect 1646 3088 1650 3092
rect 1710 3088 1714 3092
rect 1822 3088 1826 3092
rect 1934 3088 1938 3092
rect 2310 3088 2314 3092
rect 2486 3088 2490 3092
rect 2526 3088 2530 3092
rect 2566 3088 2570 3092
rect 2782 3088 2786 3092
rect 3206 3088 3210 3092
rect 3630 3088 3634 3092
rect 3662 3088 3666 3092
rect 3990 3088 3994 3092
rect 4038 3088 4042 3092
rect 4238 3088 4242 3092
rect 4918 3088 4922 3092
rect 4990 3088 4994 3092
rect 126 3078 130 3082
rect 214 3078 218 3082
rect 358 3078 362 3082
rect 390 3078 394 3082
rect 486 3078 490 3082
rect 574 3078 578 3082
rect 6 3068 10 3072
rect 86 3068 90 3072
rect 174 3068 178 3072
rect 222 3068 226 3072
rect 302 3068 306 3072
rect 630 3078 634 3082
rect 598 3068 602 3072
rect 814 3078 818 3082
rect 958 3078 962 3082
rect 1278 3078 1282 3082
rect 1286 3078 1290 3082
rect 1438 3078 1442 3082
rect 1478 3078 1482 3082
rect 1542 3078 1546 3082
rect 1654 3078 1658 3082
rect 1718 3078 1722 3082
rect 1926 3078 1930 3082
rect 2030 3078 2034 3082
rect 654 3068 658 3072
rect 678 3068 682 3072
rect 774 3068 778 3072
rect 798 3068 802 3072
rect 846 3068 850 3072
rect 942 3068 946 3072
rect 1038 3068 1042 3072
rect 1150 3068 1154 3072
rect 1198 3068 1202 3072
rect 1326 3068 1330 3072
rect 1334 3068 1338 3072
rect 1382 3068 1386 3072
rect 1414 3068 1418 3072
rect 1470 3068 1474 3072
rect 1598 3068 1602 3072
rect 1638 3068 1642 3072
rect 1654 3068 1658 3072
rect 1702 3068 1706 3072
rect 1846 3068 1850 3072
rect 1854 3068 1858 3072
rect 1894 3068 1898 3072
rect 2054 3068 2058 3072
rect 2070 3068 2074 3072
rect 2142 3068 2146 3072
rect 2294 3068 2298 3072
rect 2342 3068 2346 3072
rect 2390 3068 2394 3072
rect 2430 3068 2434 3072
rect 2454 3078 2458 3082
rect 2478 3078 2482 3082
rect 3198 3078 3202 3082
rect 3302 3078 3306 3082
rect 3438 3078 3442 3082
rect 3574 3078 3578 3082
rect 3670 3078 3674 3082
rect 3758 3078 3762 3082
rect 3766 3078 3770 3082
rect 3902 3078 3906 3082
rect 3934 3078 3938 3082
rect 3982 3078 3986 3082
rect 4134 3078 4138 3082
rect 4350 3078 4354 3082
rect 4638 3078 4642 3082
rect 4654 3078 4658 3082
rect 4694 3078 4698 3082
rect 5126 3078 5130 3082
rect 2494 3068 2498 3072
rect 2558 3068 2562 3072
rect 2590 3068 2594 3072
rect 2638 3068 2642 3072
rect 2718 3068 2722 3072
rect 2726 3068 2730 3072
rect 2758 3068 2762 3072
rect 2838 3068 2842 3072
rect 2982 3068 2986 3072
rect 3022 3068 3026 3072
rect 3134 3068 3138 3072
rect 3174 3068 3178 3072
rect 3182 3068 3186 3072
rect 3286 3068 3290 3072
rect 3326 3068 3330 3072
rect 3390 3068 3394 3072
rect 3422 3068 3426 3072
rect 78 3058 82 3062
rect 110 3058 114 3062
rect 158 3058 162 3062
rect 166 3058 170 3062
rect 198 3058 202 3062
rect 286 3058 290 3062
rect 294 3058 298 3062
rect 326 3058 330 3062
rect 398 3058 402 3062
rect 494 3058 498 3062
rect 558 3058 562 3062
rect 606 3058 610 3062
rect 614 3058 618 3062
rect 646 3058 650 3062
rect 662 3058 666 3062
rect 694 3059 698 3063
rect 766 3058 770 3062
rect 798 3058 802 3062
rect 862 3059 866 3063
rect 966 3058 970 3062
rect 1062 3058 1066 3062
rect 1126 3058 1130 3062
rect 1142 3058 1146 3062
rect 1174 3058 1178 3062
rect 1182 3058 1186 3062
rect 1222 3058 1226 3062
rect 1302 3058 1306 3062
rect 1310 3058 1314 3062
rect 1342 3058 1346 3062
rect 1390 3058 1394 3062
rect 1406 3058 1410 3062
rect 1422 3058 1426 3062
rect 1446 3058 1450 3062
rect 1462 3058 1466 3062
rect 1502 3058 1506 3062
rect 1526 3058 1530 3062
rect 1534 3058 1538 3062
rect 1558 3058 1562 3062
rect 1574 3058 1578 3062
rect 1606 3058 1610 3062
rect 1630 3058 1634 3062
rect 1670 3058 1674 3062
rect 1678 3058 1682 3062
rect 1694 3058 1698 3062
rect 1766 3058 1770 3062
rect 1782 3058 1786 3062
rect 1838 3058 1842 3062
rect 1862 3058 1866 3062
rect 1894 3058 1898 3062
rect 1902 3058 1906 3062
rect 1918 3058 1922 3062
rect 1966 3058 1970 3062
rect 1998 3059 2002 3063
rect 2046 3058 2050 3062
rect 2078 3058 2082 3062
rect 2094 3058 2098 3062
rect 2118 3058 2122 3062
rect 2126 3058 2130 3062
rect 2134 3058 2138 3062
rect 2182 3058 2186 3062
rect 2278 3059 2282 3063
rect 2374 3059 2378 3063
rect 2414 3058 2418 3062
rect 2438 3058 2442 3062
rect 2470 3058 2474 3062
rect 2502 3058 2506 3062
rect 2510 3058 2514 3062
rect 2582 3058 2586 3062
rect 2598 3058 2602 3062
rect 2606 3058 2610 3062
rect 2630 3058 2634 3062
rect 2718 3058 2722 3062
rect 2774 3058 2778 3062
rect 2814 3058 2818 3062
rect 2830 3058 2834 3062
rect 2846 3058 2850 3062
rect 2854 3058 2858 3062
rect 2878 3058 2882 3062
rect 2894 3058 2898 3062
rect 2982 3058 2986 3062
rect 3030 3058 3034 3062
rect 3062 3058 3066 3062
rect 3086 3058 3090 3062
rect 3094 3058 3098 3062
rect 3142 3058 3146 3062
rect 3174 3058 3178 3062
rect 3270 3059 3274 3063
rect 3494 3068 3498 3072
rect 3558 3068 3562 3072
rect 3598 3068 3602 3072
rect 3614 3068 3618 3072
rect 3654 3068 3658 3072
rect 3678 3068 3682 3072
rect 3710 3068 3714 3072
rect 3750 3068 3754 3072
rect 3782 3068 3786 3072
rect 3846 3068 3850 3072
rect 3894 3068 3898 3072
rect 3926 3068 3930 3072
rect 3974 3068 3978 3072
rect 4030 3068 4034 3072
rect 4118 3068 4122 3072
rect 4198 3068 4202 3072
rect 4262 3068 4266 3072
rect 4318 3068 4322 3072
rect 4494 3068 4498 3072
rect 4518 3068 4522 3072
rect 4526 3068 4530 3072
rect 4590 3068 4594 3072
rect 4598 3068 4602 3072
rect 4638 3068 4642 3072
rect 4742 3068 4746 3072
rect 4782 3068 4786 3072
rect 4870 3068 4874 3072
rect 4910 3068 4914 3072
rect 4942 3068 4946 3072
rect 4966 3068 4970 3072
rect 5030 3068 5034 3072
rect 5078 3068 5082 3072
rect 5198 3068 5202 3072
rect 5238 3068 5242 3072
rect 3318 3058 3322 3062
rect 3326 3058 3330 3062
rect 3350 3058 3354 3062
rect 3358 3058 3362 3062
rect 3390 3058 3394 3062
rect 3414 3058 3418 3062
rect 3454 3058 3458 3062
rect 3470 3058 3474 3062
rect 3542 3059 3546 3063
rect 3590 3058 3594 3062
rect 3622 3058 3626 3062
rect 3646 3058 3650 3062
rect 3686 3058 3690 3062
rect 3718 3058 3722 3062
rect 3742 3058 3746 3062
rect 3806 3058 3810 3062
rect 3902 3058 3906 3062
rect 3918 3058 3922 3062
rect 3966 3058 3970 3062
rect 3998 3058 4002 3062
rect 4022 3058 4026 3062
rect 4102 3059 4106 3063
rect 4182 3058 4186 3062
rect 4190 3058 4194 3062
rect 4206 3058 4210 3062
rect 4222 3058 4226 3062
rect 4262 3058 4266 3062
rect 4270 3058 4274 3062
rect 4310 3058 4314 3062
rect 4350 3059 4354 3063
rect 4438 3058 4442 3062
rect 4486 3058 4490 3062
rect 4606 3058 4610 3062
rect 4622 3058 4626 3062
rect 4638 3058 4642 3062
rect 4726 3059 4730 3063
rect 4766 3058 4770 3062
rect 4782 3058 4786 3062
rect 4854 3059 4858 3063
rect 4902 3058 4906 3062
rect 4934 3058 4938 3062
rect 4974 3058 4978 3062
rect 5038 3058 5042 3062
rect 5150 3058 5154 3062
rect 5214 3059 5218 3063
rect 1358 3048 1362 3052
rect 1406 3048 1410 3052
rect 1438 3048 1442 3052
rect 1446 3048 1450 3052
rect 1478 3048 1482 3052
rect 1590 3048 1594 3052
rect 1622 3048 1626 3052
rect 1686 3048 1690 3052
rect 1822 3048 1826 3052
rect 1878 3048 1882 3052
rect 2166 3048 2170 3052
rect 2542 3048 2546 3052
rect 2566 3048 2570 3052
rect 2622 3048 2626 3052
rect 2774 3048 2778 3052
rect 2814 3048 2818 3052
rect 3046 3048 3050 3052
rect 3366 3048 3370 3052
rect 3382 3048 3386 3052
rect 3470 3048 3474 3052
rect 3630 3048 3634 3052
rect 3702 3048 3706 3052
rect 3718 3048 3722 3052
rect 3734 3048 3738 3052
rect 3886 3048 3890 3052
rect 3902 3048 3906 3052
rect 3934 3048 3938 3052
rect 4006 3048 4010 3052
rect 4166 3048 4170 3052
rect 4222 3048 4226 3052
rect 4286 3048 4290 3052
rect 4454 3048 4458 3052
rect 4470 3048 4474 3052
rect 4502 3048 4506 3052
rect 4758 3048 4762 3052
rect 4918 3048 4922 3052
rect 534 3038 538 3042
rect 926 3038 930 3042
rect 1006 3038 1010 3042
rect 1102 3038 1106 3042
rect 1726 3038 1730 3042
rect 2782 3038 2786 3042
rect 2870 3038 2874 3042
rect 2942 3038 2946 3042
rect 4310 3038 4314 3042
rect 4790 3038 4794 3042
rect 4886 3038 4890 3042
rect 4902 3038 4906 3042
rect 550 3028 554 3032
rect 2102 3028 2106 3032
rect 4414 3028 4418 3032
rect 4510 3028 4514 3032
rect 62 3018 66 3022
rect 142 3018 146 3022
rect 454 3018 458 3022
rect 758 3018 762 3022
rect 1302 3018 1306 3022
rect 1318 3018 1322 3022
rect 1510 3018 1514 3022
rect 1574 3018 1578 3022
rect 1606 3018 1610 3022
rect 2158 3018 2162 3022
rect 2198 3018 2202 3022
rect 2526 3018 2530 3022
rect 2550 3018 2554 3022
rect 3030 3018 3034 3022
rect 3070 3018 3074 3022
rect 3110 3018 3114 3022
rect 3158 3018 3162 3022
rect 3198 3018 3202 3022
rect 3478 3018 3482 3022
rect 3686 3018 3690 3022
rect 3998 3018 4002 3022
rect 4022 3018 4026 3022
rect 4486 3018 4490 3022
rect 4614 3018 4618 3022
rect 4998 3018 5002 3022
rect 5094 3018 5098 3022
rect 5278 3018 5282 3022
rect 330 3003 334 3007
rect 337 3003 341 3007
rect 1354 3003 1358 3007
rect 1361 3003 1365 3007
rect 2386 3003 2390 3007
rect 2393 3003 2397 3007
rect 3402 3003 3406 3007
rect 3409 3003 3413 3007
rect 4426 3003 4430 3007
rect 4433 3003 4437 3007
rect 734 2988 738 2992
rect 782 2988 786 2992
rect 926 2988 930 2992
rect 1454 2988 1458 2992
rect 1582 2988 1586 2992
rect 1606 2988 1610 2992
rect 1798 2988 1802 2992
rect 1958 2988 1962 2992
rect 1990 2988 1994 2992
rect 2366 2988 2370 2992
rect 2470 2988 2474 2992
rect 2926 2988 2930 2992
rect 3014 2988 3018 2992
rect 3046 2988 3050 2992
rect 3454 2988 3458 2992
rect 3494 2988 3498 2992
rect 3710 2988 3714 2992
rect 3814 2988 3818 2992
rect 4062 2988 4066 2992
rect 4710 2988 4714 2992
rect 5110 2988 5114 2992
rect 5198 2988 5202 2992
rect 5262 2988 5266 2992
rect 3518 2978 3522 2982
rect 4006 2978 4010 2982
rect 4990 2978 4994 2982
rect 598 2968 602 2972
rect 1078 2968 1082 2972
rect 1686 2968 1690 2972
rect 2678 2968 2682 2972
rect 2710 2968 2714 2972
rect 2726 2968 2730 2972
rect 3190 2968 3194 2972
rect 3438 2968 3442 2972
rect 3678 2968 3682 2972
rect 3926 2968 3930 2972
rect 4158 2968 4162 2972
rect 4222 2968 4226 2972
rect 758 2958 762 2962
rect 1286 2958 1290 2962
rect 1342 2958 1346 2962
rect 1646 2958 1650 2962
rect 70 2947 74 2951
rect 150 2948 154 2952
rect 246 2948 250 2952
rect 310 2948 314 2952
rect 350 2948 354 2952
rect 374 2948 378 2952
rect 446 2948 450 2952
rect 542 2948 546 2952
rect 606 2948 610 2952
rect 638 2948 642 2952
rect 678 2948 682 2952
rect 686 2948 690 2952
rect 718 2948 722 2952
rect 750 2948 754 2952
rect 798 2948 802 2952
rect 854 2948 858 2952
rect 942 2948 946 2952
rect 982 2948 986 2952
rect 1006 2948 1010 2952
rect 1070 2948 1074 2952
rect 1150 2948 1154 2952
rect 1158 2948 1162 2952
rect 1190 2947 1194 2951
rect 1270 2948 1274 2952
rect 1318 2948 1322 2952
rect 1374 2948 1378 2952
rect 1390 2948 1394 2952
rect 1422 2948 1426 2952
rect 1470 2948 1474 2952
rect 1510 2948 1514 2952
rect 1590 2948 1594 2952
rect 1622 2948 1626 2952
rect 2022 2958 2026 2962
rect 2054 2958 2058 2962
rect 2102 2958 2106 2962
rect 2950 2958 2954 2962
rect 3254 2958 3258 2962
rect 4046 2958 4050 2962
rect 1662 2948 1666 2952
rect 1670 2948 1674 2952
rect 1726 2948 1730 2952
rect 1782 2948 1786 2952
rect 1830 2948 1834 2952
rect 1886 2948 1890 2952
rect 1910 2948 1914 2952
rect 1974 2948 1978 2952
rect 2006 2948 2010 2952
rect 2030 2948 2034 2952
rect 2174 2947 2178 2951
rect 2214 2948 2218 2952
rect 2238 2948 2242 2952
rect 2246 2948 2250 2952
rect 2254 2948 2258 2952
rect 2302 2948 2306 2952
rect 2334 2948 2338 2952
rect 2342 2948 2346 2952
rect 2350 2948 2354 2952
rect 2406 2948 2410 2952
rect 2422 2948 2426 2952
rect 2454 2948 2458 2952
rect 2502 2948 2506 2952
rect 2534 2948 2538 2952
rect 2566 2948 2570 2952
rect 2574 2948 2578 2952
rect 2582 2948 2586 2952
rect 2614 2948 2618 2952
rect 2646 2948 2650 2952
rect 2654 2948 2658 2952
rect 2702 2948 2706 2952
rect 2766 2948 2770 2952
rect 2838 2948 2842 2952
rect 2862 2948 2866 2952
rect 2966 2948 2970 2952
rect 2990 2948 2994 2952
rect 2998 2948 3002 2952
rect 3030 2948 3034 2952
rect 3070 2948 3074 2952
rect 3142 2948 3146 2952
rect 3198 2948 3202 2952
rect 3246 2948 3250 2952
rect 3302 2947 3306 2951
rect 3382 2948 3386 2952
rect 3478 2948 3482 2952
rect 3534 2948 3538 2952
rect 3566 2948 3570 2952
rect 3574 2948 3578 2952
rect 3638 2948 3642 2952
rect 3654 2948 3658 2952
rect 3750 2948 3754 2952
rect 3758 2948 3762 2952
rect 3766 2948 3770 2952
rect 3798 2948 3802 2952
rect 3862 2948 3866 2952
rect 3942 2948 3946 2952
rect 3990 2948 3994 2952
rect 4022 2948 4026 2952
rect 4078 2948 4082 2952
rect 4086 2948 4090 2952
rect 4142 2948 4146 2952
rect 4198 2958 4202 2962
rect 4342 2958 4346 2962
rect 4374 2958 4378 2962
rect 4430 2958 4434 2962
rect 4486 2958 4490 2962
rect 4678 2958 4682 2962
rect 4910 2958 4914 2962
rect 4198 2948 4202 2952
rect 4278 2948 4282 2952
rect 4334 2948 4338 2952
rect 4358 2948 4362 2952
rect 4390 2948 4394 2952
rect 4414 2948 4418 2952
rect 4422 2948 4426 2952
rect 4478 2948 4482 2952
rect 4502 2948 4506 2952
rect 4518 2948 4522 2952
rect 4526 2948 4530 2952
rect 4558 2948 4562 2952
rect 4622 2948 4626 2952
rect 4694 2948 4698 2952
rect 4758 2948 4762 2952
rect 4838 2948 4842 2952
rect 4846 2948 4850 2952
rect 4870 2948 4874 2952
rect 4894 2948 4898 2952
rect 4966 2958 4970 2962
rect 4926 2948 4930 2952
rect 4934 2948 4938 2952
rect 5038 2948 5042 2952
rect 5086 2948 5090 2952
rect 5094 2948 5098 2952
rect 5118 2948 5122 2952
rect 5150 2948 5154 2952
rect 5182 2948 5186 2952
rect 5302 2948 5306 2952
rect 62 2938 66 2942
rect 126 2938 130 2942
rect 222 2938 226 2942
rect 318 2938 322 2942
rect 390 2938 394 2942
rect 534 2938 538 2942
rect 614 2938 618 2942
rect 694 2938 698 2942
rect 814 2938 818 2942
rect 1094 2938 1098 2942
rect 1198 2938 1202 2942
rect 1262 2938 1266 2942
rect 1310 2938 1314 2942
rect 1326 2938 1330 2942
rect 1350 2938 1354 2942
rect 1366 2938 1370 2942
rect 1398 2938 1402 2942
rect 1486 2938 1490 2942
rect 1678 2938 1682 2942
rect 1766 2938 1770 2942
rect 1862 2938 1866 2942
rect 1998 2938 2002 2942
rect 2078 2938 2082 2942
rect 2206 2938 2210 2942
rect 2326 2938 2330 2942
rect 2446 2938 2450 2942
rect 2494 2938 2498 2942
rect 2510 2938 2514 2942
rect 2558 2938 2562 2942
rect 2638 2938 2642 2942
rect 2702 2938 2706 2942
rect 2934 2938 2938 2942
rect 2950 2938 2954 2942
rect 3094 2938 3098 2942
rect 3206 2938 3210 2942
rect 3222 2938 3226 2942
rect 3270 2938 3274 2942
rect 3286 2938 3290 2942
rect 3310 2938 3314 2942
rect 3374 2938 3378 2942
rect 3390 2938 3394 2942
rect 3422 2938 3426 2942
rect 3598 2938 3602 2942
rect 3718 2938 3722 2942
rect 3854 2938 3858 2942
rect 3950 2938 3954 2942
rect 4030 2938 4034 2942
rect 4134 2938 4138 2942
rect 4174 2938 4178 2942
rect 4190 2938 4194 2942
rect 4302 2938 4306 2942
rect 4350 2938 4354 2942
rect 4366 2938 4370 2942
rect 4398 2938 4402 2942
rect 4406 2938 4410 2942
rect 4510 2938 4514 2942
rect 4550 2938 4554 2942
rect 4574 2938 4578 2942
rect 4662 2938 4666 2942
rect 4734 2938 4738 2942
rect 4822 2938 4826 2942
rect 4886 2938 4890 2942
rect 4942 2938 4946 2942
rect 4958 2938 4962 2942
rect 4982 2938 4986 2942
rect 5046 2938 5050 2942
rect 5134 2938 5138 2942
rect 5174 2938 5178 2942
rect 5254 2938 5258 2942
rect 5294 2938 5298 2942
rect 102 2928 106 2932
rect 326 2928 330 2932
rect 374 2928 378 2932
rect 406 2928 410 2932
rect 438 2928 442 2932
rect 622 2928 626 2932
rect 654 2928 658 2932
rect 710 2928 714 2932
rect 766 2928 770 2932
rect 1054 2928 1058 2932
rect 1110 2928 1114 2932
rect 1142 2928 1146 2932
rect 1326 2928 1330 2932
rect 1438 2928 1442 2932
rect 1814 2928 1818 2932
rect 1982 2928 1986 2932
rect 2062 2928 2066 2932
rect 2174 2928 2178 2932
rect 2286 2928 2290 2932
rect 2390 2928 2394 2932
rect 2526 2928 2530 2932
rect 2558 2928 2562 2932
rect 2622 2928 2626 2932
rect 2670 2928 2674 2932
rect 3126 2928 3130 2932
rect 3222 2928 3226 2932
rect 3230 2928 3234 2932
rect 3246 2928 3250 2932
rect 3974 2928 3978 2932
rect 4102 2928 4106 2932
rect 4126 2928 4130 2932
rect 4318 2928 4322 2932
rect 4334 2928 4338 2932
rect 4374 2928 4378 2932
rect 4686 2928 4690 2932
rect 4854 2928 4858 2932
rect 5270 2928 5274 2932
rect 5278 2928 5282 2932
rect 6 2918 10 2922
rect 110 2918 114 2922
rect 206 2918 210 2922
rect 302 2918 306 2922
rect 398 2918 402 2922
rect 502 2918 506 2922
rect 670 2918 674 2922
rect 702 2918 706 2922
rect 910 2918 914 2922
rect 926 2918 930 2922
rect 1038 2918 1042 2922
rect 1086 2918 1090 2922
rect 1254 2918 1258 2922
rect 1302 2918 1306 2922
rect 1406 2918 1410 2922
rect 1798 2918 1802 2922
rect 1822 2918 1826 2922
rect 1942 2918 1946 2922
rect 2270 2918 2274 2922
rect 2318 2918 2322 2922
rect 2438 2918 2442 2922
rect 2486 2918 2490 2922
rect 2598 2918 2602 2922
rect 2630 2918 2634 2922
rect 2950 2918 2954 2922
rect 3014 2918 3018 2922
rect 3254 2918 3258 2922
rect 3366 2918 3370 2922
rect 3494 2918 3498 2922
rect 3550 2918 3554 2922
rect 3590 2918 3594 2922
rect 3782 2918 3786 2922
rect 3958 2918 3962 2922
rect 4046 2918 4050 2922
rect 4094 2918 4098 2922
rect 4118 2918 4122 2922
rect 4206 2918 4210 2922
rect 4462 2918 4466 2922
rect 4486 2918 4490 2922
rect 4710 2918 4714 2922
rect 4974 2918 4978 2922
rect 5166 2918 5170 2922
rect 5286 2918 5290 2922
rect 850 2903 854 2907
rect 857 2903 861 2907
rect 1874 2903 1878 2907
rect 1881 2903 1885 2907
rect 2890 2903 2894 2907
rect 2897 2903 2901 2907
rect 3922 2903 3926 2907
rect 3929 2903 3933 2907
rect 4938 2903 4942 2907
rect 4945 2903 4949 2907
rect 94 2888 98 2892
rect 166 2888 170 2892
rect 398 2888 402 2892
rect 494 2888 498 2892
rect 558 2888 562 2892
rect 646 2888 650 2892
rect 870 2888 874 2892
rect 902 2888 906 2892
rect 982 2888 986 2892
rect 1254 2888 1258 2892
rect 1894 2888 1898 2892
rect 2030 2888 2034 2892
rect 2094 2888 2098 2892
rect 2182 2888 2186 2892
rect 2350 2888 2354 2892
rect 2382 2888 2386 2892
rect 2478 2888 2482 2892
rect 2606 2888 2610 2892
rect 3150 2888 3154 2892
rect 3262 2888 3266 2892
rect 3286 2888 3290 2892
rect 3334 2888 3338 2892
rect 3470 2888 3474 2892
rect 3510 2888 3514 2892
rect 3526 2888 3530 2892
rect 3566 2888 3570 2892
rect 3638 2888 3642 2892
rect 3806 2888 3810 2892
rect 3838 2888 3842 2892
rect 4166 2888 4170 2892
rect 4190 2888 4194 2892
rect 4446 2888 4450 2892
rect 4518 2888 4522 2892
rect 4982 2888 4986 2892
rect 5102 2888 5106 2892
rect 5294 2888 5298 2892
rect 326 2878 330 2882
rect 342 2878 346 2882
rect 534 2878 538 2882
rect 198 2868 202 2872
rect 214 2868 218 2872
rect 254 2868 258 2872
rect 262 2868 266 2872
rect 318 2868 322 2872
rect 374 2868 378 2872
rect 430 2868 434 2872
rect 438 2868 442 2872
rect 526 2868 530 2872
rect 582 2868 586 2872
rect 590 2868 594 2872
rect 622 2868 626 2872
rect 638 2868 642 2872
rect 662 2878 666 2882
rect 686 2878 690 2882
rect 934 2878 938 2882
rect 942 2878 946 2882
rect 1014 2878 1018 2882
rect 1038 2878 1042 2882
rect 1078 2878 1082 2882
rect 1502 2878 1506 2882
rect 1582 2878 1586 2882
rect 1798 2878 1802 2882
rect 2086 2878 2090 2882
rect 2574 2878 2578 2882
rect 2806 2878 2810 2882
rect 3318 2878 3322 2882
rect 3558 2878 3562 2882
rect 3734 2878 3738 2882
rect 4158 2878 4162 2882
rect 4334 2878 4338 2882
rect 4494 2878 4498 2882
rect 4510 2878 4514 2882
rect 4558 2878 4562 2882
rect 742 2868 746 2872
rect 782 2868 786 2872
rect 798 2868 802 2872
rect 894 2868 898 2872
rect 958 2868 962 2872
rect 974 2868 978 2872
rect 1046 2868 1050 2872
rect 1102 2868 1106 2872
rect 1142 2868 1146 2872
rect 1158 2868 1162 2872
rect 1174 2868 1178 2872
rect 1278 2868 1282 2872
rect 1310 2868 1314 2872
rect 1318 2868 1322 2872
rect 1438 2868 1442 2872
rect 1486 2868 1490 2872
rect 1598 2868 1602 2872
rect 1758 2868 1762 2872
rect 1966 2868 1970 2872
rect 2046 2868 2050 2872
rect 2110 2868 2114 2872
rect 2142 2868 2146 2872
rect 2150 2868 2154 2872
rect 2278 2868 2282 2872
rect 2294 2868 2298 2872
rect 2366 2868 2370 2872
rect 2558 2868 2562 2872
rect 2614 2868 2618 2872
rect 2638 2868 2642 2872
rect 2726 2868 2730 2872
rect 2862 2868 2866 2872
rect 2870 2868 2874 2872
rect 3006 2868 3010 2872
rect 3054 2868 3058 2872
rect 3166 2868 3170 2872
rect 3238 2868 3242 2872
rect 3278 2868 3282 2872
rect 3342 2868 3346 2872
rect 3550 2868 3554 2872
rect 3574 2868 3578 2872
rect 3750 2868 3754 2872
rect 3830 2868 3834 2872
rect 3870 2868 3874 2872
rect 3990 2868 3994 2872
rect 4054 2868 4058 2872
rect 4158 2868 4162 2872
rect 4174 2868 4178 2872
rect 4414 2868 4418 2872
rect 4486 2868 4490 2872
rect 4526 2868 4530 2872
rect 4598 2878 4602 2882
rect 4750 2878 4754 2882
rect 5046 2878 5050 2882
rect 4582 2868 4586 2872
rect 4678 2868 4682 2872
rect 4694 2868 4698 2872
rect 4766 2868 4770 2872
rect 4806 2868 4810 2872
rect 4846 2868 4850 2872
rect 4862 2868 4866 2872
rect 4894 2868 4898 2872
rect 4942 2868 4946 2872
rect 5062 2868 5066 2872
rect 5078 2868 5082 2872
rect 38 2858 42 2862
rect 62 2858 66 2862
rect 110 2858 114 2862
rect 134 2858 138 2862
rect 142 2858 146 2862
rect 158 2858 162 2862
rect 182 2858 186 2862
rect 190 2858 194 2862
rect 206 2858 210 2862
rect 246 2858 250 2862
rect 270 2858 274 2862
rect 310 2858 314 2862
rect 358 2858 362 2862
rect 382 2858 386 2862
rect 446 2858 450 2862
rect 502 2858 506 2862
rect 534 2858 538 2862
rect 558 2858 562 2862
rect 574 2858 578 2862
rect 598 2858 602 2862
rect 614 2858 618 2862
rect 630 2858 634 2862
rect 678 2858 682 2862
rect 702 2858 706 2862
rect 718 2858 722 2862
rect 750 2858 754 2862
rect 806 2858 810 2862
rect 870 2858 874 2862
rect 918 2858 922 2862
rect 958 2858 962 2862
rect 966 2858 970 2862
rect 998 2858 1002 2862
rect 1014 2858 1018 2862
rect 1094 2858 1098 2862
rect 1110 2858 1114 2862
rect 1150 2858 1154 2862
rect 1190 2859 1194 2863
rect 1286 2858 1290 2862
rect 1302 2858 1306 2862
rect 1374 2858 1378 2862
rect 1390 2858 1394 2862
rect 1454 2859 1458 2863
rect 1526 2858 1530 2862
rect 1558 2858 1562 2862
rect 1566 2858 1570 2862
rect 1622 2858 1626 2862
rect 1638 2858 1642 2862
rect 1702 2858 1706 2862
rect 1710 2858 1714 2862
rect 1734 2858 1738 2862
rect 1742 2858 1746 2862
rect 1750 2858 1754 2862
rect 1782 2858 1786 2862
rect 1830 2859 1834 2863
rect 1862 2858 1866 2862
rect 1934 2858 1938 2862
rect 1974 2858 1978 2862
rect 1998 2858 2002 2862
rect 2038 2858 2042 2862
rect 2070 2858 2074 2862
rect 2110 2858 2114 2862
rect 2134 2858 2138 2862
rect 2158 2858 2162 2862
rect 2214 2858 2218 2862
rect 2246 2859 2250 2863
rect 2326 2858 2330 2862
rect 2342 2858 2346 2862
rect 2422 2858 2426 2862
rect 2438 2858 2442 2862
rect 2510 2858 2514 2862
rect 2542 2859 2546 2863
rect 2590 2858 2594 2862
rect 2622 2858 2626 2862
rect 2654 2859 2658 2863
rect 2686 2858 2690 2862
rect 2750 2858 2754 2862
rect 2766 2858 2770 2862
rect 2790 2858 2794 2862
rect 2822 2858 2826 2862
rect 2830 2858 2834 2862
rect 2838 2858 2842 2862
rect 2862 2858 2866 2862
rect 2942 2858 2946 2862
rect 2966 2858 2970 2862
rect 3094 2858 3098 2862
rect 3158 2858 3162 2862
rect 3190 2858 3194 2862
rect 3198 2858 3202 2862
rect 3206 2858 3210 2862
rect 3246 2858 3250 2862
rect 3270 2858 3274 2862
rect 3302 2858 3306 2862
rect 3350 2858 3354 2862
rect 3366 2858 3370 2862
rect 3382 2858 3386 2862
rect 3390 2858 3394 2862
rect 3414 2858 3418 2862
rect 3422 2858 3426 2862
rect 3446 2858 3450 2862
rect 3494 2858 3498 2862
rect 3542 2858 3546 2862
rect 3582 2858 3586 2862
rect 3590 2858 3594 2862
rect 3622 2858 3626 2862
rect 3630 2858 3634 2862
rect 3678 2858 3682 2862
rect 3694 2858 3698 2862
rect 3782 2858 3786 2862
rect 3790 2858 3794 2862
rect 3854 2858 3858 2862
rect 3902 2858 3906 2862
rect 3998 2858 4002 2862
rect 4022 2858 4026 2862
rect 4030 2858 4034 2862
rect 4102 2858 4106 2862
rect 4126 2859 4130 2863
rect 4182 2858 4186 2862
rect 4222 2858 4226 2862
rect 4230 2858 4234 2862
rect 4294 2858 4298 2862
rect 4318 2858 4322 2862
rect 4326 2858 4330 2862
rect 4406 2858 4410 2862
rect 4478 2858 4482 2862
rect 4534 2858 4538 2862
rect 4542 2858 4546 2862
rect 4574 2858 4578 2862
rect 4590 2858 4594 2862
rect 4646 2858 4650 2862
rect 4774 2858 4778 2862
rect 4798 2858 4802 2862
rect 4830 2858 4834 2862
rect 4838 2858 4842 2862
rect 4854 2858 4858 2862
rect 4902 2858 4906 2862
rect 4958 2858 4962 2862
rect 5022 2858 5026 2862
rect 5086 2858 5090 2862
rect 5142 2858 5146 2862
rect 5166 2858 5170 2862
rect 5230 2859 5234 2863
rect 230 2848 234 2852
rect 270 2848 274 2852
rect 294 2848 298 2852
rect 358 2848 362 2852
rect 398 2848 402 2852
rect 502 2848 506 2852
rect 558 2848 562 2852
rect 734 2848 738 2852
rect 766 2848 770 2852
rect 1070 2848 1074 2852
rect 1126 2848 1130 2852
rect 1262 2848 1266 2852
rect 1686 2848 1690 2852
rect 1774 2848 1778 2852
rect 2094 2848 2098 2852
rect 2118 2848 2122 2852
rect 2174 2848 2178 2852
rect 2342 2848 2346 2852
rect 2766 2848 2770 2852
rect 2774 2848 2778 2852
rect 3222 2848 3226 2852
rect 3262 2848 3266 2852
rect 3326 2848 3330 2852
rect 3526 2848 3530 2852
rect 4038 2848 4042 2852
rect 4790 2848 4794 2852
rect 4878 2848 4882 2852
rect 4958 2848 4962 2852
rect 4974 2848 4978 2852
rect 550 2838 554 2842
rect 846 2838 850 2842
rect 2062 2838 2066 2842
rect 3654 2838 3658 2842
rect 4310 2838 4314 2842
rect 4774 2828 4778 2832
rect 118 2818 122 2822
rect 494 2818 498 2822
rect 614 2818 618 2822
rect 718 2818 722 2822
rect 750 2818 754 2822
rect 862 2818 866 2822
rect 1054 2818 1058 2822
rect 1094 2818 1098 2822
rect 1422 2818 1426 2822
rect 1518 2818 1522 2822
rect 1550 2818 1554 2822
rect 1574 2818 1578 2822
rect 1926 2818 1930 2822
rect 2158 2818 2162 2822
rect 2790 2818 2794 2822
rect 3030 2818 3034 2822
rect 3438 2818 3442 2822
rect 3606 2818 3610 2822
rect 3806 2818 3810 2822
rect 3982 2818 3986 2822
rect 4046 2818 4050 2822
rect 4062 2818 4066 2822
rect 4502 2818 4506 2822
rect 4918 2818 4922 2822
rect 5110 2818 5114 2822
rect 330 2803 334 2807
rect 337 2803 341 2807
rect 1354 2803 1358 2807
rect 1361 2803 1365 2807
rect 2386 2803 2390 2807
rect 2393 2803 2397 2807
rect 3402 2803 3406 2807
rect 3409 2803 3413 2807
rect 4426 2803 4430 2807
rect 4433 2803 4437 2807
rect 110 2788 114 2792
rect 710 2788 714 2792
rect 1382 2788 1386 2792
rect 1534 2788 1538 2792
rect 1822 2788 1826 2792
rect 2118 2788 2122 2792
rect 2206 2788 2210 2792
rect 2774 2788 2778 2792
rect 2854 2788 2858 2792
rect 3014 2788 3018 2792
rect 3038 2788 3042 2792
rect 3078 2788 3082 2792
rect 3134 2788 3138 2792
rect 3278 2788 3282 2792
rect 3638 2788 3642 2792
rect 3782 2788 3786 2792
rect 4190 2788 4194 2792
rect 5014 2788 5018 2792
rect 5094 2788 5098 2792
rect 5214 2788 5218 2792
rect 5222 2788 5226 2792
rect 5302 2788 5306 2792
rect 334 2778 338 2782
rect 3646 2778 3650 2782
rect 382 2768 386 2772
rect 510 2768 514 2772
rect 574 2768 578 2772
rect 854 2768 858 2772
rect 1350 2768 1354 2772
rect 1406 2768 1410 2772
rect 1446 2768 1450 2772
rect 1742 2768 1746 2772
rect 2150 2768 2154 2772
rect 2390 2768 2394 2772
rect 3470 2768 3474 2772
rect 3910 2768 3914 2772
rect 4558 2768 4562 2772
rect 4742 2768 4746 2772
rect 4798 2768 4802 2772
rect 4926 2768 4930 2772
rect 4990 2768 4994 2772
rect 142 2758 146 2762
rect 38 2748 42 2752
rect 62 2748 66 2752
rect 134 2748 138 2752
rect 198 2748 202 2752
rect 278 2748 282 2752
rect 366 2748 370 2752
rect 646 2758 650 2762
rect 694 2758 698 2762
rect 902 2758 906 2762
rect 934 2758 938 2762
rect 950 2758 954 2762
rect 966 2758 970 2762
rect 1078 2758 1082 2762
rect 1094 2758 1098 2762
rect 1126 2758 1130 2762
rect 1158 2758 1162 2762
rect 406 2748 410 2752
rect 454 2748 458 2752
rect 518 2748 522 2752
rect 566 2748 570 2752
rect 582 2748 586 2752
rect 590 2748 594 2752
rect 630 2748 634 2752
rect 662 2748 666 2752
rect 686 2748 690 2752
rect 710 2748 714 2752
rect 734 2748 738 2752
rect 750 2748 754 2752
rect 806 2748 810 2752
rect 878 2748 882 2752
rect 894 2748 898 2752
rect 918 2748 922 2752
rect 926 2748 930 2752
rect 950 2748 954 2752
rect 1006 2748 1010 2752
rect 1070 2748 1074 2752
rect 1110 2748 1114 2752
rect 1142 2748 1146 2752
rect 1158 2748 1162 2752
rect 118 2738 122 2742
rect 158 2738 162 2742
rect 270 2738 274 2742
rect 358 2738 362 2742
rect 390 2738 394 2742
rect 414 2738 418 2742
rect 430 2738 434 2742
rect 478 2738 482 2742
rect 526 2738 530 2742
rect 598 2738 602 2742
rect 622 2738 626 2742
rect 718 2738 722 2742
rect 726 2738 730 2742
rect 742 2738 746 2742
rect 758 2738 762 2742
rect 798 2738 802 2742
rect 870 2738 874 2742
rect 910 2738 914 2742
rect 1190 2747 1194 2751
rect 1294 2748 1298 2752
rect 1318 2748 1322 2752
rect 1382 2748 1386 2752
rect 1422 2748 1426 2752
rect 1438 2748 1442 2752
rect 1470 2758 1474 2762
rect 1574 2758 1578 2762
rect 1486 2748 1490 2752
rect 1518 2748 1522 2752
rect 1542 2748 1546 2752
rect 1558 2748 1562 2752
rect 1574 2748 1578 2752
rect 1614 2748 1618 2752
rect 1638 2748 1642 2752
rect 1686 2748 1690 2752
rect 1758 2758 1762 2762
rect 2030 2758 2034 2762
rect 2038 2758 2042 2762
rect 2166 2758 2170 2762
rect 2174 2758 2178 2762
rect 2294 2758 2298 2762
rect 2502 2758 2506 2762
rect 2518 2758 2522 2762
rect 2558 2758 2562 2762
rect 2758 2758 2762 2762
rect 2822 2758 2826 2762
rect 3182 2758 3186 2762
rect 3222 2758 3226 2762
rect 1734 2748 1738 2752
rect 1774 2748 1778 2752
rect 1790 2748 1794 2752
rect 1806 2748 1810 2752
rect 1830 2748 1834 2752
rect 1886 2748 1890 2752
rect 1942 2748 1946 2752
rect 1966 2748 1970 2752
rect 2014 2748 2018 2752
rect 2038 2748 2042 2752
rect 2062 2748 2066 2752
rect 2094 2748 2098 2752
rect 2126 2748 2130 2752
rect 2134 2748 2138 2752
rect 2150 2748 2154 2752
rect 2270 2748 2274 2752
rect 2278 2748 2282 2752
rect 982 2738 986 2742
rect 1070 2738 1074 2742
rect 1102 2738 1106 2742
rect 1134 2738 1138 2742
rect 1174 2738 1178 2742
rect 1270 2738 1274 2742
rect 1374 2738 1378 2742
rect 1430 2738 1434 2742
rect 1438 2738 1442 2742
rect 1494 2738 1498 2742
rect 1542 2738 1546 2742
rect 1550 2738 1554 2742
rect 1678 2738 1682 2742
rect 1710 2738 1714 2742
rect 1758 2738 1762 2742
rect 1782 2738 1786 2742
rect 1798 2738 1802 2742
rect 1838 2738 1842 2742
rect 2006 2738 2010 2742
rect 2070 2738 2074 2742
rect 2142 2738 2146 2742
rect 2190 2738 2194 2742
rect 2262 2738 2266 2742
rect 2326 2747 2330 2751
rect 2406 2748 2410 2752
rect 2446 2748 2450 2752
rect 2478 2748 2482 2752
rect 2486 2748 2490 2752
rect 2494 2748 2498 2752
rect 2534 2748 2538 2752
rect 2542 2748 2546 2752
rect 2582 2748 2586 2752
rect 2598 2748 2602 2752
rect 2606 2748 2610 2752
rect 2630 2748 2634 2752
rect 2678 2748 2682 2752
rect 2758 2748 2762 2752
rect 2774 2748 2778 2752
rect 2790 2748 2794 2752
rect 2870 2748 2874 2752
rect 2918 2748 2922 2752
rect 2926 2748 2930 2752
rect 2958 2748 2962 2752
rect 2966 2748 2970 2752
rect 2998 2748 3002 2752
rect 3062 2748 3066 2752
rect 3094 2748 3098 2752
rect 3150 2748 3154 2752
rect 3158 2748 3162 2752
rect 3230 2748 3234 2752
rect 3262 2748 3266 2752
rect 3302 2748 3306 2752
rect 3414 2748 3418 2752
rect 3478 2748 3482 2752
rect 3502 2748 3506 2752
rect 3526 2748 3530 2752
rect 3566 2748 3570 2752
rect 3678 2748 3682 2752
rect 3710 2747 3714 2751
rect 3766 2748 3770 2752
rect 3798 2748 3802 2752
rect 3870 2748 3874 2752
rect 3886 2748 3890 2752
rect 3942 2748 3946 2752
rect 3950 2748 3954 2752
rect 3998 2748 4002 2752
rect 4022 2758 4026 2762
rect 4094 2758 4098 2762
rect 4126 2758 4130 2762
rect 4142 2758 4146 2762
rect 4158 2758 4162 2762
rect 4206 2758 4210 2762
rect 4222 2758 4226 2762
rect 4238 2758 4242 2762
rect 4294 2758 4298 2762
rect 4054 2748 4058 2752
rect 4078 2748 4082 2752
rect 4086 2748 4090 2752
rect 4110 2748 4114 2752
rect 4142 2748 4146 2752
rect 4166 2748 4170 2752
rect 4174 2748 4178 2752
rect 4230 2748 4234 2752
rect 4254 2748 4258 2752
rect 4278 2748 4282 2752
rect 4334 2758 4338 2762
rect 4606 2758 4610 2762
rect 4670 2758 4674 2762
rect 4686 2758 4690 2762
rect 4702 2758 4706 2762
rect 4758 2758 4762 2762
rect 4318 2748 4322 2752
rect 4374 2748 4378 2752
rect 4486 2748 4490 2752
rect 4542 2748 4546 2752
rect 4574 2748 4578 2752
rect 4582 2748 4586 2752
rect 4614 2748 4618 2752
rect 4654 2748 4658 2752
rect 4686 2748 4690 2752
rect 4710 2748 4714 2752
rect 2286 2738 2290 2742
rect 2310 2738 2314 2742
rect 2438 2738 2442 2742
rect 2526 2738 2530 2742
rect 2542 2738 2546 2742
rect 2590 2738 2594 2742
rect 2638 2738 2642 2742
rect 2686 2738 2690 2742
rect 2782 2738 2786 2742
rect 2790 2738 2794 2742
rect 2846 2738 2850 2742
rect 2886 2738 2890 2742
rect 2934 2738 2938 2742
rect 2950 2738 2954 2742
rect 2990 2738 2994 2742
rect 3126 2738 3130 2742
rect 3206 2738 3210 2742
rect 3358 2738 3362 2742
rect 3390 2738 3394 2742
rect 3518 2738 3522 2742
rect 3542 2738 3546 2742
rect 3806 2738 3810 2742
rect 3878 2738 3882 2742
rect 3958 2738 3962 2742
rect 3966 2738 3970 2742
rect 3982 2738 3986 2742
rect 4022 2738 4026 2742
rect 4038 2738 4042 2742
rect 4118 2738 4122 2742
rect 4150 2738 4154 2742
rect 4182 2738 4186 2742
rect 4230 2738 4234 2742
rect 4246 2738 4250 2742
rect 4262 2738 4266 2742
rect 4270 2738 4274 2742
rect 4310 2738 4314 2742
rect 4326 2738 4330 2742
rect 4414 2738 4418 2742
rect 174 2728 178 2732
rect 534 2728 538 2732
rect 550 2728 554 2732
rect 606 2728 610 2732
rect 638 2728 642 2732
rect 1502 2728 1506 2732
rect 1526 2728 1530 2732
rect 1702 2728 1706 2732
rect 1854 2728 1858 2732
rect 1902 2728 1906 2732
rect 2086 2728 2090 2732
rect 2510 2728 2514 2732
rect 2558 2728 2562 2732
rect 2814 2728 2818 2732
rect 3174 2728 3178 2732
rect 3494 2728 3498 2732
rect 4526 2738 4530 2742
rect 4590 2738 4594 2742
rect 4622 2738 4626 2742
rect 4646 2738 4650 2742
rect 4710 2738 4714 2742
rect 4734 2738 4738 2742
rect 4758 2748 4762 2752
rect 4894 2758 4898 2762
rect 4958 2758 4962 2762
rect 4782 2748 4786 2752
rect 4854 2748 4858 2752
rect 4910 2748 4914 2752
rect 4974 2748 4978 2752
rect 5054 2758 5058 2762
rect 5014 2748 5018 2752
rect 5038 2748 5042 2752
rect 5070 2748 5074 2752
rect 5086 2748 5090 2752
rect 5126 2748 5130 2752
rect 5134 2748 5138 2752
rect 5190 2748 5194 2752
rect 5254 2748 5258 2752
rect 5262 2748 5266 2752
rect 4790 2738 4794 2742
rect 4878 2738 4882 2742
rect 4918 2738 4922 2742
rect 4926 2738 4930 2742
rect 4966 2738 4970 2742
rect 5022 2738 5026 2742
rect 5030 2738 5034 2742
rect 5086 2738 5090 2742
rect 5198 2738 5202 2742
rect 5238 2738 5242 2742
rect 5278 2738 5282 2742
rect 3662 2728 3666 2732
rect 3982 2728 3986 2732
rect 4094 2728 4098 2732
rect 4198 2728 4202 2732
rect 4478 2728 4482 2732
rect 4638 2728 4642 2732
rect 5214 2728 5218 2732
rect 5230 2728 5234 2732
rect 5238 2728 5242 2732
rect 5286 2728 5290 2732
rect 238 2718 242 2722
rect 614 2718 618 2722
rect 670 2718 674 2722
rect 1062 2718 1066 2722
rect 1126 2718 1130 2722
rect 1254 2718 1258 2722
rect 1510 2718 1514 2722
rect 1742 2718 1746 2722
rect 1998 2718 2002 2722
rect 2046 2718 2050 2722
rect 2078 2718 2082 2722
rect 2182 2718 2186 2722
rect 2470 2718 2474 2722
rect 2566 2718 2570 2722
rect 2806 2718 2810 2722
rect 2830 2718 2834 2722
rect 2854 2718 2858 2722
rect 2934 2718 2938 2722
rect 3166 2718 3170 2722
rect 3182 2718 3186 2722
rect 3222 2718 3226 2722
rect 3246 2718 3250 2722
rect 3750 2718 3754 2722
rect 3910 2718 3914 2722
rect 3974 2718 3978 2722
rect 4062 2718 4066 2722
rect 4446 2718 4450 2722
rect 4598 2718 4602 2722
rect 4630 2718 4634 2722
rect 4750 2718 4754 2722
rect 4766 2718 4770 2722
rect 4894 2718 4898 2722
rect 850 2703 854 2707
rect 857 2703 861 2707
rect 1874 2703 1878 2707
rect 1881 2703 1885 2707
rect 2890 2703 2894 2707
rect 2897 2703 2901 2707
rect 3922 2703 3926 2707
rect 3929 2703 3933 2707
rect 4938 2703 4942 2707
rect 4945 2703 4949 2707
rect 94 2688 98 2692
rect 142 2688 146 2692
rect 198 2688 202 2692
rect 550 2688 554 2692
rect 590 2688 594 2692
rect 750 2688 754 2692
rect 822 2688 826 2692
rect 902 2688 906 2692
rect 1070 2688 1074 2692
rect 1142 2688 1146 2692
rect 1206 2688 1210 2692
rect 1326 2688 1330 2692
rect 1582 2688 1586 2692
rect 1614 2688 1618 2692
rect 1726 2688 1730 2692
rect 1750 2688 1754 2692
rect 1790 2688 1794 2692
rect 1814 2688 1818 2692
rect 2190 2688 2194 2692
rect 2478 2688 2482 2692
rect 2582 2688 2586 2692
rect 2598 2688 2602 2692
rect 2638 2688 2642 2692
rect 2742 2688 2746 2692
rect 2846 2688 2850 2692
rect 2862 2688 2866 2692
rect 2942 2688 2946 2692
rect 3014 2688 3018 2692
rect 3110 2688 3114 2692
rect 3238 2688 3242 2692
rect 3270 2688 3274 2692
rect 3334 2688 3338 2692
rect 3446 2688 3450 2692
rect 3702 2688 3706 2692
rect 3942 2688 3946 2692
rect 3958 2688 3962 2692
rect 4278 2688 4282 2692
rect 4438 2688 4442 2692
rect 4694 2688 4698 2692
rect 4742 2688 4746 2692
rect 5078 2688 5082 2692
rect 5286 2688 5290 2692
rect 190 2678 194 2682
rect 222 2678 226 2682
rect 238 2678 242 2682
rect 350 2678 354 2682
rect 478 2678 482 2682
rect 582 2678 586 2682
rect 638 2678 642 2682
rect 742 2678 746 2682
rect 758 2678 762 2682
rect 798 2678 802 2682
rect 814 2678 818 2682
rect 854 2678 858 2682
rect 942 2678 946 2682
rect 1022 2678 1026 2682
rect 102 2668 106 2672
rect 126 2668 130 2672
rect 150 2668 154 2672
rect 190 2668 194 2672
rect 206 2668 210 2672
rect 246 2668 250 2672
rect 270 2668 274 2672
rect 302 2668 306 2672
rect 422 2668 426 2672
rect 574 2668 578 2672
rect 598 2668 602 2672
rect 710 2668 714 2672
rect 1150 2678 1154 2682
rect 1406 2678 1410 2682
rect 1574 2678 1578 2682
rect 1622 2678 1626 2682
rect 1646 2678 1650 2682
rect 1686 2678 1690 2682
rect 1734 2678 1738 2682
rect 1782 2678 1786 2682
rect 1822 2678 1826 2682
rect 1878 2678 1882 2682
rect 2046 2678 2050 2682
rect 2054 2678 2058 2682
rect 2070 2678 2074 2682
rect 2166 2678 2170 2682
rect 2182 2678 2186 2682
rect 2342 2678 2346 2682
rect 2670 2678 2674 2682
rect 2750 2678 2754 2682
rect 3510 2678 3514 2682
rect 3686 2678 3690 2682
rect 3934 2678 3938 2682
rect 4382 2678 4386 2682
rect 4518 2678 4522 2682
rect 4758 2678 4762 2682
rect 4806 2678 4810 2682
rect 4894 2678 4898 2682
rect 5086 2678 5090 2682
rect 790 2668 794 2672
rect 854 2668 858 2672
rect 870 2668 874 2672
rect 910 2668 914 2672
rect 1094 2668 1098 2672
rect 1110 2668 1114 2672
rect 1118 2668 1122 2672
rect 1174 2668 1178 2672
rect 1190 2668 1194 2672
rect 1302 2668 1306 2672
rect 1334 2668 1338 2672
rect 1358 2668 1362 2672
rect 1390 2668 1394 2672
rect 1406 2668 1410 2672
rect 1414 2668 1418 2672
rect 1470 2668 1474 2672
rect 1518 2668 1522 2672
rect 1606 2668 1610 2672
rect 1654 2668 1658 2672
rect 1710 2668 1714 2672
rect 1774 2668 1778 2672
rect 1838 2668 1842 2672
rect 1910 2668 1914 2672
rect 1998 2668 2002 2672
rect 2102 2668 2106 2672
rect 2110 2668 2114 2672
rect 2126 2668 2130 2672
rect 2142 2668 2146 2672
rect 2206 2668 2210 2672
rect 2214 2668 2218 2672
rect 2246 2668 2250 2672
rect 2278 2668 2282 2672
rect 2422 2668 2426 2672
rect 2446 2668 2450 2672
rect 2502 2668 2506 2672
rect 2686 2668 2690 2672
rect 2766 2668 2770 2672
rect 3030 2668 3034 2672
rect 3078 2668 3082 2672
rect 3134 2668 3138 2672
rect 3294 2668 3298 2672
rect 3342 2668 3346 2672
rect 3526 2668 3530 2672
rect 3542 2668 3546 2672
rect 3590 2668 3594 2672
rect 3726 2668 3730 2672
rect 3758 2668 3762 2672
rect 3830 2668 3834 2672
rect 3854 2668 3858 2672
rect 3862 2668 3866 2672
rect 3878 2668 3882 2672
rect 3910 2668 3914 2672
rect 4166 2668 4170 2672
rect 4382 2668 4386 2672
rect 4462 2668 4466 2672
rect 4558 2668 4562 2672
rect 4582 2668 4586 2672
rect 4630 2668 4634 2672
rect 4670 2668 4674 2672
rect 4718 2668 4722 2672
rect 4782 2668 4786 2672
rect 4838 2668 4842 2672
rect 4870 2668 4874 2672
rect 4950 2668 4954 2672
rect 5062 2668 5066 2672
rect 38 2658 42 2662
rect 62 2658 66 2662
rect 110 2658 114 2662
rect 158 2658 162 2662
rect 182 2658 186 2662
rect 214 2658 218 2662
rect 222 2658 226 2662
rect 238 2658 242 2662
rect 302 2658 306 2662
rect 350 2659 354 2663
rect 430 2658 434 2662
rect 446 2658 450 2662
rect 478 2659 482 2663
rect 566 2658 570 2662
rect 606 2658 610 2662
rect 646 2658 650 2662
rect 718 2658 722 2662
rect 726 2658 730 2662
rect 758 2658 762 2662
rect 782 2658 786 2662
rect 830 2658 834 2662
rect 838 2658 842 2662
rect 886 2658 890 2662
rect 918 2658 922 2662
rect 958 2658 962 2662
rect 990 2659 994 2663
rect 1022 2658 1026 2662
rect 1078 2658 1082 2662
rect 1102 2658 1106 2662
rect 1126 2658 1130 2662
rect 1142 2658 1146 2662
rect 1166 2658 1170 2662
rect 1182 2658 1186 2662
rect 1246 2658 1250 2662
rect 1270 2659 1274 2663
rect 1310 2658 1314 2662
rect 1326 2658 1330 2662
rect 1350 2658 1354 2662
rect 1366 2658 1370 2662
rect 1422 2658 1426 2662
rect 1454 2658 1458 2662
rect 1462 2658 1466 2662
rect 1502 2659 1506 2663
rect 1590 2658 1594 2662
rect 1598 2658 1602 2662
rect 1630 2658 1634 2662
rect 1686 2658 1690 2662
rect 1702 2658 1706 2662
rect 1750 2658 1754 2662
rect 1766 2658 1770 2662
rect 1798 2658 1802 2662
rect 1806 2658 1810 2662
rect 1830 2658 1834 2662
rect 1862 2658 1866 2662
rect 1926 2659 1930 2663
rect 2022 2658 2026 2662
rect 2030 2658 2034 2662
rect 2046 2658 2050 2662
rect 2054 2658 2058 2662
rect 2094 2658 2098 2662
rect 2118 2658 2122 2662
rect 2158 2658 2162 2662
rect 2182 2658 2186 2662
rect 2222 2658 2226 2662
rect 2270 2658 2274 2662
rect 2286 2658 2290 2662
rect 2294 2658 2298 2662
rect 2422 2658 2426 2662
rect 2462 2658 2466 2662
rect 2518 2659 2522 2663
rect 2622 2658 2626 2662
rect 2646 2658 2650 2662
rect 2726 2658 2730 2662
rect 2782 2659 2786 2663
rect 2878 2658 2882 2662
rect 2902 2658 2906 2662
rect 2966 2658 2970 2662
rect 2990 2658 2994 2662
rect 2998 2658 3002 2662
rect 3062 2658 3066 2662
rect 3150 2658 3154 2662
rect 3158 2658 3162 2662
rect 3214 2658 3218 2662
rect 3254 2658 3258 2662
rect 3310 2658 3314 2662
rect 3318 2658 3322 2662
rect 3382 2658 3386 2662
rect 3430 2658 3434 2662
rect 3454 2658 3458 2662
rect 3486 2658 3490 2662
rect 3550 2658 3554 2662
rect 3606 2658 3610 2662
rect 3614 2658 3618 2662
rect 3654 2658 3658 2662
rect 3662 2658 3666 2662
rect 3718 2658 3722 2662
rect 3750 2658 3754 2662
rect 3790 2658 3794 2662
rect 3814 2658 3818 2662
rect 3822 2658 3826 2662
rect 3846 2658 3850 2662
rect 3878 2658 3882 2662
rect 3950 2658 3954 2662
rect 3998 2658 4002 2662
rect 4014 2658 4018 2662
rect 4102 2658 4106 2662
rect 4134 2659 4138 2663
rect 4174 2658 4178 2662
rect 4198 2658 4202 2662
rect 4206 2658 4210 2662
rect 4214 2658 4218 2662
rect 4222 2658 4226 2662
rect 4246 2658 4250 2662
rect 4262 2658 4266 2662
rect 4302 2658 4306 2662
rect 4326 2658 4330 2662
rect 4334 2658 4338 2662
rect 4342 2658 4346 2662
rect 4358 2658 4362 2662
rect 4398 2658 4402 2662
rect 4454 2658 4458 2662
rect 4470 2658 4474 2662
rect 4478 2658 4482 2662
rect 4502 2658 4506 2662
rect 4534 2658 4538 2662
rect 4550 2658 4554 2662
rect 4566 2658 4570 2662
rect 4622 2658 4626 2662
rect 4686 2658 4690 2662
rect 4710 2658 4714 2662
rect 4726 2658 4730 2662
rect 4750 2658 4754 2662
rect 4774 2658 4778 2662
rect 4830 2658 4834 2662
rect 4862 2658 4866 2662
rect 4878 2658 4882 2662
rect 4902 2658 4906 2662
rect 4910 2658 4914 2662
rect 4942 2658 4946 2662
rect 5038 2658 5042 2662
rect 5126 2658 5130 2662
rect 5150 2658 5154 2662
rect 5238 2658 5242 2662
rect 126 2648 130 2652
rect 134 2648 138 2652
rect 150 2648 154 2652
rect 446 2648 450 2652
rect 550 2648 554 2652
rect 734 2648 738 2652
rect 798 2648 802 2652
rect 902 2648 906 2652
rect 934 2648 938 2652
rect 1086 2648 1090 2652
rect 1142 2648 1146 2652
rect 1198 2648 1202 2652
rect 1326 2648 1330 2652
rect 1438 2648 1442 2652
rect 1678 2648 1682 2652
rect 1726 2648 1730 2652
rect 1750 2648 1754 2652
rect 1854 2648 1858 2652
rect 2078 2648 2082 2652
rect 2134 2648 2138 2652
rect 2158 2648 2162 2652
rect 2190 2648 2194 2652
rect 2238 2648 2242 2652
rect 2310 2648 2314 2652
rect 2702 2648 2706 2652
rect 2726 2648 2730 2652
rect 3542 2648 3546 2652
rect 3646 2648 3650 2652
rect 3830 2648 3834 2652
rect 3862 2648 3866 2652
rect 4062 2648 4066 2652
rect 4342 2648 4346 2652
rect 4414 2648 4418 2652
rect 4646 2648 4650 2652
rect 4830 2648 4834 2652
rect 4846 2648 4850 2652
rect 4926 2648 4930 2652
rect 278 2638 282 2642
rect 414 2638 418 2642
rect 542 2638 546 2642
rect 702 2638 706 2642
rect 766 2638 770 2642
rect 918 2638 922 2642
rect 1566 2638 1570 2642
rect 2942 2638 2946 2642
rect 4814 2638 4818 2642
rect 4310 2628 4314 2632
rect 830 2618 834 2622
rect 846 2618 850 2622
rect 950 2618 954 2622
rect 1662 2618 1666 2622
rect 1990 2618 1994 2622
rect 2094 2618 2098 2622
rect 2254 2618 2258 2622
rect 2918 2618 2922 2622
rect 2974 2618 2978 2622
rect 3174 2618 3178 2622
rect 3198 2618 3202 2622
rect 3398 2618 3402 2622
rect 3566 2618 3570 2622
rect 3630 2618 3634 2622
rect 3702 2618 3706 2622
rect 3766 2618 3770 2622
rect 3798 2618 3802 2622
rect 4230 2618 4234 2622
rect 4494 2618 4498 2622
rect 4790 2618 4794 2622
rect 4862 2618 4866 2622
rect 4886 2618 4890 2622
rect 5094 2618 5098 2622
rect 330 2603 334 2607
rect 337 2603 341 2607
rect 1354 2603 1358 2607
rect 1361 2603 1365 2607
rect 2386 2603 2390 2607
rect 2393 2603 2397 2607
rect 3402 2603 3406 2607
rect 3409 2603 3413 2607
rect 4426 2603 4430 2607
rect 4433 2603 4437 2607
rect 486 2588 490 2592
rect 1046 2588 1050 2592
rect 1086 2588 1090 2592
rect 1542 2588 1546 2592
rect 1758 2588 1762 2592
rect 2126 2588 2130 2592
rect 2238 2588 2242 2592
rect 2278 2588 2282 2592
rect 2822 2588 2826 2592
rect 3326 2588 3330 2592
rect 3470 2588 3474 2592
rect 3502 2588 3506 2592
rect 4038 2588 4042 2592
rect 4062 2588 4066 2592
rect 4102 2588 4106 2592
rect 4262 2588 4266 2592
rect 4510 2588 4514 2592
rect 4806 2588 4810 2592
rect 5166 2588 5170 2592
rect 5270 2588 5274 2592
rect 94 2578 98 2582
rect 3294 2578 3298 2582
rect 4350 2578 4354 2582
rect 4606 2578 4610 2582
rect 134 2568 138 2572
rect 254 2568 258 2572
rect 294 2568 298 2572
rect 350 2568 354 2572
rect 702 2568 706 2572
rect 798 2568 802 2572
rect 966 2568 970 2572
rect 1006 2568 1010 2572
rect 1294 2568 1298 2572
rect 1310 2568 1314 2572
rect 1582 2568 1586 2572
rect 1918 2568 1922 2572
rect 2294 2568 2298 2572
rect 4238 2568 4242 2572
rect 110 2558 114 2562
rect 126 2558 130 2562
rect 150 2558 154 2562
rect 270 2558 274 2562
rect 38 2548 42 2552
rect 62 2548 66 2552
rect 110 2548 114 2552
rect 150 2548 154 2552
rect 198 2548 202 2552
rect 270 2548 274 2552
rect 374 2558 378 2562
rect 470 2558 474 2562
rect 502 2558 506 2562
rect 814 2558 818 2562
rect 830 2558 834 2562
rect 982 2558 986 2562
rect 318 2548 322 2552
rect 382 2548 386 2552
rect 414 2548 418 2552
rect 454 2548 458 2552
rect 486 2548 490 2552
rect 534 2547 538 2551
rect 646 2548 650 2552
rect 766 2547 770 2551
rect 822 2548 826 2552
rect 830 2548 834 2552
rect 846 2548 850 2552
rect 910 2548 914 2552
rect 982 2548 986 2552
rect 1126 2558 1130 2562
rect 1158 2558 1162 2562
rect 1358 2558 1362 2562
rect 1374 2558 1378 2562
rect 1390 2558 1394 2562
rect 1526 2558 1530 2562
rect 1550 2558 1554 2562
rect 1614 2558 1618 2562
rect 1902 2558 1906 2562
rect 2070 2558 2074 2562
rect 2406 2558 2410 2562
rect 2430 2558 2434 2562
rect 2638 2558 2642 2562
rect 2798 2558 2802 2562
rect 3014 2558 3018 2562
rect 3038 2558 3042 2562
rect 3190 2558 3194 2562
rect 3214 2558 3218 2562
rect 3558 2558 3562 2562
rect 3750 2558 3754 2562
rect 4158 2558 4162 2562
rect 4182 2558 4186 2562
rect 4382 2558 4386 2562
rect 4398 2558 4402 2562
rect 1062 2548 1066 2552
rect 1070 2548 1074 2552
rect 1102 2548 1106 2552
rect 1134 2548 1138 2552
rect 1182 2548 1186 2552
rect 1190 2548 1194 2552
rect 1262 2548 1266 2552
rect 1326 2548 1330 2552
rect 1342 2548 1346 2552
rect 1422 2548 1426 2552
rect 1430 2548 1434 2552
rect 1454 2548 1458 2552
rect 1510 2548 1514 2552
rect 1526 2548 1530 2552
rect 1566 2548 1570 2552
rect 1582 2548 1586 2552
rect 1598 2548 1602 2552
rect 1622 2548 1626 2552
rect 1630 2548 1634 2552
rect 1654 2548 1658 2552
rect 1662 2548 1666 2552
rect 102 2538 106 2542
rect 158 2538 162 2542
rect 174 2538 178 2542
rect 214 2538 218 2542
rect 262 2538 266 2542
rect 326 2538 330 2542
rect 358 2538 362 2542
rect 374 2538 378 2542
rect 390 2538 394 2542
rect 438 2538 442 2542
rect 446 2538 450 2542
rect 478 2538 482 2542
rect 550 2538 554 2542
rect 750 2538 754 2542
rect 822 2538 826 2542
rect 854 2538 858 2542
rect 974 2538 978 2542
rect 1030 2538 1034 2542
rect 1694 2547 1698 2551
rect 1718 2548 1722 2552
rect 1766 2548 1770 2552
rect 1822 2548 1826 2552
rect 1926 2548 1930 2552
rect 1974 2547 1978 2551
rect 2006 2548 2010 2552
rect 2046 2548 2050 2552
rect 2110 2548 2114 2552
rect 2134 2548 2138 2552
rect 2214 2548 2218 2552
rect 2246 2548 2250 2552
rect 2286 2548 2290 2552
rect 2334 2548 2338 2552
rect 2494 2548 2498 2552
rect 2502 2548 2506 2552
rect 2550 2548 2554 2552
rect 2566 2548 2570 2552
rect 2574 2548 2578 2552
rect 2598 2548 2602 2552
rect 2622 2548 2626 2552
rect 2638 2548 2642 2552
rect 2670 2548 2674 2552
rect 2694 2548 2698 2552
rect 2726 2548 2730 2552
rect 2734 2548 2738 2552
rect 2758 2548 2762 2552
rect 2790 2548 2794 2552
rect 2838 2548 2842 2552
rect 2878 2548 2882 2552
rect 2902 2548 2906 2552
rect 2950 2548 2954 2552
rect 2982 2548 2986 2552
rect 2998 2548 3002 2552
rect 3014 2548 3018 2552
rect 3030 2548 3034 2552
rect 3046 2548 3050 2552
rect 3086 2548 3090 2552
rect 3134 2548 3138 2552
rect 3150 2548 3154 2552
rect 3166 2548 3170 2552
rect 3174 2548 3178 2552
rect 3246 2548 3250 2552
rect 3254 2548 3258 2552
rect 3310 2548 3314 2552
rect 3342 2548 3346 2552
rect 3374 2548 3378 2552
rect 3406 2548 3410 2552
rect 3486 2548 3490 2552
rect 3518 2548 3522 2552
rect 3582 2548 3586 2552
rect 3638 2548 3642 2552
rect 3678 2548 3682 2552
rect 3702 2548 3706 2552
rect 3734 2548 3738 2552
rect 3742 2548 3746 2552
rect 3774 2548 3778 2552
rect 3806 2548 3810 2552
rect 3870 2548 3874 2552
rect 3958 2548 3962 2552
rect 3982 2548 3986 2552
rect 4022 2548 4026 2552
rect 4078 2548 4082 2552
rect 4134 2548 4138 2552
rect 4166 2548 4170 2552
rect 4190 2548 4194 2552
rect 4198 2548 4202 2552
rect 4278 2548 4282 2552
rect 4310 2548 4314 2552
rect 4318 2548 4322 2552
rect 4430 2548 4434 2552
rect 4462 2548 4466 2552
rect 4486 2558 4490 2562
rect 4622 2558 4626 2562
rect 4902 2558 4906 2562
rect 5070 2558 5074 2562
rect 4550 2548 4554 2552
rect 4638 2548 4642 2552
rect 4710 2548 4714 2552
rect 4766 2548 4770 2552
rect 4798 2548 4802 2552
rect 4862 2548 4866 2552
rect 4910 2548 4914 2552
rect 4918 2548 4922 2552
rect 4990 2548 4994 2552
rect 5046 2548 5050 2552
rect 5134 2558 5138 2562
rect 5094 2548 5098 2552
rect 5126 2548 5130 2552
rect 5134 2548 5138 2552
rect 5158 2548 5162 2552
rect 5206 2548 5210 2552
rect 5222 2548 5226 2552
rect 5262 2548 5266 2552
rect 1094 2538 1098 2542
rect 1158 2538 1162 2542
rect 1182 2538 1186 2542
rect 1214 2538 1218 2542
rect 1230 2538 1234 2542
rect 1246 2538 1250 2542
rect 1278 2538 1282 2542
rect 1318 2538 1322 2542
rect 1334 2538 1338 2542
rect 1366 2538 1370 2542
rect 1398 2538 1402 2542
rect 1478 2538 1482 2542
rect 1534 2538 1538 2542
rect 1550 2538 1554 2542
rect 1558 2538 1562 2542
rect 1590 2538 1594 2542
rect 1830 2538 1834 2542
rect 1918 2538 1922 2542
rect 2046 2538 2050 2542
rect 2086 2538 2090 2542
rect 2206 2538 2210 2542
rect 2222 2538 2226 2542
rect 2358 2538 2362 2542
rect 2430 2538 2434 2542
rect 2446 2538 2450 2542
rect 2670 2538 2674 2542
rect 326 2528 330 2532
rect 406 2528 410 2532
rect 438 2528 442 2532
rect 630 2528 634 2532
rect 902 2528 906 2532
rect 1134 2528 1138 2532
rect 1150 2528 1154 2532
rect 1446 2528 1450 2532
rect 1486 2528 1490 2532
rect 1782 2528 1786 2532
rect 1942 2528 1946 2532
rect 1974 2528 1978 2532
rect 2102 2528 2106 2532
rect 2270 2528 2274 2532
rect 2478 2528 2482 2532
rect 2582 2528 2586 2532
rect 2694 2538 2698 2542
rect 2718 2538 2722 2542
rect 2766 2538 2770 2542
rect 2790 2538 2794 2542
rect 2846 2538 2850 2542
rect 2910 2538 2914 2542
rect 2942 2538 2946 2542
rect 2950 2538 2954 2542
rect 2974 2538 2978 2542
rect 2990 2538 2994 2542
rect 3022 2538 3026 2542
rect 3054 2538 3058 2542
rect 3078 2538 3082 2542
rect 3102 2538 3106 2542
rect 3118 2538 3122 2542
rect 3166 2538 3170 2542
rect 3198 2538 3202 2542
rect 3222 2538 3226 2542
rect 3390 2538 3394 2542
rect 3454 2538 3458 2542
rect 3574 2538 3578 2542
rect 3646 2538 3650 2542
rect 3750 2538 3754 2542
rect 3798 2538 3802 2542
rect 3878 2538 3882 2542
rect 4142 2538 4146 2542
rect 4166 2538 4170 2542
rect 4342 2538 4346 2542
rect 4398 2538 4402 2542
rect 4454 2538 4458 2542
rect 4478 2538 4482 2542
rect 4590 2538 4594 2542
rect 4646 2538 4650 2542
rect 4734 2538 4738 2542
rect 4790 2538 4794 2542
rect 4838 2538 4842 2542
rect 4886 2538 4890 2542
rect 4926 2538 4930 2542
rect 5006 2538 5010 2542
rect 5046 2538 5050 2542
rect 5102 2538 5106 2542
rect 5158 2538 5162 2542
rect 2750 2528 2754 2532
rect 2782 2528 2786 2532
rect 2806 2528 2810 2532
rect 2926 2528 2930 2532
rect 2958 2528 2962 2532
rect 3062 2528 3066 2532
rect 3118 2528 3122 2532
rect 3190 2528 3194 2532
rect 3598 2528 3602 2532
rect 3782 2528 3786 2532
rect 4118 2528 4122 2532
rect 4134 2528 4138 2532
rect 4238 2528 4242 2532
rect 4294 2528 4298 2532
rect 4334 2528 4338 2532
rect 4614 2528 4618 2532
rect 4750 2528 4754 2532
rect 4782 2528 4786 2532
rect 5110 2528 5114 2532
rect 5278 2528 5282 2532
rect 470 2518 474 2522
rect 598 2518 602 2522
rect 694 2518 698 2522
rect 1126 2518 1130 2522
rect 1438 2518 1442 2522
rect 1638 2518 1642 2522
rect 1774 2518 1778 2522
rect 1894 2518 1898 2522
rect 1934 2518 1938 2522
rect 2038 2518 2042 2522
rect 2094 2518 2098 2522
rect 2126 2518 2130 2522
rect 2406 2518 2410 2522
rect 2438 2518 2442 2522
rect 2742 2518 2746 2522
rect 2886 2518 2890 2522
rect 3070 2518 3074 2522
rect 3110 2518 3114 2522
rect 3134 2518 3138 2522
rect 3214 2518 3218 2522
rect 3270 2518 3274 2522
rect 3326 2518 3330 2522
rect 3358 2518 3362 2522
rect 3542 2518 3546 2522
rect 3558 2518 3562 2522
rect 3622 2518 3626 2522
rect 3686 2518 3690 2522
rect 3718 2518 3722 2522
rect 3814 2518 3818 2522
rect 3926 2518 3930 2522
rect 4062 2518 4066 2522
rect 4150 2518 4154 2522
rect 4206 2518 4210 2522
rect 4262 2518 4266 2522
rect 4326 2518 4330 2522
rect 4382 2518 4386 2522
rect 4622 2518 4626 2522
rect 4654 2518 4658 2522
rect 4942 2518 4946 2522
rect 5078 2518 5082 2522
rect 5118 2518 5122 2522
rect 850 2503 854 2507
rect 857 2503 861 2507
rect 1874 2503 1878 2507
rect 1881 2503 1885 2507
rect 2890 2503 2894 2507
rect 2897 2503 2901 2507
rect 3922 2503 3926 2507
rect 3929 2503 3933 2507
rect 4938 2503 4942 2507
rect 4945 2503 4949 2507
rect 94 2488 98 2492
rect 470 2488 474 2492
rect 494 2488 498 2492
rect 526 2488 530 2492
rect 646 2488 650 2492
rect 1174 2488 1178 2492
rect 1366 2488 1370 2492
rect 1406 2488 1410 2492
rect 1526 2488 1530 2492
rect 1558 2488 1562 2492
rect 1798 2488 1802 2492
rect 2014 2488 2018 2492
rect 2046 2488 2050 2492
rect 2094 2488 2098 2492
rect 2190 2488 2194 2492
rect 2254 2488 2258 2492
rect 2302 2488 2306 2492
rect 2342 2488 2346 2492
rect 2478 2488 2482 2492
rect 2654 2488 2658 2492
rect 2670 2488 2674 2492
rect 2878 2488 2882 2492
rect 2990 2488 2994 2492
rect 3030 2488 3034 2492
rect 3102 2488 3106 2492
rect 3262 2488 3266 2492
rect 3446 2488 3450 2492
rect 3766 2488 3770 2492
rect 3902 2488 3906 2492
rect 3990 2488 3994 2492
rect 4110 2488 4114 2492
rect 4142 2488 4146 2492
rect 4246 2488 4250 2492
rect 4342 2488 4346 2492
rect 4358 2488 4362 2492
rect 4510 2488 4514 2492
rect 4670 2488 4674 2492
rect 4838 2488 4842 2492
rect 4974 2488 4978 2492
rect 5086 2488 5090 2492
rect 5190 2488 5194 2492
rect 214 2478 218 2482
rect 398 2478 402 2482
rect 598 2478 602 2482
rect 606 2478 610 2482
rect 686 2478 690 2482
rect 702 2478 706 2482
rect 998 2478 1002 2482
rect 102 2468 106 2472
rect 150 2468 154 2472
rect 182 2468 186 2472
rect 286 2468 290 2472
rect 302 2468 306 2472
rect 350 2468 354 2472
rect 518 2468 522 2472
rect 558 2468 562 2472
rect 566 2468 570 2472
rect 614 2468 618 2472
rect 654 2468 658 2472
rect 1646 2478 1650 2482
rect 1774 2478 1778 2482
rect 1830 2478 1834 2482
rect 1918 2478 1922 2482
rect 1998 2478 2002 2482
rect 710 2468 714 2472
rect 742 2468 746 2472
rect 814 2468 818 2472
rect 846 2468 850 2472
rect 870 2468 874 2472
rect 910 2468 914 2472
rect 958 2468 962 2472
rect 966 2468 970 2472
rect 982 2468 986 2472
rect 1054 2468 1058 2472
rect 1094 2468 1098 2472
rect 1182 2468 1186 2472
rect 1214 2468 1218 2472
rect 38 2458 42 2462
rect 62 2458 66 2462
rect 110 2458 114 2462
rect 158 2458 162 2462
rect 174 2458 178 2462
rect 222 2458 226 2462
rect 294 2458 298 2462
rect 334 2458 338 2462
rect 1246 2468 1250 2472
rect 1286 2468 1290 2472
rect 1390 2468 1394 2472
rect 1414 2468 1418 2472
rect 1502 2468 1506 2472
rect 1622 2468 1626 2472
rect 1662 2468 1666 2472
rect 1758 2468 1762 2472
rect 1790 2468 1794 2472
rect 1862 2468 1866 2472
rect 1886 2468 1890 2472
rect 1982 2468 1986 2472
rect 2038 2478 2042 2482
rect 2078 2478 2082 2482
rect 2022 2468 2026 2472
rect 2558 2478 2562 2482
rect 2870 2478 2874 2482
rect 2926 2478 2930 2482
rect 3198 2478 3202 2482
rect 3246 2478 3250 2482
rect 3270 2478 3274 2482
rect 3358 2478 3362 2482
rect 3550 2478 3554 2482
rect 3654 2478 3658 2482
rect 3702 2478 3706 2482
rect 3830 2478 3834 2482
rect 4070 2478 4074 2482
rect 4118 2478 4122 2482
rect 4478 2478 4482 2482
rect 4638 2478 4642 2482
rect 4766 2478 4770 2482
rect 4782 2478 4786 2482
rect 5094 2478 5098 2482
rect 5270 2478 5274 2482
rect 2102 2468 2106 2472
rect 2118 2468 2122 2472
rect 2382 2468 2386 2472
rect 2430 2468 2434 2472
rect 2534 2468 2538 2472
rect 2574 2468 2578 2472
rect 2678 2468 2682 2472
rect 2686 2468 2690 2472
rect 2702 2468 2706 2472
rect 2718 2468 2722 2472
rect 2734 2468 2738 2472
rect 2750 2468 2754 2472
rect 2766 2468 2770 2472
rect 2798 2468 2802 2472
rect 2838 2468 2842 2472
rect 2854 2468 2858 2472
rect 2918 2468 2922 2472
rect 2950 2468 2954 2472
rect 2974 2468 2978 2472
rect 3014 2468 3018 2472
rect 3174 2468 3178 2472
rect 3190 2468 3194 2472
rect 3230 2468 3234 2472
rect 3294 2468 3298 2472
rect 3302 2468 3306 2472
rect 3326 2468 3330 2472
rect 3334 2468 3338 2472
rect 3366 2468 3370 2472
rect 3374 2468 3378 2472
rect 3406 2468 3410 2472
rect 3486 2468 3490 2472
rect 390 2458 394 2462
rect 422 2458 426 2462
rect 454 2458 458 2462
rect 478 2458 482 2462
rect 510 2458 514 2462
rect 542 2458 546 2462
rect 574 2458 578 2462
rect 614 2458 618 2462
rect 630 2458 634 2462
rect 662 2458 666 2462
rect 702 2458 706 2462
rect 718 2458 722 2462
rect 726 2458 730 2462
rect 742 2458 746 2462
rect 750 2458 754 2462
rect 758 2458 762 2462
rect 782 2458 786 2462
rect 822 2458 826 2462
rect 838 2458 842 2462
rect 870 2458 874 2462
rect 894 2458 898 2462
rect 926 2458 930 2462
rect 950 2458 954 2462
rect 974 2458 978 2462
rect 998 2458 1002 2462
rect 1014 2458 1018 2462
rect 1030 2458 1034 2462
rect 1062 2458 1066 2462
rect 1126 2458 1130 2462
rect 1142 2458 1146 2462
rect 1190 2458 1194 2462
rect 1222 2458 1226 2462
rect 1238 2458 1242 2462
rect 1254 2458 1258 2462
rect 1302 2459 1306 2463
rect 3518 2468 3522 2472
rect 3526 2468 3530 2472
rect 3574 2468 3578 2472
rect 3606 2468 3610 2472
rect 3694 2468 3698 2472
rect 3710 2468 3714 2472
rect 3742 2468 3746 2472
rect 3750 2468 3754 2472
rect 3806 2468 3810 2472
rect 3838 2468 3842 2472
rect 3894 2468 3898 2472
rect 3926 2468 3930 2472
rect 4046 2468 4050 2472
rect 4062 2468 4066 2472
rect 4094 2468 4098 2472
rect 4198 2468 4202 2472
rect 4254 2468 4258 2472
rect 4286 2468 4290 2472
rect 4294 2468 4298 2472
rect 4318 2468 4322 2472
rect 4326 2468 4330 2472
rect 4350 2468 4354 2472
rect 4382 2468 4386 2472
rect 4414 2468 4418 2472
rect 4454 2466 4458 2470
rect 4462 2468 4466 2472
rect 4470 2468 4474 2472
rect 4502 2468 4506 2472
rect 4590 2468 4594 2472
rect 4678 2468 4682 2472
rect 4694 2468 4698 2472
rect 4710 2468 4714 2472
rect 4790 2468 4794 2472
rect 4822 2468 4826 2472
rect 4894 2468 4898 2472
rect 4910 2468 4914 2472
rect 4926 2468 4930 2472
rect 4934 2468 4938 2472
rect 5054 2468 5058 2472
rect 5078 2468 5082 2472
rect 5206 2468 5210 2472
rect 1430 2458 1434 2462
rect 1438 2458 1442 2462
rect 1470 2458 1474 2462
rect 1510 2458 1514 2462
rect 1542 2458 1546 2462
rect 1582 2458 1586 2462
rect 1606 2458 1610 2462
rect 1614 2458 1618 2462
rect 1630 2458 1634 2462
rect 1686 2458 1690 2462
rect 1750 2458 1754 2462
rect 1782 2458 1786 2462
rect 1814 2458 1818 2462
rect 1854 2458 1858 2462
rect 1894 2458 1898 2462
rect 1934 2458 1938 2462
rect 1942 2458 1946 2462
rect 2030 2458 2034 2462
rect 2054 2458 2058 2462
rect 2062 2458 2066 2462
rect 2110 2458 2114 2462
rect 2126 2458 2130 2462
rect 2142 2458 2146 2462
rect 2166 2458 2170 2462
rect 2214 2458 2218 2462
rect 2238 2458 2242 2462
rect 2270 2458 2274 2462
rect 2278 2458 2282 2462
rect 2286 2458 2290 2462
rect 2318 2458 2322 2462
rect 2326 2458 2330 2462
rect 2374 2458 2378 2462
rect 2414 2458 2418 2462
rect 2422 2458 2426 2462
rect 2462 2458 2466 2462
rect 2542 2458 2546 2462
rect 2598 2458 2602 2462
rect 2694 2458 2698 2462
rect 2710 2458 2714 2462
rect 2726 2458 2730 2462
rect 2758 2458 2762 2462
rect 2774 2458 2778 2462
rect 2790 2458 2794 2462
rect 2846 2458 2850 2462
rect 2862 2458 2866 2462
rect 2894 2458 2898 2462
rect 2942 2458 2946 2462
rect 2950 2458 2954 2462
rect 2982 2458 2986 2462
rect 3006 2458 3010 2462
rect 3054 2458 3058 2462
rect 3078 2458 3082 2462
rect 3118 2458 3122 2462
rect 3126 2458 3130 2462
rect 3150 2458 3154 2462
rect 3190 2458 3194 2462
rect 3222 2458 3226 2462
rect 3230 2458 3234 2462
rect 3254 2458 3258 2462
rect 3318 2458 3322 2462
rect 3342 2458 3346 2462
rect 3358 2458 3362 2462
rect 3382 2458 3386 2462
rect 3446 2458 3450 2462
rect 3478 2458 3482 2462
rect 3494 2458 3498 2462
rect 3510 2458 3514 2462
rect 3518 2458 3522 2462
rect 3598 2458 3602 2462
rect 3630 2458 3634 2462
rect 3678 2458 3682 2462
rect 3734 2458 3738 2462
rect 3782 2458 3786 2462
rect 3886 2458 3890 2462
rect 3918 2458 3922 2462
rect 3982 2458 3986 2462
rect 4006 2458 4010 2462
rect 4038 2458 4042 2462
rect 4094 2458 4098 2462
rect 4102 2458 4106 2462
rect 4126 2458 4130 2462
rect 4206 2458 4210 2462
rect 4254 2458 4258 2462
rect 4278 2458 4282 2462
rect 4310 2458 4314 2462
rect 4358 2458 4362 2462
rect 4406 2458 4410 2462
rect 4438 2458 4442 2462
rect 4478 2458 4482 2462
rect 4494 2458 4498 2462
rect 4566 2458 4570 2462
rect 4622 2458 4626 2462
rect 4654 2458 4658 2462
rect 4686 2458 4690 2462
rect 4702 2458 4706 2462
rect 4718 2458 4722 2462
rect 4750 2458 4754 2462
rect 4766 2458 4770 2462
rect 4790 2458 4794 2462
rect 4814 2458 4818 2462
rect 4926 2458 4930 2462
rect 4934 2458 4938 2462
rect 5038 2459 5042 2463
rect 5070 2458 5074 2462
rect 5134 2458 5138 2462
rect 5150 2458 5154 2462
rect 5222 2459 5226 2463
rect 110 2448 114 2452
rect 126 2448 130 2452
rect 134 2448 138 2452
rect 150 2448 154 2452
rect 318 2448 322 2452
rect 438 2448 442 2452
rect 470 2448 474 2452
rect 646 2448 650 2452
rect 662 2448 666 2452
rect 678 2448 682 2452
rect 798 2448 802 2452
rect 894 2448 898 2452
rect 934 2448 938 2452
rect 990 2448 994 2452
rect 1022 2448 1026 2452
rect 1078 2448 1082 2452
rect 1206 2448 1210 2452
rect 1254 2448 1258 2452
rect 1270 2448 1274 2452
rect 1350 2448 1354 2452
rect 1406 2448 1410 2452
rect 1462 2448 1466 2452
rect 1646 2448 1650 2452
rect 1838 2448 1842 2452
rect 1910 2448 1914 2452
rect 1966 2448 1970 2452
rect 2142 2448 2146 2452
rect 2174 2448 2178 2452
rect 2358 2448 2362 2452
rect 2406 2448 2410 2452
rect 2662 2448 2666 2452
rect 2878 2448 2882 2452
rect 2958 2448 2962 2452
rect 2990 2448 2994 2452
rect 3166 2448 3170 2452
rect 3302 2448 3306 2452
rect 3398 2448 3402 2452
rect 3462 2448 3466 2452
rect 3494 2448 3498 2452
rect 3550 2448 3554 2452
rect 3582 2448 3586 2452
rect 3614 2448 3618 2452
rect 3662 2448 3666 2452
rect 3694 2448 3698 2452
rect 3718 2448 3722 2452
rect 3766 2448 3770 2452
rect 3862 2448 3866 2452
rect 3870 2448 3874 2452
rect 3886 2448 3890 2452
rect 3902 2448 3906 2452
rect 4062 2448 4066 2452
rect 4294 2448 4298 2452
rect 4390 2448 4394 2452
rect 4606 2448 4610 2452
rect 4622 2448 4626 2452
rect 4734 2448 4738 2452
rect 4798 2448 4802 2452
rect 4902 2448 4906 2452
rect 5174 2448 5178 2452
rect 590 2438 594 2442
rect 1038 2438 1042 2442
rect 1062 2438 1066 2442
rect 1238 2438 1242 2442
rect 1478 2438 1482 2442
rect 2158 2438 2162 2442
rect 4342 2438 4346 2442
rect 774 2428 778 2432
rect 950 2428 954 2432
rect 2374 2428 2378 2432
rect 2550 2428 2554 2432
rect 2734 2428 2738 2432
rect 2830 2428 2834 2432
rect 4070 2428 4074 2432
rect 142 2418 146 2422
rect 278 2418 282 2422
rect 574 2418 578 2422
rect 1030 2418 1034 2422
rect 1190 2418 1194 2422
rect 1526 2418 1530 2422
rect 1598 2418 1602 2422
rect 1742 2418 1746 2422
rect 1774 2418 1778 2422
rect 1854 2418 1858 2422
rect 1894 2418 1898 2422
rect 2166 2418 2170 2422
rect 2190 2418 2194 2422
rect 2222 2418 2226 2422
rect 2446 2418 2450 2422
rect 2790 2418 2794 2422
rect 2934 2418 2938 2422
rect 3070 2418 3074 2422
rect 3142 2418 3146 2422
rect 3198 2418 3202 2422
rect 3238 2418 3242 2422
rect 3286 2418 3290 2422
rect 3630 2418 3634 2422
rect 3678 2418 3682 2422
rect 3734 2418 3738 2422
rect 3846 2418 3850 2422
rect 3958 2418 3962 2422
rect 3990 2418 3994 2422
rect 4022 2418 4026 2422
rect 4262 2418 4266 2422
rect 5286 2418 5290 2422
rect 330 2403 334 2407
rect 337 2403 341 2407
rect 1354 2403 1358 2407
rect 1361 2403 1365 2407
rect 2386 2403 2390 2407
rect 2393 2403 2397 2407
rect 3402 2403 3406 2407
rect 3409 2403 3413 2407
rect 4426 2403 4430 2407
rect 4433 2403 4437 2407
rect 638 2388 642 2392
rect 654 2388 658 2392
rect 742 2388 746 2392
rect 886 2388 890 2392
rect 1310 2388 1314 2392
rect 1382 2388 1386 2392
rect 1454 2388 1458 2392
rect 1486 2388 1490 2392
rect 1510 2388 1514 2392
rect 1686 2388 1690 2392
rect 1710 2388 1714 2392
rect 1806 2388 1810 2392
rect 2022 2388 2026 2392
rect 2118 2388 2122 2392
rect 2166 2388 2170 2392
rect 2310 2388 2314 2392
rect 2462 2388 2466 2392
rect 2486 2388 2490 2392
rect 2534 2388 2538 2392
rect 2558 2388 2562 2392
rect 2622 2388 2626 2392
rect 2662 2388 2666 2392
rect 2750 2388 2754 2392
rect 2782 2388 2786 2392
rect 2982 2388 2986 2392
rect 3686 2388 3690 2392
rect 3766 2388 3770 2392
rect 4054 2388 4058 2392
rect 4110 2388 4114 2392
rect 4134 2388 4138 2392
rect 4166 2388 4170 2392
rect 4462 2388 4466 2392
rect 4542 2388 4546 2392
rect 5118 2388 5122 2392
rect 5222 2388 5226 2392
rect 4294 2378 4298 2382
rect 510 2368 514 2372
rect 622 2368 626 2372
rect 942 2368 946 2372
rect 966 2368 970 2372
rect 1118 2368 1122 2372
rect 2422 2368 2426 2372
rect 2630 2368 2634 2372
rect 4190 2368 4194 2372
rect 5110 2368 5114 2372
rect 5278 2368 5282 2372
rect 142 2358 146 2362
rect 542 2358 546 2362
rect 670 2358 674 2362
rect 678 2358 682 2362
rect 758 2358 762 2362
rect 38 2348 42 2352
rect 62 2348 66 2352
rect 126 2348 130 2352
rect 142 2348 146 2352
rect 150 2348 154 2352
rect 158 2348 162 2352
rect 182 2348 186 2352
rect 118 2338 122 2342
rect 222 2347 226 2351
rect 318 2348 322 2352
rect 390 2348 394 2352
rect 454 2348 458 2352
rect 462 2348 466 2352
rect 510 2348 514 2352
rect 526 2348 530 2352
rect 574 2347 578 2351
rect 654 2348 658 2352
rect 718 2348 722 2352
rect 742 2348 746 2352
rect 766 2348 770 2352
rect 830 2348 834 2352
rect 926 2348 930 2352
rect 942 2348 946 2352
rect 1022 2358 1026 2362
rect 1134 2358 1138 2362
rect 1150 2358 1154 2362
rect 1166 2358 1170 2362
rect 1182 2358 1186 2362
rect 1214 2358 1218 2362
rect 1502 2358 1506 2362
rect 1606 2358 1610 2362
rect 1742 2358 1746 2362
rect 1774 2358 1778 2362
rect 1886 2358 1890 2362
rect 1934 2358 1938 2362
rect 982 2348 986 2352
rect 1006 2348 1010 2352
rect 1062 2348 1066 2352
rect 1134 2348 1138 2352
rect 1166 2348 1170 2352
rect 1190 2348 1194 2352
rect 1214 2348 1218 2352
rect 1254 2348 1258 2352
rect 1318 2348 1322 2352
rect 1382 2348 1386 2352
rect 1422 2348 1426 2352
rect 1430 2348 1434 2352
rect 1438 2348 1442 2352
rect 1462 2348 1466 2352
rect 1550 2348 1554 2352
rect 1558 2348 1562 2352
rect 1590 2348 1594 2352
rect 1598 2348 1602 2352
rect 1622 2348 1626 2352
rect 1638 2348 1642 2352
rect 1670 2348 1674 2352
rect 1678 2348 1682 2352
rect 1718 2348 1722 2352
rect 1750 2348 1754 2352
rect 1766 2348 1770 2352
rect 1790 2348 1794 2352
rect 1798 2348 1802 2352
rect 1830 2348 1834 2352
rect 1838 2348 1842 2352
rect 1878 2348 1882 2352
rect 1982 2347 1986 2351
rect 2022 2348 2026 2352
rect 2046 2358 2050 2362
rect 2110 2358 2114 2362
rect 2158 2358 2162 2362
rect 2646 2358 2650 2362
rect 2702 2358 2706 2362
rect 2766 2358 2770 2362
rect 2862 2358 2866 2362
rect 2950 2358 2954 2362
rect 3126 2358 3130 2362
rect 3334 2358 3338 2362
rect 3358 2358 3362 2362
rect 3390 2358 3394 2362
rect 3406 2358 3410 2362
rect 3726 2358 3730 2362
rect 2062 2348 2066 2352
rect 2126 2348 2130 2352
rect 2190 2348 2194 2352
rect 2222 2348 2226 2352
rect 2238 2348 2242 2352
rect 2254 2348 2258 2352
rect 2262 2348 2266 2352
rect 2294 2348 2298 2352
rect 2326 2348 2330 2352
rect 2334 2348 2338 2352
rect 2342 2348 2346 2352
rect 2366 2348 2370 2352
rect 2406 2348 2410 2352
rect 2430 2348 2434 2352
rect 2438 2348 2442 2352
rect 2446 2348 2450 2352
rect 2502 2348 2506 2352
rect 2510 2348 2514 2352
rect 2542 2348 2546 2352
rect 2550 2348 2554 2352
rect 2566 2348 2570 2352
rect 2606 2348 2610 2352
rect 2614 2348 2618 2352
rect 2638 2348 2642 2352
rect 2654 2348 2658 2352
rect 2686 2348 2690 2352
rect 2734 2348 2738 2352
rect 2750 2348 2754 2352
rect 2774 2348 2778 2352
rect 2798 2348 2802 2352
rect 2830 2348 2834 2352
rect 2846 2348 2850 2352
rect 2862 2348 2866 2352
rect 2886 2348 2890 2352
rect 2910 2348 2914 2352
rect 2934 2348 2938 2352
rect 2966 2348 2970 2352
rect 2990 2348 2994 2352
rect 2998 2348 3002 2352
rect 3030 2348 3034 2352
rect 3062 2348 3066 2352
rect 3094 2348 3098 2352
rect 3110 2348 3114 2352
rect 3158 2348 3162 2352
rect 3174 2348 3178 2352
rect 3206 2348 3210 2352
rect 3214 2348 3218 2352
rect 3246 2348 3250 2352
rect 3278 2348 3282 2352
rect 3286 2348 3290 2352
rect 3294 2348 3298 2352
rect 3318 2348 3322 2352
rect 3366 2348 3370 2352
rect 3374 2348 3378 2352
rect 3438 2348 3442 2352
rect 3486 2348 3490 2352
rect 238 2338 242 2342
rect 310 2338 314 2342
rect 350 2338 354 2342
rect 438 2338 442 2342
rect 470 2338 474 2342
rect 518 2338 522 2342
rect 542 2338 546 2342
rect 646 2338 650 2342
rect 694 2338 698 2342
rect 726 2338 730 2342
rect 734 2338 738 2342
rect 806 2338 810 2342
rect 854 2338 858 2342
rect 934 2338 938 2342
rect 990 2338 994 2342
rect 998 2338 1002 2342
rect 1014 2338 1018 2342
rect 1038 2338 1042 2342
rect 1126 2338 1130 2342
rect 1158 2338 1162 2342
rect 1190 2338 1194 2342
rect 1230 2338 1234 2342
rect 1326 2338 1330 2342
rect 1390 2338 1394 2342
rect 1478 2338 1482 2342
rect 1518 2338 1522 2342
rect 1614 2338 1618 2342
rect 1630 2338 1634 2342
rect 1646 2338 1650 2342
rect 1662 2338 1666 2342
rect 1838 2338 1842 2342
rect 1910 2338 1914 2342
rect 1974 2338 1978 2342
rect 2014 2338 2018 2342
rect 2070 2338 2074 2342
rect 2078 2338 2082 2342
rect 2126 2338 2130 2342
rect 2134 2338 2138 2342
rect 2182 2338 2186 2342
rect 2198 2338 2202 2342
rect 2246 2338 2250 2342
rect 2270 2338 2274 2342
rect 2286 2338 2290 2342
rect 2518 2338 2522 2342
rect 2534 2338 2538 2342
rect 2678 2338 2682 2342
rect 2726 2338 2730 2342
rect 2742 2338 2746 2342
rect 2806 2338 2810 2342
rect 2822 2338 2826 2342
rect 2838 2338 2842 2342
rect 2870 2338 2874 2342
rect 2894 2338 2898 2342
rect 2926 2338 2930 2342
rect 2990 2338 2994 2342
rect 3006 2338 3010 2342
rect 3022 2338 3026 2342
rect 3062 2338 3066 2342
rect 3086 2338 3090 2342
rect 3094 2338 3098 2342
rect 3134 2338 3138 2342
rect 3166 2338 3170 2342
rect 3182 2338 3186 2342
rect 3198 2338 3202 2342
rect 3222 2338 3226 2342
rect 3270 2338 3274 2342
rect 3326 2338 3330 2342
rect 3334 2338 3338 2342
rect 3350 2338 3354 2342
rect 3382 2338 3386 2342
rect 3422 2338 3426 2342
rect 3430 2338 3434 2342
rect 3446 2338 3450 2342
rect 3478 2338 3482 2342
rect 3494 2338 3498 2342
rect 3510 2348 3514 2352
rect 3542 2348 3546 2352
rect 3574 2348 3578 2352
rect 3590 2348 3594 2352
rect 3614 2348 3618 2352
rect 3622 2348 3626 2352
rect 3630 2348 3634 2352
rect 3646 2348 3650 2352
rect 3662 2348 3666 2352
rect 3694 2348 3698 2352
rect 3742 2348 3746 2352
rect 3766 2348 3770 2352
rect 3790 2358 3794 2362
rect 3846 2358 3850 2362
rect 4094 2358 4098 2362
rect 4102 2358 4106 2362
rect 3806 2348 3810 2352
rect 3814 2348 3818 2352
rect 3830 2348 3834 2352
rect 3838 2348 3842 2352
rect 3846 2348 3850 2352
rect 3878 2348 3882 2352
rect 3894 2348 3898 2352
rect 3910 2348 3914 2352
rect 3950 2348 3954 2352
rect 3982 2348 3986 2352
rect 3990 2348 3994 2352
rect 4038 2348 4042 2352
rect 4078 2348 4082 2352
rect 4150 2348 4154 2352
rect 4182 2348 4186 2352
rect 4222 2348 4226 2352
rect 3518 2338 3522 2342
rect 3638 2338 3642 2342
rect 3670 2338 3674 2342
rect 3686 2338 3690 2342
rect 3750 2338 3754 2342
rect 3758 2338 3762 2342
rect 3814 2338 3818 2342
rect 4254 2347 4258 2351
rect 4294 2348 4298 2352
rect 4318 2358 4322 2362
rect 4398 2358 4402 2362
rect 4510 2358 4514 2362
rect 4638 2358 4642 2362
rect 4814 2358 4818 2362
rect 5238 2358 5242 2362
rect 5270 2358 5274 2362
rect 4334 2348 4338 2352
rect 4374 2348 4378 2352
rect 4406 2348 4410 2352
rect 4478 2348 4482 2352
rect 4486 2348 4490 2352
rect 4534 2348 4538 2352
rect 4574 2348 4578 2352
rect 4582 2348 4586 2352
rect 4662 2348 4666 2352
rect 4710 2348 4714 2352
rect 4758 2348 4762 2352
rect 4822 2348 4826 2352
rect 4830 2348 4834 2352
rect 4886 2348 4890 2352
rect 4902 2348 4906 2352
rect 4958 2348 4962 2352
rect 4966 2348 4970 2352
rect 4990 2348 4994 2352
rect 4998 2348 5002 2352
rect 3870 2338 3874 2342
rect 3902 2338 3906 2342
rect 3958 2338 3962 2342
rect 3974 2338 3978 2342
rect 3998 2338 4002 2342
rect 4078 2338 4082 2342
rect 4118 2338 4122 2342
rect 4286 2338 4290 2342
rect 4342 2338 4346 2342
rect 4382 2338 4386 2342
rect 4454 2338 4458 2342
rect 4526 2338 4530 2342
rect 4598 2338 4602 2342
rect 4654 2338 4658 2342
rect 4702 2338 4706 2342
rect 4750 2338 4754 2342
rect 4782 2338 4786 2342
rect 4838 2338 4842 2342
rect 4926 2338 4930 2342
rect 4990 2338 4994 2342
rect 5046 2347 5050 2351
rect 5150 2348 5154 2352
rect 5158 2348 5162 2352
rect 5222 2348 5226 2352
rect 5254 2348 5258 2352
rect 5262 2348 5266 2352
rect 5278 2348 5282 2352
rect 5294 2348 5298 2352
rect 5030 2338 5034 2342
rect 5126 2338 5130 2342
rect 5174 2338 5178 2342
rect 5214 2338 5218 2342
rect 5246 2338 5250 2342
rect 5302 2338 5306 2342
rect 166 2328 170 2332
rect 294 2328 298 2332
rect 486 2328 490 2332
rect 574 2328 578 2332
rect 782 2328 786 2332
rect 910 2328 914 2332
rect 1342 2328 1346 2332
rect 1582 2328 1586 2332
rect 1694 2328 1698 2332
rect 1702 2328 1706 2332
rect 1750 2328 1754 2332
rect 1766 2328 1770 2332
rect 2166 2328 2170 2332
rect 2230 2328 2234 2332
rect 2286 2328 2290 2332
rect 2566 2328 2570 2332
rect 2598 2328 2602 2332
rect 2670 2328 2674 2332
rect 2790 2328 2794 2332
rect 2814 2328 2818 2332
rect 3022 2328 3026 2332
rect 3054 2328 3058 2332
rect 3086 2328 3090 2332
rect 3158 2328 3162 2332
rect 3190 2328 3194 2332
rect 3238 2328 3242 2332
rect 3270 2328 3274 2332
rect 3462 2328 3466 2332
rect 3550 2328 3554 2332
rect 3654 2328 3658 2332
rect 3686 2328 3690 2332
rect 3710 2328 3714 2332
rect 3854 2328 3858 2332
rect 3886 2328 3890 2332
rect 3934 2328 3938 2332
rect 4022 2328 4026 2332
rect 4502 2328 4506 2332
rect 4678 2328 4682 2332
rect 4686 2328 4690 2332
rect 5014 2328 5018 2332
rect 286 2318 290 2322
rect 302 2318 306 2322
rect 446 2318 450 2322
rect 702 2318 706 2322
rect 918 2318 922 2322
rect 1406 2318 1410 2322
rect 1534 2318 1538 2322
rect 1662 2318 1666 2322
rect 1742 2318 1746 2322
rect 2102 2318 2106 2322
rect 2158 2318 2162 2322
rect 2358 2318 2362 2322
rect 2718 2318 2722 2322
rect 2862 2318 2866 2322
rect 3014 2318 3018 2322
rect 3046 2318 3050 2322
rect 3518 2318 3522 2322
rect 4006 2318 4010 2322
rect 4054 2318 4058 2322
rect 4094 2318 4098 2322
rect 4102 2318 4106 2322
rect 4134 2318 4138 2322
rect 4358 2318 4362 2322
rect 4390 2318 4394 2322
rect 4462 2318 4466 2322
rect 4638 2318 4642 2322
rect 4670 2318 4674 2322
rect 4694 2318 4698 2322
rect 4718 2318 4722 2322
rect 4846 2318 4850 2322
rect 850 2303 854 2307
rect 857 2303 861 2307
rect 1874 2303 1878 2307
rect 1881 2303 1885 2307
rect 2890 2303 2894 2307
rect 2897 2303 2901 2307
rect 3922 2303 3926 2307
rect 3929 2303 3933 2307
rect 4938 2303 4942 2307
rect 4945 2303 4949 2307
rect 198 2288 202 2292
rect 246 2288 250 2292
rect 270 2288 274 2292
rect 398 2288 402 2292
rect 558 2288 562 2292
rect 1198 2288 1202 2292
rect 1382 2288 1386 2292
rect 1470 2288 1474 2292
rect 1734 2288 1738 2292
rect 1934 2288 1938 2292
rect 1958 2288 1962 2292
rect 2118 2288 2122 2292
rect 2142 2288 2146 2292
rect 2174 2288 2178 2292
rect 2230 2288 2234 2292
rect 2334 2288 2338 2292
rect 2486 2288 2490 2292
rect 2622 2288 2626 2292
rect 2646 2288 2650 2292
rect 2702 2288 2706 2292
rect 2726 2288 2730 2292
rect 2806 2288 2810 2292
rect 2846 2288 2850 2292
rect 2894 2288 2898 2292
rect 2918 2288 2922 2292
rect 2942 2288 2946 2292
rect 2974 2288 2978 2292
rect 3070 2288 3074 2292
rect 3262 2288 3266 2292
rect 3286 2288 3290 2292
rect 3310 2288 3314 2292
rect 3414 2288 3418 2292
rect 3454 2288 3458 2292
rect 3486 2288 3490 2292
rect 3598 2288 3602 2292
rect 3750 2288 3754 2292
rect 3766 2288 3770 2292
rect 3782 2288 3786 2292
rect 4222 2288 4226 2292
rect 4254 2288 4258 2292
rect 4510 2288 4514 2292
rect 4766 2288 4770 2292
rect 4838 2288 4842 2292
rect 4862 2288 4866 2292
rect 5142 2288 5146 2292
rect 5254 2288 5258 2292
rect 182 2278 186 2282
rect 126 2268 130 2272
rect 278 2278 282 2282
rect 406 2278 410 2282
rect 462 2278 466 2282
rect 838 2278 842 2282
rect 886 2278 890 2282
rect 1286 2278 1290 2282
rect 1294 2278 1298 2282
rect 1334 2278 1338 2282
rect 1390 2278 1394 2282
rect 1478 2278 1482 2282
rect 1486 2278 1490 2282
rect 1502 2278 1506 2282
rect 1534 2278 1538 2282
rect 1862 2278 1866 2282
rect 1918 2278 1922 2282
rect 1926 2278 1930 2282
rect 1966 2278 1970 2282
rect 1974 2278 1978 2282
rect 1990 2278 1994 2282
rect 206 2268 210 2272
rect 222 2268 226 2272
rect 262 2268 266 2272
rect 286 2268 290 2272
rect 302 2268 306 2272
rect 390 2268 394 2272
rect 422 2268 426 2272
rect 574 2268 578 2272
rect 726 2268 730 2272
rect 758 2268 762 2272
rect 38 2258 42 2262
rect 62 2258 66 2262
rect 118 2258 122 2262
rect 126 2258 130 2262
rect 150 2258 154 2262
rect 158 2258 162 2262
rect 166 2258 170 2262
rect 214 2258 218 2262
rect 230 2258 234 2262
rect 254 2258 258 2262
rect 286 2258 290 2262
rect 310 2258 314 2262
rect 366 2258 370 2262
rect 374 2258 378 2262
rect 382 2258 386 2262
rect 414 2258 418 2262
rect 446 2258 450 2262
rect 494 2259 498 2263
rect 798 2268 802 2272
rect 814 2268 818 2272
rect 1006 2268 1010 2272
rect 1062 2268 1066 2272
rect 1078 2268 1082 2272
rect 1102 2268 1106 2272
rect 1118 2268 1122 2272
rect 1142 2268 1146 2272
rect 1206 2268 1210 2272
rect 1262 2268 1266 2272
rect 1350 2268 1354 2272
rect 1398 2268 1402 2272
rect 1430 2268 1434 2272
rect 1446 2268 1450 2272
rect 1462 2268 1466 2272
rect 1502 2268 1506 2272
rect 1566 2268 1570 2272
rect 1654 2268 1658 2272
rect 1670 2268 1674 2272
rect 1702 2268 1706 2272
rect 1758 2268 1762 2272
rect 1774 2268 1778 2272
rect 1918 2268 1922 2272
rect 1998 2268 2002 2272
rect 2022 2268 2026 2272
rect 2038 2268 2042 2272
rect 2166 2268 2170 2272
rect 2278 2278 2282 2282
rect 2494 2278 2498 2282
rect 2614 2278 2618 2282
rect 2654 2278 2658 2282
rect 2854 2278 2858 2282
rect 3446 2278 3450 2282
rect 3478 2278 3482 2282
rect 3758 2278 3762 2282
rect 3934 2278 3938 2282
rect 4022 2278 4026 2282
rect 4070 2278 4074 2282
rect 4230 2278 4234 2282
rect 4350 2278 4354 2282
rect 2262 2268 2266 2272
rect 2286 2268 2290 2272
rect 2358 2268 2362 2272
rect 2374 2268 2378 2272
rect 2438 2268 2442 2272
rect 2478 2268 2482 2272
rect 2494 2268 2498 2272
rect 2534 2268 2538 2272
rect 2606 2268 2610 2272
rect 2694 2268 2698 2272
rect 2710 2268 2714 2272
rect 2750 2268 2754 2272
rect 2822 2268 2826 2272
rect 2838 2268 2842 2272
rect 2862 2268 2866 2272
rect 2958 2268 2962 2272
rect 3118 2268 3122 2272
rect 3150 2268 3154 2272
rect 3238 2268 3242 2272
rect 3318 2268 3322 2272
rect 3326 2268 3330 2272
rect 526 2258 530 2262
rect 598 2258 602 2262
rect 662 2258 666 2262
rect 678 2258 682 2262
rect 686 2258 690 2262
rect 710 2258 714 2262
rect 718 2258 722 2262
rect 734 2258 738 2262
rect 766 2258 770 2262
rect 782 2258 786 2262
rect 790 2258 794 2262
rect 822 2258 826 2262
rect 886 2259 890 2263
rect 966 2258 970 2262
rect 990 2258 994 2262
rect 998 2258 1002 2262
rect 1014 2258 1018 2262
rect 1038 2258 1042 2262
rect 1046 2258 1050 2262
rect 1054 2258 1058 2262
rect 1086 2258 1090 2262
rect 1134 2259 1138 2263
rect 1214 2258 1218 2262
rect 1254 2258 1258 2262
rect 1270 2258 1274 2262
rect 1294 2258 1298 2262
rect 1310 2258 1314 2262
rect 1318 2258 1322 2262
rect 1366 2258 1370 2262
rect 1406 2258 1410 2262
rect 1454 2258 1458 2262
rect 1486 2258 1490 2262
rect 1518 2258 1522 2262
rect 1558 2258 1562 2262
rect 1630 2258 1634 2262
rect 1678 2258 1682 2262
rect 1694 2258 1698 2262
rect 1750 2258 1754 2262
rect 1790 2259 1794 2263
rect 1822 2258 1826 2262
rect 1894 2258 1898 2262
rect 1910 2258 1914 2262
rect 1942 2258 1946 2262
rect 1950 2258 1954 2262
rect 1990 2258 1994 2262
rect 1998 2258 2002 2262
rect 2054 2259 2058 2263
rect 2126 2258 2130 2262
rect 2150 2258 2154 2262
rect 2214 2258 2218 2262
rect 2246 2258 2250 2262
rect 2254 2258 2258 2262
rect 2294 2258 2298 2262
rect 2318 2258 2322 2262
rect 2350 2258 2354 2262
rect 2382 2258 2386 2262
rect 2430 2258 2434 2262
rect 2462 2258 2466 2262
rect 2470 2258 2474 2262
rect 2510 2258 2514 2262
rect 2526 2258 2530 2262
rect 2566 2258 2570 2262
rect 2582 2258 2586 2262
rect 2630 2258 2634 2262
rect 2662 2258 2666 2262
rect 2686 2258 2690 2262
rect 2718 2258 2722 2262
rect 2726 2258 2730 2262
rect 2742 2258 2746 2262
rect 2758 2258 2762 2262
rect 2766 2258 2770 2262
rect 2790 2258 2794 2262
rect 310 2248 314 2252
rect 438 2248 442 2252
rect 782 2248 786 2252
rect 1238 2248 1242 2252
rect 1430 2248 1434 2252
rect 1694 2248 1698 2252
rect 1726 2248 1730 2252
rect 2022 2248 2026 2252
rect 2310 2248 2314 2252
rect 2374 2248 2378 2252
rect 2414 2248 2418 2252
rect 3430 2266 3434 2270
rect 3438 2268 3442 2272
rect 3462 2268 3466 2272
rect 3494 2268 3498 2272
rect 3526 2268 3530 2272
rect 3550 2268 3554 2272
rect 3558 2268 3562 2272
rect 3598 2268 3602 2272
rect 3614 2268 3618 2272
rect 3638 2268 3642 2272
rect 3726 2268 3730 2272
rect 3734 2266 3738 2270
rect 3862 2268 3866 2272
rect 2830 2258 2834 2262
rect 2870 2258 2874 2262
rect 2942 2258 2946 2262
rect 2990 2258 2994 2262
rect 3022 2258 3026 2262
rect 3086 2258 3090 2262
rect 3094 2258 3098 2262
rect 3126 2258 3130 2262
rect 3158 2258 3162 2262
rect 3198 2258 3202 2262
rect 3222 2258 3226 2262
rect 3230 2258 3234 2262
rect 3238 2258 3242 2262
rect 3270 2258 3274 2262
rect 3470 2258 3474 2262
rect 3502 2258 3506 2262
rect 3510 2258 3514 2262
rect 3566 2258 3570 2262
rect 3582 2258 3586 2262
rect 3622 2258 3626 2262
rect 3662 2258 3666 2262
rect 3774 2258 3778 2262
rect 3846 2259 3850 2263
rect 3910 2268 3914 2272
rect 3926 2268 3930 2272
rect 3974 2268 3978 2272
rect 3982 2268 3986 2272
rect 4142 2268 4146 2272
rect 4198 2268 4202 2272
rect 4206 2268 4210 2272
rect 4238 2268 4242 2272
rect 4262 2268 4266 2272
rect 4318 2268 4322 2272
rect 4446 2268 4450 2272
rect 4470 2268 4474 2272
rect 4486 2268 4490 2272
rect 4502 2268 4506 2272
rect 4526 2278 4530 2282
rect 4686 2278 4690 2282
rect 4774 2278 4778 2282
rect 4782 2278 4786 2282
rect 4822 2278 4826 2282
rect 4542 2268 4546 2272
rect 4758 2268 4762 2272
rect 4926 2278 4930 2282
rect 5022 2278 5026 2282
rect 5030 2278 5034 2282
rect 5126 2278 5130 2282
rect 4846 2268 4850 2272
rect 5038 2268 5042 2272
rect 5102 2268 5106 2272
rect 5294 2278 5298 2282
rect 5150 2268 5154 2272
rect 5174 2268 5178 2272
rect 3878 2258 3882 2262
rect 3894 2258 3898 2262
rect 3910 2258 3914 2262
rect 3966 2258 3970 2262
rect 3990 2258 3994 2262
rect 4014 2258 4018 2262
rect 4038 2258 4042 2262
rect 4078 2258 4082 2262
rect 4150 2258 4154 2262
rect 4158 2258 4162 2262
rect 4190 2258 4194 2262
rect 4206 2258 4210 2262
rect 4270 2258 4274 2262
rect 4310 2258 4314 2262
rect 4350 2259 4354 2263
rect 4478 2258 4482 2262
rect 4494 2258 4498 2262
rect 4550 2258 4554 2262
rect 4558 2258 4562 2262
rect 4566 2258 4570 2262
rect 4582 2258 4586 2262
rect 4590 2258 4594 2262
rect 4678 2258 4682 2262
rect 4718 2258 4722 2262
rect 4726 2258 4730 2262
rect 4774 2258 4778 2262
rect 4798 2258 4802 2262
rect 4806 2258 4810 2262
rect 4854 2258 4858 2262
rect 4918 2258 4922 2262
rect 4958 2258 4962 2262
rect 4982 2258 4986 2262
rect 5006 2258 5010 2262
rect 5110 2258 5114 2262
rect 5158 2258 5162 2262
rect 5198 2258 5202 2262
rect 5222 2258 5226 2262
rect 5262 2258 5266 2262
rect 2886 2248 2890 2252
rect 2942 2248 2946 2252
rect 3262 2248 3266 2252
rect 3302 2248 3306 2252
rect 3526 2248 3530 2252
rect 3534 2248 3538 2252
rect 3582 2248 3586 2252
rect 3878 2248 3882 2252
rect 3942 2248 3946 2252
rect 4174 2248 4178 2252
rect 4254 2248 4258 2252
rect 4286 2248 4290 2252
rect 4310 2248 4314 2252
rect 4398 2248 4402 2252
rect 4614 2248 4618 2252
rect 950 2238 954 2242
rect 1542 2238 1546 2242
rect 1862 2238 1866 2242
rect 3382 2238 3386 2242
rect 4134 2238 4138 2242
rect 750 2228 754 2232
rect 358 2218 362 2222
rect 982 2218 986 2222
rect 1214 2218 1218 2222
rect 1278 2218 1282 2222
rect 1574 2218 1578 2222
rect 1678 2218 1682 2222
rect 2198 2218 2202 2222
rect 2278 2218 2282 2222
rect 2294 2218 2298 2222
rect 2446 2218 2450 2222
rect 2526 2218 2530 2222
rect 2550 2218 2554 2222
rect 3006 2218 3010 2222
rect 3046 2218 3050 2222
rect 3174 2218 3178 2222
rect 3214 2218 3218 2222
rect 3542 2218 3546 2222
rect 3566 2218 3570 2222
rect 3718 2218 3722 2222
rect 3990 2218 3994 2222
rect 4998 2218 5002 2222
rect 5262 2218 5266 2222
rect 5286 2218 5290 2222
rect 330 2203 334 2207
rect 337 2203 341 2207
rect 1354 2203 1358 2207
rect 1361 2203 1365 2207
rect 2386 2203 2390 2207
rect 2393 2203 2397 2207
rect 3402 2203 3406 2207
rect 3409 2203 3413 2207
rect 4426 2203 4430 2207
rect 4433 2203 4437 2207
rect 62 2188 66 2192
rect 542 2188 546 2192
rect 614 2188 618 2192
rect 654 2188 658 2192
rect 742 2188 746 2192
rect 766 2188 770 2192
rect 782 2188 786 2192
rect 1206 2188 1210 2192
rect 1614 2188 1618 2192
rect 1678 2188 1682 2192
rect 1958 2188 1962 2192
rect 2118 2188 2122 2192
rect 2150 2188 2154 2192
rect 2190 2188 2194 2192
rect 2214 2188 2218 2192
rect 2246 2188 2250 2192
rect 2374 2188 2378 2192
rect 2414 2188 2418 2192
rect 2502 2188 2506 2192
rect 2542 2188 2546 2192
rect 2686 2188 2690 2192
rect 2718 2188 2722 2192
rect 2742 2188 2746 2192
rect 2814 2188 2818 2192
rect 3294 2188 3298 2192
rect 3334 2188 3338 2192
rect 3374 2188 3378 2192
rect 3558 2188 3562 2192
rect 3654 2188 3658 2192
rect 3774 2188 3778 2192
rect 3902 2188 3906 2192
rect 3966 2188 3970 2192
rect 3998 2188 4002 2192
rect 4454 2188 4458 2192
rect 4854 2188 4858 2192
rect 5070 2188 5074 2192
rect 5150 2188 5154 2192
rect 5182 2188 5186 2192
rect 5198 2188 5202 2192
rect 686 2178 690 2182
rect 3430 2178 3434 2182
rect 4310 2178 4314 2182
rect 4942 2178 4946 2182
rect 150 2168 154 2172
rect 166 2168 170 2172
rect 358 2168 362 2172
rect 862 2168 866 2172
rect 1550 2168 1554 2172
rect 1686 2168 1690 2172
rect 1742 2168 1746 2172
rect 1982 2168 1986 2172
rect 2302 2168 2306 2172
rect 2598 2168 2602 2172
rect 3142 2168 3146 2172
rect 3862 2168 3866 2172
rect 4174 2168 4178 2172
rect 5134 2168 5138 2172
rect 342 2158 346 2162
rect 670 2158 674 2162
rect 774 2158 778 2162
rect 822 2158 826 2162
rect 110 2148 114 2152
rect 174 2148 178 2152
rect 190 2148 194 2152
rect 222 2148 226 2152
rect 262 2148 266 2152
rect 358 2148 362 2152
rect 422 2148 426 2152
rect 446 2148 450 2152
rect 686 2148 690 2152
rect 806 2148 810 2152
rect 846 2158 850 2162
rect 1438 2158 1442 2162
rect 1566 2158 1570 2162
rect 1702 2158 1706 2162
rect 1710 2158 1714 2162
rect 1838 2158 1842 2162
rect 1886 2158 1890 2162
rect 1974 2158 1978 2162
rect 2318 2158 2322 2162
rect 2470 2158 2474 2162
rect 2854 2158 2858 2162
rect 3246 2158 3250 2162
rect 3310 2158 3314 2162
rect 846 2148 850 2152
rect 934 2148 938 2152
rect 1014 2148 1018 2152
rect 1070 2148 1074 2152
rect 1094 2148 1098 2152
rect 1110 2148 1114 2152
rect 1158 2148 1162 2152
rect 1270 2148 1274 2152
rect 1358 2148 1362 2152
rect 1374 2148 1378 2152
rect 1398 2148 1402 2152
rect 1406 2148 1410 2152
rect 1422 2148 1426 2152
rect 1430 2148 1434 2152
rect 1478 2148 1482 2152
rect 1550 2148 1554 2152
rect 1574 2148 1578 2152
rect 1590 2148 1594 2152
rect 1606 2148 1610 2152
rect 1646 2148 1650 2152
rect 1694 2148 1698 2152
rect 1726 2148 1730 2152
rect 1798 2148 1802 2152
rect 1846 2148 1850 2152
rect 1854 2148 1858 2152
rect 1902 2148 1906 2152
rect 1910 2148 1914 2152
rect 1934 2148 1938 2152
rect 1958 2148 1962 2152
rect 2030 2148 2034 2152
rect 2102 2148 2106 2152
rect 2142 2148 2146 2152
rect 2174 2148 2178 2152
rect 2230 2148 2234 2152
rect 2238 2148 2242 2152
rect 2254 2148 2258 2152
rect 2302 2148 2306 2152
rect 2326 2148 2330 2152
rect 2350 2148 2354 2152
rect 2358 2148 2362 2152
rect 2430 2148 2434 2152
rect 2438 2148 2442 2152
rect 2518 2148 2522 2152
rect 2574 2148 2578 2152
rect 2630 2148 2634 2152
rect 2670 2148 2674 2152
rect 2702 2148 2706 2152
rect 2758 2148 2762 2152
rect 2766 2148 2770 2152
rect 2918 2148 2922 2152
rect 2966 2148 2970 2152
rect 2974 2148 2978 2152
rect 6 2138 10 2142
rect 86 2138 90 2142
rect 182 2138 186 2142
rect 238 2138 242 2142
rect 366 2138 370 2142
rect 470 2138 474 2142
rect 486 2138 490 2142
rect 558 2138 562 2142
rect 662 2138 666 2142
rect 750 2138 754 2142
rect 758 2138 762 2142
rect 790 2138 794 2142
rect 798 2138 802 2142
rect 854 2138 858 2142
rect 870 2138 874 2142
rect 1006 2138 1010 2142
rect 1230 2138 1234 2142
rect 1246 2138 1250 2142
rect 1366 2138 1370 2142
rect 1374 2138 1378 2142
rect 1414 2138 1418 2142
rect 1454 2138 1458 2142
rect 1542 2138 1546 2142
rect 1574 2138 1578 2142
rect 1718 2138 1722 2142
rect 1734 2138 1738 2142
rect 1822 2138 1826 2142
rect 1942 2138 1946 2142
rect 1950 2138 1954 2142
rect 2038 2138 2042 2142
rect 2270 2138 2274 2142
rect 2278 2138 2282 2142
rect 2294 2138 2298 2142
rect 2462 2138 2466 2142
rect 2486 2138 2490 2142
rect 2494 2138 2498 2142
rect 2558 2138 2562 2142
rect 2574 2138 2578 2142
rect 2726 2138 2730 2142
rect 2782 2138 2786 2142
rect 3054 2147 3058 2151
rect 3126 2148 3130 2152
rect 3182 2148 3186 2152
rect 3230 2148 3234 2152
rect 3278 2148 3282 2152
rect 3294 2148 3298 2152
rect 3326 2148 3330 2152
rect 3350 2148 3354 2152
rect 3358 2148 3362 2152
rect 3390 2148 3394 2152
rect 3470 2148 3474 2152
rect 3534 2148 3538 2152
rect 3598 2148 3602 2152
rect 3630 2148 3634 2152
rect 3702 2148 3706 2152
rect 3814 2148 3818 2152
rect 3822 2148 3826 2152
rect 3838 2148 3842 2152
rect 3950 2158 3954 2162
rect 4230 2158 4234 2162
rect 4438 2158 4442 2162
rect 4630 2158 4634 2162
rect 4662 2158 4666 2162
rect 4702 2158 4706 2162
rect 3894 2148 3898 2152
rect 3918 2148 3922 2152
rect 3926 2148 3930 2152
rect 3950 2148 3954 2152
rect 3966 2148 3970 2152
rect 3982 2148 3986 2152
rect 4014 2148 4018 2152
rect 4022 2148 4026 2152
rect 4126 2148 4130 2152
rect 4214 2148 4218 2152
rect 4222 2148 4226 2152
rect 4246 2148 4250 2152
rect 4270 2148 4274 2152
rect 4294 2148 4298 2152
rect 4302 2148 4306 2152
rect 4382 2148 4386 2152
rect 4470 2148 4474 2152
rect 4502 2148 4506 2152
rect 4518 2148 4522 2152
rect 4526 2148 4530 2152
rect 4582 2148 4586 2152
rect 4646 2148 4650 2152
rect 4686 2148 4690 2152
rect 4814 2158 4818 2162
rect 5086 2158 5090 2162
rect 5166 2158 5170 2162
rect 4718 2148 4722 2152
rect 4726 2148 4730 2152
rect 2830 2138 2834 2142
rect 2878 2138 2882 2142
rect 3006 2138 3010 2142
rect 3062 2138 3066 2142
rect 3222 2138 3226 2142
rect 3286 2138 3290 2142
rect 3710 2138 3714 2142
rect 3782 2138 3786 2142
rect 3830 2138 3834 2142
rect 3862 2138 3866 2142
rect 3878 2138 3882 2142
rect 3974 2138 3978 2142
rect 4046 2138 4050 2142
rect 4054 2138 4058 2142
rect 4158 2138 4162 2142
rect 4190 2138 4194 2142
rect 4222 2138 4226 2142
rect 4766 2147 4770 2151
rect 4838 2148 4842 2152
rect 4886 2148 4890 2152
rect 4918 2148 4922 2152
rect 4926 2148 4930 2152
rect 4974 2148 4978 2152
rect 4982 2148 4986 2152
rect 5014 2148 5018 2152
rect 5022 2148 5026 2152
rect 5030 2148 5034 2152
rect 5054 2148 5058 2152
rect 5118 2148 5122 2152
rect 5134 2148 5138 2152
rect 5150 2148 5154 2152
rect 5174 2148 5178 2152
rect 5230 2148 5234 2152
rect 5254 2148 5258 2152
rect 4374 2138 4378 2142
rect 4462 2138 4466 2142
rect 4598 2138 4602 2142
rect 4654 2138 4658 2142
rect 4678 2138 4682 2142
rect 4734 2138 4738 2142
rect 4750 2138 4754 2142
rect 4910 2138 4914 2142
rect 5102 2138 5106 2142
rect 5110 2138 5114 2142
rect 5142 2138 5146 2142
rect 206 2128 210 2132
rect 286 2128 290 2132
rect 710 2128 714 2132
rect 1086 2128 1090 2132
rect 1142 2128 1146 2132
rect 1606 2128 1610 2132
rect 1630 2128 1634 2132
rect 1654 2128 1658 2132
rect 1670 2128 1674 2132
rect 1806 2128 1810 2132
rect 1886 2128 1890 2132
rect 2254 2128 2258 2132
rect 2286 2128 2290 2132
rect 2614 2128 2618 2132
rect 3022 2128 3026 2132
rect 3494 2128 3498 2132
rect 4286 2128 4290 2132
rect 4470 2128 4474 2132
rect 4670 2128 4674 2132
rect 4870 2128 4874 2132
rect 4990 2128 4994 2132
rect 5078 2128 5082 2132
rect 5190 2128 5194 2132
rect 318 2118 322 2122
rect 638 2118 642 2122
rect 1062 2118 1066 2122
rect 1222 2118 1226 2122
rect 1534 2118 1538 2122
rect 2086 2118 2090 2122
rect 2414 2118 2418 2122
rect 2478 2118 2482 2122
rect 2542 2118 2546 2122
rect 2622 2118 2626 2122
rect 2646 2118 2650 2122
rect 2742 2118 2746 2122
rect 2814 2118 2818 2122
rect 2846 2118 2850 2122
rect 2958 2118 2962 2122
rect 3118 2118 3122 2122
rect 3166 2118 3170 2122
rect 3206 2118 3210 2122
rect 3246 2118 3250 2122
rect 3262 2118 3266 2122
rect 3454 2118 3458 2122
rect 3518 2118 3522 2122
rect 3582 2118 3586 2122
rect 3614 2118 3618 2122
rect 4198 2118 4202 2122
rect 4534 2118 4538 2122
rect 4630 2118 4634 2122
rect 4854 2118 4858 2122
rect 4902 2118 4906 2122
rect 5046 2118 5050 2122
rect 5086 2118 5090 2122
rect 850 2103 854 2107
rect 857 2103 861 2107
rect 1874 2103 1878 2107
rect 1881 2103 1885 2107
rect 2890 2103 2894 2107
rect 2897 2103 2901 2107
rect 3922 2103 3926 2107
rect 3929 2103 3933 2107
rect 4938 2103 4942 2107
rect 4945 2103 4949 2107
rect 254 2088 258 2092
rect 350 2088 354 2092
rect 534 2088 538 2092
rect 574 2088 578 2092
rect 830 2088 834 2092
rect 934 2088 938 2092
rect 1070 2088 1074 2092
rect 1102 2088 1106 2092
rect 1270 2088 1274 2092
rect 1366 2088 1370 2092
rect 1390 2088 1394 2092
rect 1438 2088 1442 2092
rect 1598 2088 1602 2092
rect 1710 2088 1714 2092
rect 1854 2088 1858 2092
rect 1910 2088 1914 2092
rect 2246 2088 2250 2092
rect 2310 2088 2314 2092
rect 2422 2088 2426 2092
rect 3110 2088 3114 2092
rect 3166 2088 3170 2092
rect 3238 2088 3242 2092
rect 3270 2088 3274 2092
rect 3342 2088 3346 2092
rect 3398 2088 3402 2092
rect 3606 2088 3610 2092
rect 3646 2088 3650 2092
rect 3662 2088 3666 2092
rect 3710 2088 3714 2092
rect 3734 2088 3738 2092
rect 3774 2088 3778 2092
rect 3886 2088 3890 2092
rect 4014 2088 4018 2092
rect 4206 2088 4210 2092
rect 4366 2088 4370 2092
rect 4982 2088 4986 2092
rect 5022 2088 5026 2092
rect 5118 2088 5122 2092
rect 5222 2088 5226 2092
rect 286 2078 290 2082
rect 382 2078 386 2082
rect 462 2078 466 2082
rect 542 2078 546 2082
rect 550 2078 554 2082
rect 558 2078 562 2082
rect 566 2078 570 2082
rect 606 2078 610 2082
rect 942 2078 946 2082
rect 1158 2078 1162 2082
rect 1238 2078 1242 2082
rect 1334 2078 1338 2082
rect 1398 2078 1402 2082
rect 1582 2078 1586 2082
rect 6 2068 10 2072
rect 70 2068 74 2072
rect 86 2068 90 2072
rect 190 2068 194 2072
rect 246 2068 250 2072
rect 318 2068 322 2072
rect 326 2068 330 2072
rect 398 2068 402 2072
rect 606 2068 610 2072
rect 662 2068 666 2072
rect 734 2068 738 2072
rect 790 2068 794 2072
rect 822 2068 826 2072
rect 862 2068 866 2072
rect 878 2068 882 2072
rect 910 2068 914 2072
rect 926 2068 930 2072
rect 1006 2068 1010 2072
rect 1078 2068 1082 2072
rect 110 2058 114 2062
rect 198 2058 202 2062
rect 222 2058 226 2062
rect 230 2058 234 2062
rect 238 2058 242 2062
rect 270 2058 274 2062
rect 286 2058 290 2062
rect 310 2058 314 2062
rect 1086 2066 1090 2070
rect 1118 2068 1122 2072
rect 1166 2068 1170 2072
rect 1198 2068 1202 2072
rect 1214 2068 1218 2072
rect 1294 2068 1298 2072
rect 1310 2068 1314 2072
rect 1326 2068 1330 2072
rect 1366 2068 1370 2072
rect 1398 2068 1402 2072
rect 1438 2068 1442 2072
rect 1454 2068 1458 2072
rect 1462 2068 1466 2072
rect 1494 2068 1498 2072
rect 1558 2068 1562 2072
rect 1606 2078 1610 2082
rect 1630 2078 1634 2082
rect 1654 2078 1658 2082
rect 2238 2078 2242 2082
rect 2414 2078 2418 2082
rect 2470 2078 2474 2082
rect 2734 2078 2738 2082
rect 2758 2078 2762 2082
rect 2822 2078 2826 2082
rect 2838 2078 2842 2082
rect 1630 2068 1634 2072
rect 1646 2068 1650 2072
rect 1806 2068 1810 2072
rect 1846 2068 1850 2072
rect 1878 2068 1882 2072
rect 1886 2068 1890 2072
rect 1918 2068 1922 2072
rect 1974 2068 1978 2072
rect 2038 2068 2042 2072
rect 2078 2068 2082 2072
rect 2102 2068 2106 2072
rect 2110 2068 2114 2072
rect 2150 2068 2154 2072
rect 2254 2068 2258 2072
rect 2302 2068 2306 2072
rect 2558 2068 2562 2072
rect 2662 2068 2666 2072
rect 2710 2068 2714 2072
rect 2774 2068 2778 2072
rect 2910 2078 2914 2082
rect 2966 2078 2970 2082
rect 3078 2078 3082 2082
rect 3334 2078 3338 2082
rect 3390 2078 3394 2082
rect 3614 2078 3618 2082
rect 3654 2078 3658 2082
rect 3814 2078 3818 2082
rect 2918 2068 2922 2072
rect 3062 2068 3066 2072
rect 3190 2068 3194 2072
rect 3326 2068 3330 2072
rect 3358 2068 3362 2072
rect 3406 2068 3410 2072
rect 3470 2068 3474 2072
rect 3478 2068 3482 2072
rect 3550 2068 3554 2072
rect 3622 2068 3626 2072
rect 3670 2068 3674 2072
rect 3686 2068 3690 2072
rect 3718 2068 3722 2072
rect 3726 2068 3730 2072
rect 3758 2068 3762 2072
rect 3806 2068 3810 2072
rect 3838 2068 3842 2072
rect 3878 2068 3882 2072
rect 3910 2068 3914 2072
rect 4038 2068 4042 2072
rect 4062 2078 4066 2082
rect 4166 2078 4170 2082
rect 4238 2078 4242 2082
rect 4862 2078 4866 2082
rect 5214 2078 5218 2082
rect 4142 2068 4146 2072
rect 4190 2068 4194 2072
rect 4206 2068 4210 2072
rect 4230 2068 4234 2072
rect 4286 2068 4290 2072
rect 4358 2068 4362 2072
rect 4390 2068 4394 2072
rect 4398 2068 4402 2072
rect 4462 2068 4466 2072
rect 4470 2068 4474 2072
rect 4550 2068 4554 2072
rect 4598 2068 4602 2072
rect 4606 2068 4610 2072
rect 4630 2068 4634 2072
rect 4662 2068 4666 2072
rect 4694 2068 4698 2072
rect 4830 2068 4834 2072
rect 5054 2068 5058 2072
rect 5070 2068 5074 2072
rect 470 2058 474 2062
rect 494 2059 498 2063
rect 526 2058 530 2062
rect 582 2058 586 2062
rect 614 2058 618 2062
rect 726 2058 730 2062
rect 790 2058 794 2062
rect 814 2058 818 2062
rect 870 2058 874 2062
rect 878 2058 882 2062
rect 926 2058 930 2062
rect 950 2058 954 2062
rect 1014 2058 1018 2062
rect 1110 2058 1114 2062
rect 1126 2058 1130 2062
rect 1142 2058 1146 2062
rect 1174 2058 1178 2062
rect 1222 2058 1226 2062
rect 1246 2058 1250 2062
rect 1254 2058 1258 2062
rect 1278 2058 1282 2062
rect 1294 2058 1298 2062
rect 1318 2058 1322 2062
rect 1358 2058 1362 2062
rect 1374 2058 1378 2062
rect 1422 2058 1426 2062
rect 1462 2058 1466 2062
rect 1518 2058 1522 2062
rect 1558 2058 1562 2062
rect 1566 2058 1570 2062
rect 1606 2058 1610 2062
rect 1654 2058 1658 2062
rect 1670 2058 1674 2062
rect 1694 2058 1698 2062
rect 1790 2059 1794 2063
rect 1838 2058 1842 2062
rect 1870 2058 1874 2062
rect 1902 2058 1906 2062
rect 1918 2058 1922 2062
rect 1942 2058 1946 2062
rect 1966 2058 1970 2062
rect 2030 2058 2034 2062
rect 2086 2058 2090 2062
rect 2118 2058 2122 2062
rect 2126 2058 2130 2062
rect 2166 2059 2170 2063
rect 2262 2058 2266 2062
rect 2270 2058 2274 2062
rect 2326 2058 2330 2062
rect 2358 2058 2362 2062
rect 2430 2058 2434 2062
rect 2438 2058 2442 2062
rect 2486 2058 2490 2062
rect 2598 2058 2602 2062
rect 2630 2059 2634 2063
rect 2678 2058 2682 2062
rect 2718 2058 2722 2062
rect 2742 2058 2746 2062
rect 2814 2058 2818 2062
rect 2878 2058 2882 2062
rect 2926 2058 2930 2062
rect 2950 2058 2954 2062
rect 3014 2058 3018 2062
rect 3046 2059 3050 2063
rect 3102 2058 3106 2062
rect 3126 2058 3130 2062
rect 3134 2058 3138 2062
rect 3150 2058 3154 2062
rect 3174 2058 3178 2062
rect 3182 2058 3186 2062
rect 3214 2058 3218 2062
rect 3246 2058 3250 2062
rect 3286 2058 3290 2062
rect 3294 2058 3298 2062
rect 3318 2058 3322 2062
rect 3350 2058 3354 2062
rect 3366 2058 3370 2062
rect 3414 2058 3418 2062
rect 3438 2058 3442 2062
rect 3446 2058 3450 2062
rect 3470 2058 3474 2062
rect 3558 2058 3562 2062
rect 3598 2058 3602 2062
rect 3630 2058 3634 2062
rect 3678 2058 3682 2062
rect 3694 2058 3698 2062
rect 3710 2058 3714 2062
rect 3734 2058 3738 2062
rect 3750 2058 3754 2062
rect 3870 2058 3874 2062
rect 3902 2058 3906 2062
rect 3998 2058 4002 2062
rect 4030 2058 4034 2062
rect 4046 2058 4050 2062
rect 4086 2058 4090 2062
rect 4102 2058 4106 2062
rect 4126 2058 4130 2062
rect 4134 2058 4138 2062
rect 4150 2058 4154 2062
rect 4198 2058 4202 2062
rect 4230 2058 4234 2062
rect 4302 2059 4306 2063
rect 5110 2068 5114 2072
rect 5198 2068 5202 2072
rect 5230 2068 5234 2072
rect 5278 2068 5282 2072
rect 4350 2058 4354 2062
rect 4382 2058 4386 2062
rect 4406 2058 4410 2062
rect 4478 2058 4482 2062
rect 4502 2058 4506 2062
rect 4510 2058 4514 2062
rect 4526 2058 4530 2062
rect 4534 2058 4538 2062
rect 4558 2058 4562 2062
rect 4566 2058 4570 2062
rect 4614 2058 4618 2062
rect 4630 2058 4634 2062
rect 4654 2058 4658 2062
rect 4670 2058 4674 2062
rect 4710 2058 4714 2062
rect 4734 2058 4738 2062
rect 4742 2058 4746 2062
rect 4806 2058 4810 2062
rect 4886 2058 4890 2062
rect 4902 2058 4906 2062
rect 4958 2058 4962 2062
rect 4966 2058 4970 2062
rect 4990 2058 4994 2062
rect 5006 2058 5010 2062
rect 5014 2058 5018 2062
rect 5038 2058 5042 2062
rect 5062 2058 5066 2062
rect 5086 2058 5090 2062
rect 5102 2058 5106 2062
rect 5158 2058 5162 2062
rect 5238 2058 5242 2062
rect 5246 2058 5250 2062
rect 5254 2058 5258 2062
rect 5278 2058 5282 2062
rect 174 2048 178 2052
rect 294 2048 298 2052
rect 342 2048 346 2052
rect 630 2048 634 2052
rect 814 2048 818 2052
rect 830 2048 834 2052
rect 1190 2048 1194 2052
rect 1238 2048 1242 2052
rect 1406 2048 1410 2052
rect 1438 2048 1442 2052
rect 1486 2048 1490 2052
rect 1534 2048 1538 2052
rect 1822 2048 1826 2052
rect 1854 2048 1858 2052
rect 1950 2048 1954 2052
rect 2102 2048 2106 2052
rect 2134 2048 2138 2052
rect 2502 2048 2506 2052
rect 2934 2048 2938 2052
rect 3214 2048 3218 2052
rect 3382 2048 3386 2052
rect 3646 2048 3650 2052
rect 3782 2048 3786 2052
rect 3790 2048 3794 2052
rect 3846 2048 3850 2052
rect 4174 2048 4178 2052
rect 4334 2048 4338 2052
rect 4350 2048 4354 2052
rect 4366 2048 4370 2052
rect 4446 2048 4450 2052
rect 4494 2048 4498 2052
rect 4582 2048 4586 2052
rect 4638 2048 4642 2052
rect 4654 2048 4658 2052
rect 5078 2048 5082 2052
rect 5086 2048 5090 2052
rect 358 2038 362 2042
rect 670 2038 674 2042
rect 766 2038 770 2042
rect 798 2038 802 2042
rect 902 2038 906 2042
rect 1726 2038 1730 2042
rect 1838 2038 1842 2042
rect 1926 2038 1930 2042
rect 1966 2038 1970 2042
rect 1982 2038 1986 2042
rect 2950 2038 2954 2042
rect 3078 2038 3082 2042
rect 3366 2038 3370 2042
rect 3518 2038 3522 2042
rect 4406 2038 4410 2042
rect 4750 2038 4754 2042
rect 5134 2038 5138 2042
rect 1174 2028 1178 2032
rect 1686 2028 1690 2032
rect 2382 2028 2386 2032
rect 3198 2028 3202 2032
rect 3982 2028 3986 2032
rect 782 2018 786 2022
rect 886 2018 890 2022
rect 966 2018 970 2022
rect 1206 2018 1210 2022
rect 1518 2018 1522 2022
rect 2230 2018 2234 2022
rect 2310 2018 2314 2022
rect 2342 2018 2346 2022
rect 2454 2018 2458 2022
rect 2486 2018 2490 2022
rect 2566 2018 2570 2022
rect 2726 2018 2730 2022
rect 2750 2018 2754 2022
rect 3238 2018 3242 2022
rect 4478 2018 4482 2022
rect 4686 2018 4690 2022
rect 4726 2018 4730 2022
rect 330 2003 334 2007
rect 337 2003 341 2007
rect 1354 2003 1358 2007
rect 1361 2003 1365 2007
rect 2386 2003 2390 2007
rect 2393 2003 2397 2007
rect 3402 2003 3406 2007
rect 3409 2003 3413 2007
rect 4426 2003 4430 2007
rect 4433 2003 4437 2007
rect 166 1988 170 1992
rect 302 1988 306 1992
rect 334 1988 338 1992
rect 750 1988 754 1992
rect 1118 1988 1122 1992
rect 1462 1988 1466 1992
rect 1598 1988 1602 1992
rect 1758 1988 1762 1992
rect 1782 1988 1786 1992
rect 1990 1988 1994 1992
rect 2030 1988 2034 1992
rect 2110 1988 2114 1992
rect 2134 1988 2138 1992
rect 2374 1988 2378 1992
rect 2622 1988 2626 1992
rect 2694 1988 2698 1992
rect 2806 1988 2810 1992
rect 3254 1988 3258 1992
rect 3278 1988 3282 1992
rect 3526 1988 3530 1992
rect 4654 1988 4658 1992
rect 4782 1988 4786 1992
rect 4870 1988 4874 1992
rect 62 1978 66 1982
rect 1134 1978 1138 1982
rect 1334 1978 1338 1982
rect 3126 1978 3130 1982
rect 230 1968 234 1972
rect 438 1968 442 1972
rect 622 1968 626 1972
rect 734 1968 738 1972
rect 1822 1968 1826 1972
rect 2062 1968 2066 1972
rect 2478 1968 2482 1972
rect 2774 1968 2778 1972
rect 3014 1968 3018 1972
rect 3030 1968 3034 1972
rect 4110 1968 4114 1972
rect 4206 1968 4210 1972
rect 5062 1968 5066 1972
rect 5262 1968 5266 1972
rect 174 1958 178 1962
rect 246 1958 250 1962
rect 278 1958 282 1962
rect 286 1958 290 1962
rect 422 1958 426 1962
rect 758 1958 762 1962
rect 814 1958 818 1962
rect 934 1958 938 1962
rect 118 1948 122 1952
rect 174 1948 178 1952
rect 190 1948 194 1952
rect 262 1948 266 1952
rect 302 1948 306 1952
rect 318 1948 322 1952
rect 374 1948 378 1952
rect 390 1948 394 1952
rect 470 1948 474 1952
rect 502 1947 506 1951
rect 574 1948 578 1952
rect 654 1948 658 1952
rect 694 1948 698 1952
rect 758 1948 762 1952
rect 774 1948 778 1952
rect 798 1948 802 1952
rect 870 1948 874 1952
rect 958 1948 962 1952
rect 982 1948 986 1952
rect 990 1948 994 1952
rect 1022 1948 1026 1952
rect 1062 1948 1066 1952
rect 1134 1948 1138 1952
rect 1158 1958 1162 1962
rect 1214 1958 1218 1962
rect 1422 1958 1426 1962
rect 1558 1958 1562 1962
rect 1614 1958 1618 1962
rect 1774 1958 1778 1962
rect 1838 1958 1842 1962
rect 1870 1958 1874 1962
rect 1886 1958 1890 1962
rect 1910 1958 1914 1962
rect 2078 1958 2082 1962
rect 2150 1958 2154 1962
rect 2598 1958 2602 1962
rect 2614 1958 2618 1962
rect 2678 1958 2682 1962
rect 2790 1958 2794 1962
rect 2798 1958 2802 1962
rect 2814 1958 2818 1962
rect 2838 1958 2842 1962
rect 2862 1958 2866 1962
rect 2934 1958 2938 1962
rect 3046 1958 3050 1962
rect 3062 1958 3066 1962
rect 3070 1958 3074 1962
rect 3086 1958 3090 1962
rect 3142 1958 3146 1962
rect 3174 1958 3178 1962
rect 3430 1958 3434 1962
rect 3510 1958 3514 1962
rect 3982 1958 3986 1962
rect 4078 1958 4082 1962
rect 4318 1958 4322 1962
rect 1174 1948 1178 1952
rect 1198 1948 1202 1952
rect 1214 1948 1218 1952
rect 6 1938 10 1942
rect 86 1938 90 1942
rect 198 1938 202 1942
rect 222 1938 226 1942
rect 254 1938 258 1942
rect 310 1938 314 1942
rect 342 1938 346 1942
rect 366 1938 370 1942
rect 398 1938 402 1942
rect 206 1928 210 1932
rect 422 1928 426 1932
rect 454 1928 458 1932
rect 646 1938 650 1942
rect 670 1938 674 1942
rect 790 1938 794 1942
rect 806 1938 810 1942
rect 862 1938 866 1942
rect 998 1938 1002 1942
rect 1038 1938 1042 1942
rect 1126 1938 1130 1942
rect 1182 1938 1186 1942
rect 1190 1938 1194 1942
rect 1246 1947 1250 1951
rect 1318 1948 1322 1952
rect 1334 1948 1338 1952
rect 1374 1948 1378 1952
rect 1398 1948 1402 1952
rect 1414 1948 1418 1952
rect 1422 1948 1426 1952
rect 1526 1947 1530 1951
rect 1566 1948 1570 1952
rect 1574 1948 1578 1952
rect 1598 1948 1602 1952
rect 1622 1948 1626 1952
rect 1654 1948 1658 1952
rect 1670 1948 1674 1952
rect 1710 1948 1714 1952
rect 1726 1948 1730 1952
rect 1742 1948 1746 1952
rect 1814 1948 1818 1952
rect 1854 1948 1858 1952
rect 1894 1948 1898 1952
rect 1342 1938 1346 1942
rect 1366 1938 1370 1942
rect 1398 1938 1402 1942
rect 1430 1938 1434 1942
rect 1454 1938 1458 1942
rect 1510 1938 1514 1942
rect 1582 1938 1586 1942
rect 1590 1938 1594 1942
rect 1630 1938 1634 1942
rect 1694 1938 1698 1942
rect 1702 1938 1706 1942
rect 1734 1938 1738 1942
rect 1790 1938 1794 1942
rect 1838 1938 1842 1942
rect 1934 1948 1938 1952
rect 1942 1948 1946 1952
rect 1974 1948 1978 1952
rect 1990 1948 1994 1952
rect 2006 1948 2010 1952
rect 2014 1948 2018 1952
rect 2046 1948 2050 1952
rect 2054 1948 2058 1952
rect 2086 1948 2090 1952
rect 2118 1948 2122 1952
rect 2126 1948 2130 1952
rect 2286 1948 2290 1952
rect 2358 1948 2362 1952
rect 2406 1948 2410 1952
rect 2438 1948 2442 1952
rect 2494 1948 2498 1952
rect 2502 1948 2506 1952
rect 2566 1948 2570 1952
rect 2590 1948 2594 1952
rect 2686 1948 2690 1952
rect 2766 1948 2770 1952
rect 1998 1938 2002 1942
rect 2054 1938 2058 1942
rect 2086 1938 2090 1942
rect 2110 1938 2114 1942
rect 2126 1938 2130 1942
rect 2222 1938 2226 1942
rect 2262 1938 2266 1942
rect 2294 1938 2298 1942
rect 2470 1938 2474 1942
rect 2502 1938 2506 1942
rect 2630 1938 2634 1942
rect 2662 1938 2666 1942
rect 2670 1938 2674 1942
rect 2774 1938 2778 1942
rect 2814 1938 2818 1942
rect 2846 1948 2850 1952
rect 2918 1948 2922 1952
rect 2966 1947 2970 1951
rect 3046 1948 3050 1952
rect 3086 1948 3090 1952
rect 3126 1948 3130 1952
rect 3158 1948 3162 1952
rect 3230 1948 3234 1952
rect 3270 1948 3274 1952
rect 3294 1948 3298 1952
rect 3366 1947 3370 1951
rect 3446 1948 3450 1952
rect 3494 1948 3498 1952
rect 3502 1948 3506 1952
rect 3526 1948 3530 1952
rect 3542 1948 3546 1952
rect 3598 1948 3602 1952
rect 3606 1948 3610 1952
rect 3734 1947 3738 1951
rect 3806 1948 3810 1952
rect 3822 1948 3826 1952
rect 3902 1948 3906 1952
rect 3998 1948 4002 1952
rect 4046 1948 4050 1952
rect 4062 1948 4066 1952
rect 4070 1948 4074 1952
rect 4094 1948 4098 1952
rect 4142 1948 4146 1952
rect 4166 1948 4170 1952
rect 4614 1958 4618 1962
rect 4270 1947 4274 1951
rect 4342 1948 4346 1952
rect 4358 1948 4362 1952
rect 4766 1958 4770 1962
rect 4798 1958 4802 1962
rect 4830 1958 4834 1962
rect 4430 1947 4434 1951
rect 4566 1947 4570 1951
rect 4630 1948 4634 1952
rect 4638 1948 4642 1952
rect 4726 1948 4730 1952
rect 4870 1948 4874 1952
rect 4982 1947 4986 1951
rect 5022 1948 5026 1952
rect 5046 1958 5050 1962
rect 5126 1948 5130 1952
rect 5222 1948 5226 1952
rect 5286 1948 5290 1952
rect 2862 1938 2866 1942
rect 2886 1938 2890 1942
rect 2902 1938 2906 1942
rect 2934 1938 2938 1942
rect 2950 1938 2954 1942
rect 3038 1938 3042 1942
rect 3102 1938 3106 1942
rect 3150 1938 3154 1942
rect 3262 1938 3266 1942
rect 3414 1938 3418 1942
rect 3454 1938 3458 1942
rect 3462 1938 3466 1942
rect 3534 1938 3538 1942
rect 3638 1938 3642 1942
rect 3654 1938 3658 1942
rect 3878 1938 3882 1942
rect 3910 1938 3914 1942
rect 4014 1938 4018 1942
rect 4078 1938 4082 1942
rect 4102 1938 4106 1942
rect 4190 1938 4194 1942
rect 4262 1938 4266 1942
rect 4286 1938 4290 1942
rect 4302 1938 4306 1942
rect 4318 1938 4322 1942
rect 4350 1938 4354 1942
rect 4390 1938 4394 1942
rect 4414 1938 4418 1942
rect 4518 1938 4522 1942
rect 4582 1938 4586 1942
rect 4598 1938 4602 1942
rect 4646 1938 4650 1942
rect 4750 1938 4754 1942
rect 4790 1938 4794 1942
rect 4822 1938 4826 1942
rect 4846 1938 4850 1942
rect 4998 1938 5002 1942
rect 5014 1938 5018 1942
rect 5046 1938 5050 1942
rect 5062 1938 5066 1942
rect 5150 1938 5154 1942
rect 5214 1938 5218 1942
rect 5278 1938 5282 1942
rect 590 1928 594 1932
rect 630 1928 634 1932
rect 638 1928 642 1932
rect 966 1928 970 1932
rect 1246 1928 1250 1932
rect 1670 1928 1674 1932
rect 1694 1928 1698 1932
rect 1798 1928 1802 1932
rect 1902 1928 1906 1932
rect 1918 1928 1922 1932
rect 1958 1928 1962 1932
rect 2534 1928 2538 1932
rect 2542 1928 2546 1932
rect 2558 1928 2562 1932
rect 2582 1928 2586 1932
rect 2606 1928 2610 1932
rect 2638 1928 2642 1932
rect 2654 1928 2658 1932
rect 2710 1928 2714 1932
rect 2750 1928 2754 1932
rect 3102 1928 3106 1932
rect 3198 1928 3202 1932
rect 3222 1928 3226 1932
rect 3366 1928 3370 1932
rect 3398 1928 3402 1932
rect 3582 1928 3586 1932
rect 3638 1928 3642 1932
rect 3862 1928 3866 1932
rect 4478 1928 4482 1932
rect 4902 1928 4906 1932
rect 5262 1928 5266 1932
rect 278 1918 282 1922
rect 430 1918 434 1922
rect 1390 1918 1394 1922
rect 1638 1918 1642 1922
rect 1710 1918 1714 1922
rect 1926 1918 1930 1922
rect 2166 1918 2170 1922
rect 2230 1918 2234 1922
rect 2334 1918 2338 1922
rect 2422 1918 2426 1922
rect 2574 1918 2578 1922
rect 2734 1918 2738 1922
rect 2790 1918 2794 1922
rect 2806 1918 2810 1922
rect 2854 1918 2858 1922
rect 2870 1918 2874 1922
rect 3302 1918 3306 1922
rect 3414 1918 3418 1922
rect 3558 1918 3562 1922
rect 3646 1918 3650 1922
rect 3670 1918 3674 1922
rect 3854 1918 3858 1922
rect 3870 1918 3874 1922
rect 3966 1918 3970 1922
rect 3982 1918 3986 1922
rect 4918 1918 4922 1922
rect 5166 1918 5170 1922
rect 850 1903 854 1907
rect 857 1903 861 1907
rect 1874 1903 1878 1907
rect 1881 1903 1885 1907
rect 2890 1903 2894 1907
rect 2897 1903 2901 1907
rect 3922 1903 3926 1907
rect 3929 1903 3933 1907
rect 4938 1903 4942 1907
rect 4945 1903 4949 1907
rect 6 1888 10 1892
rect 246 1888 250 1892
rect 270 1888 274 1892
rect 310 1888 314 1892
rect 398 1888 402 1892
rect 598 1888 602 1892
rect 622 1888 626 1892
rect 830 1888 834 1892
rect 1014 1888 1018 1892
rect 1134 1888 1138 1892
rect 1358 1888 1362 1892
rect 1526 1888 1530 1892
rect 1542 1888 1546 1892
rect 1614 1888 1618 1892
rect 1710 1888 1714 1892
rect 2022 1888 2026 1892
rect 2038 1888 2042 1892
rect 2214 1888 2218 1892
rect 2286 1888 2290 1892
rect 2326 1888 2330 1892
rect 2446 1888 2450 1892
rect 2510 1888 2514 1892
rect 2558 1888 2562 1892
rect 2646 1888 2650 1892
rect 3062 1888 3066 1892
rect 3094 1888 3098 1892
rect 3110 1888 3114 1892
rect 3206 1888 3210 1892
rect 3286 1888 3290 1892
rect 3454 1888 3458 1892
rect 3582 1888 3586 1892
rect 3606 1888 3610 1892
rect 3774 1888 3778 1892
rect 3862 1888 3866 1892
rect 3942 1888 3946 1892
rect 4006 1888 4010 1892
rect 4102 1888 4106 1892
rect 4150 1888 4154 1892
rect 4430 1888 4434 1892
rect 4470 1888 4474 1892
rect 4494 1888 4498 1892
rect 4526 1888 4530 1892
rect 4750 1888 4754 1892
rect 4838 1888 4842 1892
rect 4878 1888 4882 1892
rect 4918 1888 4922 1892
rect 4982 1888 4986 1892
rect 5134 1888 5138 1892
rect 5158 1888 5162 1892
rect 5190 1888 5194 1892
rect 5238 1888 5242 1892
rect 70 1878 74 1882
rect 102 1878 106 1882
rect 182 1878 186 1882
rect 278 1878 282 1882
rect 318 1878 322 1882
rect 462 1878 466 1882
rect 510 1878 514 1882
rect 630 1878 634 1882
rect 742 1878 746 1882
rect 934 1878 938 1882
rect 1126 1878 1130 1882
rect 1558 1878 1562 1882
rect 1574 1878 1578 1882
rect 126 1868 130 1872
rect 142 1868 146 1872
rect 262 1868 266 1872
rect 286 1868 290 1872
rect 334 1868 338 1872
rect 542 1868 546 1872
rect 614 1868 618 1872
rect 686 1868 690 1872
rect 702 1868 706 1872
rect 726 1868 730 1872
rect 750 1868 754 1872
rect 766 1868 770 1872
rect 806 1868 810 1872
rect 878 1868 882 1872
rect 1022 1868 1026 1872
rect 1070 1868 1074 1872
rect 70 1859 74 1863
rect 118 1858 122 1862
rect 150 1858 154 1862
rect 190 1858 194 1862
rect 254 1858 258 1862
rect 294 1858 298 1862
rect 342 1858 346 1862
rect 358 1858 362 1862
rect 382 1858 386 1862
rect 390 1858 394 1862
rect 462 1859 466 1863
rect 1110 1868 1114 1872
rect 1158 1868 1162 1872
rect 1190 1868 1194 1872
rect 1262 1868 1266 1872
rect 1318 1868 1322 1872
rect 1326 1868 1330 1872
rect 1430 1868 1434 1872
rect 1462 1868 1466 1872
rect 2030 1878 2034 1882
rect 2422 1878 2426 1882
rect 2462 1878 2466 1882
rect 2478 1878 2482 1882
rect 2486 1878 2490 1882
rect 2518 1878 2522 1882
rect 2638 1878 2642 1882
rect 2742 1878 2746 1882
rect 2790 1878 2794 1882
rect 3102 1878 3106 1882
rect 3254 1878 3258 1882
rect 3262 1878 3266 1882
rect 3414 1878 3418 1882
rect 3518 1878 3522 1882
rect 3614 1878 3618 1882
rect 3622 1878 3626 1882
rect 1606 1868 1610 1872
rect 1678 1868 1682 1872
rect 1726 1868 1730 1872
rect 1774 1868 1778 1872
rect 2014 1868 2018 1872
rect 2054 1868 2058 1872
rect 2158 1868 2162 1872
rect 2174 1868 2178 1872
rect 2222 1868 2226 1872
rect 2262 1868 2266 1872
rect 2270 1868 2274 1872
rect 2318 1868 2322 1872
rect 2334 1868 2338 1872
rect 2342 1868 2346 1872
rect 2414 1868 2418 1872
rect 2454 1868 2458 1872
rect 2574 1868 2578 1872
rect 2614 1868 2618 1872
rect 2814 1868 2818 1872
rect 2870 1868 2874 1872
rect 2902 1868 2906 1872
rect 2950 1868 2954 1872
rect 2990 1868 2994 1872
rect 3046 1868 3050 1872
rect 3070 1868 3074 1872
rect 3078 1868 3082 1872
rect 3126 1868 3130 1872
rect 3158 1868 3162 1872
rect 3238 1868 3242 1872
rect 3254 1868 3258 1872
rect 3366 1868 3370 1872
rect 3390 1868 3394 1872
rect 3598 1868 3602 1872
rect 3638 1868 3642 1872
rect 3646 1868 3650 1872
rect 3686 1868 3690 1872
rect 3710 1868 3714 1872
rect 3750 1868 3754 1872
rect 3798 1868 3802 1872
rect 3806 1868 3810 1872
rect 3830 1868 3834 1872
rect 3838 1868 3842 1872
rect 3886 1868 3890 1872
rect 3950 1878 3954 1882
rect 3982 1878 3986 1882
rect 4182 1878 4186 1882
rect 4190 1878 4194 1882
rect 4214 1878 4218 1882
rect 4294 1878 4298 1882
rect 4478 1878 4482 1882
rect 4486 1878 4490 1882
rect 4534 1878 4538 1882
rect 4542 1878 4546 1882
rect 4590 1878 4594 1882
rect 4846 1878 4850 1882
rect 4926 1878 4930 1882
rect 5014 1878 5018 1882
rect 5046 1878 5050 1882
rect 5278 1878 5282 1882
rect 3934 1868 3938 1872
rect 3966 1868 3970 1872
rect 4046 1868 4050 1872
rect 4094 1868 4098 1872
rect 4102 1868 4106 1872
rect 4174 1868 4178 1872
rect 4198 1868 4202 1872
rect 4214 1868 4218 1872
rect 4230 1868 4234 1872
rect 4286 1868 4290 1872
rect 4518 1868 4522 1872
rect 4534 1868 4538 1872
rect 4574 1868 4578 1872
rect 494 1858 498 1862
rect 502 1858 506 1862
rect 526 1858 530 1862
rect 550 1858 554 1862
rect 582 1858 586 1862
rect 606 1858 610 1862
rect 646 1858 650 1862
rect 670 1858 674 1862
rect 678 1858 682 1862
rect 694 1858 698 1862
rect 718 1858 722 1862
rect 758 1858 762 1862
rect 806 1858 810 1862
rect 822 1858 826 1862
rect 846 1858 850 1862
rect 854 1858 858 1862
rect 902 1858 906 1862
rect 942 1858 946 1862
rect 1054 1858 1058 1862
rect 1062 1858 1066 1862
rect 1078 1858 1082 1862
rect 1094 1858 1098 1862
rect 1102 1858 1106 1862
rect 1134 1858 1138 1862
rect 1150 1858 1154 1862
rect 1198 1858 1202 1862
rect 1270 1858 1274 1862
rect 1278 1858 1282 1862
rect 1310 1858 1314 1862
rect 1334 1858 1338 1862
rect 1390 1858 1394 1862
rect 1422 1858 1426 1862
rect 1470 1858 1474 1862
rect 1534 1858 1538 1862
rect 1558 1858 1562 1862
rect 1590 1858 1594 1862
rect 1606 1858 1610 1862
rect 1670 1858 1674 1862
rect 1742 1858 1746 1862
rect 1854 1858 1858 1862
rect 1942 1858 1946 1862
rect 1966 1858 1970 1862
rect 2006 1858 2010 1862
rect 2070 1858 2074 1862
rect 2134 1858 2138 1862
rect 2182 1858 2186 1862
rect 2230 1858 2234 1862
rect 2238 1858 2242 1862
rect 2406 1858 2410 1862
rect 2438 1858 2442 1862
rect 2534 1858 2538 1862
rect 2598 1858 2602 1862
rect 2670 1858 2674 1862
rect 2702 1858 2706 1862
rect 2766 1858 2770 1862
rect 2822 1858 2826 1862
rect 2830 1858 2834 1862
rect 2878 1858 2882 1862
rect 2942 1858 2946 1862
rect 2990 1858 2994 1862
rect 2998 1858 3002 1862
rect 3006 1858 3010 1862
rect 3038 1858 3042 1862
rect 3054 1858 3058 1862
rect 3118 1858 3122 1862
rect 3134 1858 3138 1862
rect 3150 1858 3154 1862
rect 3182 1858 3186 1862
rect 3190 1858 3194 1862
rect 3214 1858 3218 1862
rect 3230 1858 3234 1862
rect 3262 1858 3266 1862
rect 3278 1858 3282 1862
rect 3326 1858 3330 1862
rect 3382 1858 3386 1862
rect 3438 1858 3442 1862
rect 3486 1858 3490 1862
rect 3526 1858 3530 1862
rect 3590 1858 3594 1862
rect 3670 1858 3674 1862
rect 3678 1858 3682 1862
rect 3694 1858 3698 1862
rect 3726 1858 3730 1862
rect 3790 1858 3794 1862
rect 3830 1858 3834 1862
rect 3846 1858 3850 1862
rect 3910 1858 3914 1862
rect 3926 1858 3930 1862
rect 3958 1858 3962 1862
rect 3990 1858 3994 1862
rect 4014 1858 4018 1862
rect 4038 1858 4042 1862
rect 4054 1858 4058 1862
rect 4110 1858 4114 1862
rect 4166 1858 4170 1862
rect 4206 1858 4210 1862
rect 4238 1858 4242 1862
rect 4246 1858 4250 1862
rect 4254 1858 4258 1862
rect 4342 1858 4346 1862
rect 4366 1858 4370 1862
rect 4406 1858 4410 1862
rect 4414 1858 4418 1862
rect 4502 1858 4506 1862
rect 4510 1858 4514 1862
rect 4558 1858 4562 1862
rect 4566 1858 4570 1862
rect 4582 1858 4586 1862
rect 4614 1858 4618 1862
rect 4630 1868 4634 1872
rect 4758 1868 4762 1872
rect 4806 1868 4810 1872
rect 4814 1868 4818 1872
rect 4870 1868 4874 1872
rect 4950 1868 4954 1872
rect 4966 1868 4970 1872
rect 5006 1868 5010 1872
rect 5030 1868 5034 1872
rect 5062 1868 5066 1872
rect 5166 1868 5170 1872
rect 4630 1858 4634 1862
rect 4638 1858 4642 1862
rect 4694 1858 4698 1862
rect 4710 1858 4714 1862
rect 4758 1858 4762 1862
rect 4870 1858 4874 1862
rect 4894 1858 4898 1862
rect 4910 1858 4914 1862
rect 4958 1858 4962 1862
rect 5006 1858 5010 1862
rect 5038 1858 5042 1862
rect 5094 1858 5098 1862
rect 5102 1858 5106 1862
rect 5118 1858 5122 1862
rect 5142 1858 5146 1862
rect 5166 1858 5170 1862
rect 5182 1858 5186 1862
rect 5206 1858 5210 1862
rect 5222 1858 5226 1862
rect 5230 1858 5234 1862
rect 566 1848 570 1852
rect 598 1848 602 1852
rect 710 1848 714 1852
rect 782 1848 786 1852
rect 1094 1848 1098 1852
rect 1134 1848 1138 1852
rect 1350 1848 1354 1852
rect 1374 1848 1378 1852
rect 1406 1848 1410 1852
rect 1710 1848 1714 1852
rect 2038 1848 2042 1852
rect 2198 1848 2202 1852
rect 2366 1848 2370 1852
rect 2550 1848 2554 1852
rect 2558 1848 2562 1852
rect 2606 1848 2610 1852
rect 2630 1848 2634 1852
rect 2678 1848 2682 1852
rect 2710 1848 2714 1852
rect 2846 1848 2850 1852
rect 3022 1848 3026 1852
rect 3054 1848 3058 1852
rect 3094 1848 3098 1852
rect 3174 1848 3178 1852
rect 3454 1848 3458 1852
rect 3710 1848 3714 1852
rect 3718 1848 3722 1852
rect 3766 1848 3770 1852
rect 3806 1848 3810 1852
rect 3870 1848 3874 1852
rect 3982 1848 3986 1852
rect 4022 1848 4026 1852
rect 4150 1848 4154 1852
rect 4598 1848 4602 1852
rect 4654 1848 4658 1852
rect 4790 1848 4794 1852
rect 4878 1848 4882 1852
rect 4974 1848 4978 1852
rect 4982 1848 4986 1852
rect 1238 1838 1242 1842
rect 1254 1838 1258 1842
rect 1294 1838 1298 1842
rect 1510 1838 1514 1842
rect 1814 1838 1818 1842
rect 2438 1838 2442 1842
rect 2542 1838 2546 1842
rect 2590 1838 2594 1842
rect 2662 1838 2666 1842
rect 2694 1838 2698 1842
rect 3566 1838 3570 1842
rect 3734 1838 3738 1842
rect 4614 1838 4618 1842
rect 4766 1838 4770 1842
rect 654 1818 658 1822
rect 742 1818 746 1822
rect 1334 1818 1338 1822
rect 1798 1818 1802 1822
rect 1998 1818 2002 1822
rect 2406 1818 2410 1822
rect 2542 1818 2546 1822
rect 2598 1818 2602 1822
rect 2622 1818 2626 1822
rect 2670 1818 2674 1822
rect 2702 1818 2706 1822
rect 3470 1818 3474 1822
rect 3726 1818 3730 1822
rect 4006 1818 4010 1822
rect 4638 1818 4642 1822
rect 5014 1818 5018 1822
rect 330 1803 334 1807
rect 337 1803 341 1807
rect 1354 1803 1358 1807
rect 1361 1803 1365 1807
rect 2386 1803 2390 1807
rect 2393 1803 2397 1807
rect 3402 1803 3406 1807
rect 3409 1803 3413 1807
rect 4426 1803 4430 1807
rect 4433 1803 4437 1807
rect 62 1788 66 1792
rect 238 1788 242 1792
rect 430 1788 434 1792
rect 710 1788 714 1792
rect 1542 1788 1546 1792
rect 1590 1788 1594 1792
rect 1990 1788 1994 1792
rect 2022 1788 2026 1792
rect 2134 1788 2138 1792
rect 2222 1788 2226 1792
rect 2270 1788 2274 1792
rect 2326 1788 2330 1792
rect 2366 1788 2370 1792
rect 2486 1788 2490 1792
rect 2502 1788 2506 1792
rect 2550 1788 2554 1792
rect 2846 1788 2850 1792
rect 3126 1788 3130 1792
rect 3502 1788 3506 1792
rect 3910 1788 3914 1792
rect 4342 1788 4346 1792
rect 4678 1788 4682 1792
rect 4982 1788 4986 1792
rect 5054 1788 5058 1792
rect 2166 1778 2170 1782
rect 2966 1778 2970 1782
rect 4278 1778 4282 1782
rect 1070 1768 1074 1772
rect 1110 1768 1114 1772
rect 2070 1768 2074 1772
rect 2766 1768 2770 1772
rect 3438 1768 3442 1772
rect 4006 1768 4010 1772
rect 4590 1768 4594 1772
rect 374 1758 378 1762
rect 414 1758 418 1762
rect 190 1748 194 1752
rect 278 1748 282 1752
rect 374 1748 378 1752
rect 430 1748 434 1752
rect 454 1758 458 1762
rect 582 1758 586 1762
rect 598 1758 602 1762
rect 742 1758 746 1762
rect 918 1758 922 1762
rect 950 1758 954 1762
rect 510 1748 514 1752
rect 6 1738 10 1742
rect 78 1738 82 1742
rect 142 1738 146 1742
rect 158 1738 162 1742
rect 254 1738 258 1742
rect 542 1747 546 1751
rect 582 1748 586 1752
rect 654 1748 658 1752
rect 726 1748 730 1752
rect 750 1748 754 1752
rect 782 1748 786 1752
rect 798 1748 802 1752
rect 846 1747 850 1751
rect 966 1748 970 1752
rect 1014 1748 1018 1752
rect 1038 1748 1042 1752
rect 1086 1748 1090 1752
rect 1094 1748 1098 1752
rect 1334 1758 1338 1762
rect 1126 1748 1130 1752
rect 1142 1748 1146 1752
rect 1174 1748 1178 1752
rect 1206 1748 1210 1752
rect 1262 1748 1266 1752
rect 1334 1748 1338 1752
rect 1374 1758 1378 1762
rect 1526 1758 1530 1762
rect 1694 1758 1698 1762
rect 1718 1758 1722 1762
rect 1750 1758 1754 1762
rect 1798 1758 1802 1762
rect 1918 1758 1922 1762
rect 2006 1758 2010 1762
rect 2038 1758 2042 1762
rect 2054 1758 2058 1762
rect 2078 1758 2082 1762
rect 2614 1758 2618 1762
rect 2646 1758 2650 1762
rect 2798 1758 2802 1762
rect 2830 1758 2834 1762
rect 2854 1758 2858 1762
rect 1398 1748 1402 1752
rect 1422 1748 1426 1752
rect 1462 1748 1466 1752
rect 1478 1748 1482 1752
rect 1542 1748 1546 1752
rect 1558 1748 1562 1752
rect 1726 1748 1730 1752
rect 1734 1748 1738 1752
rect 1782 1748 1786 1752
rect 398 1738 402 1742
rect 422 1738 426 1742
rect 558 1738 562 1742
rect 574 1738 578 1742
rect 614 1738 618 1742
rect 662 1738 666 1742
rect 718 1738 722 1742
rect 806 1738 810 1742
rect 830 1738 834 1742
rect 926 1738 930 1742
rect 942 1738 946 1742
rect 974 1738 978 1742
rect 990 1738 994 1742
rect 1078 1738 1082 1742
rect 1134 1738 1138 1742
rect 1158 1738 1162 1742
rect 1182 1738 1186 1742
rect 1222 1738 1226 1742
rect 1238 1738 1242 1742
rect 1326 1738 1330 1742
rect 1398 1738 1402 1742
rect 1550 1738 1554 1742
rect 1574 1738 1578 1742
rect 1622 1738 1626 1742
rect 1654 1738 1658 1742
rect 1710 1738 1714 1742
rect 1742 1738 1746 1742
rect 1766 1738 1770 1742
rect 1830 1747 1834 1751
rect 1910 1748 1914 1752
rect 1934 1748 1938 1752
rect 1974 1748 1978 1752
rect 1990 1748 1994 1752
rect 2022 1748 2026 1752
rect 2046 1748 2050 1752
rect 2094 1748 2098 1752
rect 2110 1748 2114 1752
rect 2118 1748 2122 1752
rect 2142 1748 2146 1752
rect 2158 1748 2162 1752
rect 2206 1748 2210 1752
rect 2254 1748 2258 1752
rect 2310 1748 2314 1752
rect 2342 1748 2346 1752
rect 2422 1747 2426 1751
rect 2502 1748 2506 1752
rect 2518 1748 2522 1752
rect 2534 1748 2538 1752
rect 2590 1748 2594 1752
rect 2630 1748 2634 1752
rect 2638 1748 2642 1752
rect 2678 1747 2682 1751
rect 2710 1748 2714 1752
rect 2766 1748 2770 1752
rect 2814 1748 2818 1752
rect 2910 1748 2914 1752
rect 2982 1748 2986 1752
rect 2990 1748 2994 1752
rect 3006 1758 3010 1762
rect 3038 1758 3042 1762
rect 3190 1758 3194 1762
rect 3022 1748 3026 1752
rect 3054 1748 3058 1752
rect 3070 1748 3074 1752
rect 3102 1748 3106 1752
rect 3134 1748 3138 1752
rect 3142 1748 3146 1752
rect 3166 1748 3170 1752
rect 3238 1748 3242 1752
rect 3302 1748 3306 1752
rect 3326 1758 3330 1762
rect 3486 1758 3490 1762
rect 3518 1758 3522 1762
rect 3894 1758 3898 1762
rect 4230 1758 4234 1762
rect 4254 1758 4258 1762
rect 3374 1747 3378 1751
rect 3470 1748 3474 1752
rect 3502 1748 3506 1752
rect 3518 1748 3522 1752
rect 3550 1748 3554 1752
rect 3558 1748 3562 1752
rect 3646 1748 3650 1752
rect 3670 1748 3674 1752
rect 3750 1748 3754 1752
rect 3830 1748 3834 1752
rect 3854 1748 3858 1752
rect 3862 1748 3866 1752
rect 3878 1748 3882 1752
rect 3894 1748 3898 1752
rect 3918 1748 3922 1752
rect 3950 1748 3954 1752
rect 3974 1748 3978 1752
rect 3982 1748 3986 1752
rect 3990 1748 3994 1752
rect 4062 1748 4066 1752
rect 4166 1748 4170 1752
rect 4174 1748 4178 1752
rect 4182 1748 4186 1752
rect 4198 1748 4202 1752
rect 4214 1748 4218 1752
rect 4318 1758 4322 1762
rect 4366 1758 4370 1762
rect 4534 1758 4538 1762
rect 4694 1758 4698 1762
rect 4846 1758 4850 1762
rect 4278 1748 4282 1752
rect 4302 1748 4306 1752
rect 4334 1748 4338 1752
rect 4382 1748 4386 1752
rect 1798 1738 1802 1742
rect 1814 1738 1818 1742
rect 1942 1738 1946 1742
rect 1966 1738 1970 1742
rect 1982 1738 1986 1742
rect 2014 1738 2018 1742
rect 2046 1738 2050 1742
rect 2086 1738 2090 1742
rect 2102 1738 2106 1742
rect 2214 1738 2218 1742
rect 2390 1738 2394 1742
rect 2494 1738 2498 1742
rect 2526 1738 2530 1742
rect 2598 1738 2602 1742
rect 2774 1738 2778 1742
rect 2782 1738 2786 1742
rect 2806 1738 2810 1742
rect 2838 1738 2842 1742
rect 2918 1738 2922 1742
rect 2974 1738 2978 1742
rect 3030 1738 3034 1742
rect 3046 1738 3050 1742
rect 3062 1738 3066 1742
rect 3070 1738 3074 1742
rect 3094 1738 3098 1742
rect 3110 1738 3114 1742
rect 3166 1738 3170 1742
rect 3254 1738 3258 1742
rect 3294 1738 3298 1742
rect 3318 1738 3322 1742
rect 3342 1738 3346 1742
rect 3358 1738 3362 1742
rect 3462 1738 3466 1742
rect 3542 1738 3546 1742
rect 3590 1738 3594 1742
rect 3606 1738 3610 1742
rect 3742 1738 3746 1742
rect 3830 1738 3834 1742
rect 3870 1738 3874 1742
rect 3934 1738 3938 1742
rect 4030 1738 4034 1742
rect 4118 1738 4122 1742
rect 4142 1738 4146 1742
rect 4438 1747 4442 1751
rect 4510 1748 4514 1752
rect 4518 1748 4522 1752
rect 4542 1748 4546 1752
rect 4614 1748 4618 1752
rect 4678 1748 4682 1752
rect 4694 1748 4698 1752
rect 4718 1748 4722 1752
rect 4734 1748 4738 1752
rect 4974 1758 4978 1762
rect 4798 1747 4802 1751
rect 4870 1748 4874 1752
rect 5014 1748 5018 1752
rect 5046 1748 5050 1752
rect 5070 1748 5074 1752
rect 5078 1748 5082 1752
rect 5174 1748 5178 1752
rect 4206 1738 4210 1742
rect 4238 1738 4242 1742
rect 4286 1738 4290 1742
rect 4294 1738 4298 1742
rect 4358 1738 4362 1742
rect 4390 1738 4394 1742
rect 4406 1738 4410 1742
rect 4446 1738 4450 1742
rect 4614 1738 4618 1742
rect 4654 1738 4658 1742
rect 4670 1738 4674 1742
rect 4726 1738 4730 1742
rect 4814 1738 4818 1742
rect 4830 1738 4834 1742
rect 4854 1738 4858 1742
rect 4878 1738 4882 1742
rect 4886 1738 4890 1742
rect 4950 1738 4954 1742
rect 5038 1738 5042 1742
rect 5102 1738 5106 1742
rect 5214 1738 5218 1742
rect 5230 1738 5234 1742
rect 5294 1738 5298 1742
rect 206 1728 210 1732
rect 342 1728 346 1732
rect 750 1728 754 1732
rect 766 1728 770 1732
rect 1406 1728 1410 1732
rect 1422 1728 1426 1732
rect 1678 1728 1682 1732
rect 1950 1728 1954 1732
rect 1958 1728 1962 1732
rect 2174 1728 2178 1732
rect 2574 1728 2578 1732
rect 2742 1728 2746 1732
rect 2830 1728 2834 1732
rect 3094 1728 3098 1732
rect 3126 1728 3130 1732
rect 3526 1728 3530 1732
rect 3902 1728 3906 1732
rect 4198 1728 4202 1732
rect 4470 1728 4474 1732
rect 4998 1728 5002 1732
rect 5062 1728 5066 1732
rect 5126 1728 5130 1732
rect 334 1718 338 1722
rect 382 1718 386 1722
rect 406 1718 410 1722
rect 478 1718 482 1722
rect 910 1718 914 1722
rect 1190 1718 1194 1722
rect 1318 1718 1322 1722
rect 1430 1718 1434 1722
rect 1558 1718 1562 1722
rect 1630 1718 1634 1722
rect 1702 1718 1706 1722
rect 1750 1718 1754 1722
rect 2294 1718 2298 1722
rect 2606 1718 2610 1722
rect 2798 1718 2802 1722
rect 4230 1718 4234 1722
rect 5030 1718 5034 1722
rect 850 1703 854 1707
rect 857 1703 861 1707
rect 1874 1703 1878 1707
rect 1881 1703 1885 1707
rect 2890 1703 2894 1707
rect 2897 1703 2901 1707
rect 3922 1703 3926 1707
rect 3929 1703 3933 1707
rect 4938 1703 4942 1707
rect 4945 1703 4949 1707
rect 94 1688 98 1692
rect 190 1688 194 1692
rect 334 1688 338 1692
rect 358 1688 362 1692
rect 518 1688 522 1692
rect 526 1688 530 1692
rect 742 1688 746 1692
rect 902 1688 906 1692
rect 1014 1688 1018 1692
rect 1286 1688 1290 1692
rect 1326 1688 1330 1692
rect 1478 1688 1482 1692
rect 1686 1688 1690 1692
rect 1766 1688 1770 1692
rect 1918 1688 1922 1692
rect 1958 1688 1962 1692
rect 2014 1688 2018 1692
rect 2046 1688 2050 1692
rect 2078 1688 2082 1692
rect 2230 1688 2234 1692
rect 2286 1688 2290 1692
rect 2390 1688 2394 1692
rect 2830 1688 2834 1692
rect 3102 1688 3106 1692
rect 3198 1688 3202 1692
rect 3366 1688 3370 1692
rect 3390 1688 3394 1692
rect 3486 1688 3490 1692
rect 3598 1688 3602 1692
rect 3638 1688 3642 1692
rect 3822 1688 3826 1692
rect 4134 1688 4138 1692
rect 4270 1688 4274 1692
rect 4318 1688 4322 1692
rect 5206 1688 5210 1692
rect 5270 1688 5274 1692
rect 390 1678 394 1682
rect 894 1678 898 1682
rect 1142 1678 1146 1682
rect 1182 1678 1186 1682
rect 1254 1678 1258 1682
rect 1294 1678 1298 1682
rect 1422 1678 1426 1682
rect 1438 1678 1442 1682
rect 1726 1678 1730 1682
rect 1966 1678 1970 1682
rect 2086 1678 2090 1682
rect 14 1668 18 1672
rect 62 1668 66 1672
rect 102 1668 106 1672
rect 126 1668 130 1672
rect 158 1668 162 1672
rect 166 1668 170 1672
rect 222 1668 226 1672
rect 238 1668 242 1672
rect 334 1668 338 1672
rect 398 1668 402 1672
rect 438 1668 442 1672
rect 542 1666 546 1670
rect 550 1668 554 1672
rect 558 1668 562 1672
rect 598 1668 602 1672
rect 614 1668 618 1672
rect 646 1668 650 1672
rect 662 1668 666 1672
rect 750 1668 754 1672
rect 814 1668 818 1672
rect 870 1668 874 1672
rect 894 1668 898 1672
rect 942 1668 946 1672
rect 46 1658 50 1662
rect 118 1658 122 1662
rect 142 1658 146 1662
rect 150 1658 154 1662
rect 174 1658 178 1662
rect 214 1658 218 1662
rect 254 1659 258 1663
rect 342 1658 346 1662
rect 374 1658 378 1662
rect 398 1658 402 1662
rect 462 1658 466 1662
rect 582 1658 586 1662
rect 606 1658 610 1662
rect 646 1658 650 1662
rect 686 1658 690 1662
rect 758 1658 762 1662
rect 798 1658 802 1662
rect 878 1658 882 1662
rect 910 1658 914 1662
rect 950 1658 954 1662
rect 1046 1658 1050 1662
rect 1078 1659 1082 1663
rect 1142 1668 1146 1672
rect 1270 1668 1274 1672
rect 1302 1668 1306 1672
rect 1334 1668 1338 1672
rect 1366 1668 1370 1672
rect 1390 1668 1394 1672
rect 1406 1668 1410 1672
rect 1486 1668 1490 1672
rect 1510 1668 1514 1672
rect 1582 1668 1586 1672
rect 1662 1668 1666 1672
rect 1718 1668 1722 1672
rect 1814 1668 1818 1672
rect 1974 1668 1978 1672
rect 2022 1668 2026 1672
rect 2038 1668 2042 1672
rect 2070 1668 2074 1672
rect 2166 1678 2170 1682
rect 2694 1678 2698 1682
rect 2758 1678 2762 1682
rect 2822 1678 2826 1682
rect 2878 1678 2882 1682
rect 2974 1678 2978 1682
rect 2446 1668 2450 1672
rect 2510 1668 2514 1672
rect 2614 1668 2618 1672
rect 2654 1668 2658 1672
rect 2662 1668 2666 1672
rect 2710 1668 2714 1672
rect 2798 1668 2802 1672
rect 2838 1668 2842 1672
rect 2854 1668 2858 1672
rect 2934 1668 2938 1672
rect 3022 1668 3026 1672
rect 3046 1668 3050 1672
rect 3070 1678 3074 1682
rect 3118 1678 3122 1682
rect 3206 1678 3210 1682
rect 3270 1678 3274 1682
rect 3334 1678 3338 1682
rect 3566 1678 3570 1682
rect 3646 1678 3650 1682
rect 3710 1678 3714 1682
rect 3742 1678 3746 1682
rect 4070 1678 4074 1682
rect 4254 1678 4258 1682
rect 4302 1678 4306 1682
rect 3094 1668 3098 1672
rect 3142 1668 3146 1672
rect 3150 1668 3154 1672
rect 3206 1668 3210 1672
rect 3222 1668 3226 1672
rect 3374 1668 3378 1672
rect 3422 1668 3426 1672
rect 3478 1668 3482 1672
rect 3614 1668 3618 1672
rect 3630 1668 3634 1672
rect 3830 1668 3834 1672
rect 4014 1668 4018 1672
rect 4038 1668 4042 1672
rect 4166 1668 4170 1672
rect 4190 1668 4194 1672
rect 4222 1668 4226 1672
rect 4238 1668 4242 1672
rect 4254 1668 4258 1672
rect 4262 1668 4266 1672
rect 4374 1678 4378 1682
rect 4406 1678 4410 1682
rect 4614 1678 4618 1682
rect 4662 1678 4666 1682
rect 4326 1668 4330 1672
rect 4478 1668 4482 1672
rect 4518 1668 4522 1672
rect 4918 1678 4922 1682
rect 4998 1678 5002 1682
rect 5150 1678 5154 1682
rect 5238 1678 5242 1682
rect 5254 1678 5258 1682
rect 5278 1678 5282 1682
rect 4686 1668 4690 1672
rect 4726 1668 4730 1672
rect 4774 1668 4778 1672
rect 4782 1668 4786 1672
rect 4862 1668 4866 1672
rect 4902 1668 4906 1672
rect 5022 1668 5026 1672
rect 5078 1668 5082 1672
rect 1110 1658 1114 1662
rect 1126 1658 1130 1662
rect 1190 1658 1194 1662
rect 1270 1658 1274 1662
rect 1278 1658 1282 1662
rect 1310 1658 1314 1662
rect 1342 1658 1346 1662
rect 1358 1658 1362 1662
rect 1374 1658 1378 1662
rect 1422 1658 1426 1662
rect 1462 1658 1466 1662
rect 1494 1658 1498 1662
rect 1582 1659 1586 1663
rect 1622 1658 1626 1662
rect 1630 1658 1634 1662
rect 1646 1658 1650 1662
rect 1662 1658 1666 1662
rect 1670 1658 1674 1662
rect 1710 1658 1714 1662
rect 1750 1658 1754 1662
rect 1806 1658 1810 1662
rect 1910 1658 1914 1662
rect 1934 1658 1938 1662
rect 1942 1658 1946 1662
rect 1950 1658 1954 1662
rect 1974 1658 1978 1662
rect 2030 1658 2034 1662
rect 2062 1658 2066 1662
rect 2118 1658 2122 1662
rect 2126 1658 2130 1662
rect 2174 1658 2178 1662
rect 2270 1658 2274 1662
rect 2294 1658 2298 1662
rect 2334 1658 2338 1662
rect 2454 1658 2458 1662
rect 2486 1658 2490 1662
rect 2494 1658 2498 1662
rect 2526 1659 2530 1663
rect 2598 1658 2602 1662
rect 2622 1658 2626 1662
rect 2646 1658 2650 1662
rect 2678 1658 2682 1662
rect 2726 1659 2730 1663
rect 2814 1658 2818 1662
rect 2846 1658 2850 1662
rect 2862 1658 2866 1662
rect 2878 1658 2882 1662
rect 3006 1659 3010 1663
rect 3038 1658 3042 1662
rect 3054 1658 3058 1662
rect 3086 1658 3090 1662
rect 3134 1658 3138 1662
rect 3158 1658 3162 1662
rect 3230 1658 3234 1662
rect 3270 1658 3274 1662
rect 3302 1659 3306 1663
rect 3350 1658 3354 1662
rect 3382 1658 3386 1662
rect 3406 1658 3410 1662
rect 3414 1658 3418 1662
rect 3446 1658 3450 1662
rect 3558 1658 3562 1662
rect 3622 1658 3626 1662
rect 3654 1658 3658 1662
rect 3662 1658 3666 1662
rect 3694 1658 3698 1662
rect 3710 1658 3714 1662
rect 3750 1658 3754 1662
rect 3862 1658 3866 1662
rect 3870 1658 3874 1662
rect 3934 1658 3938 1662
rect 3950 1658 3954 1662
rect 4030 1658 4034 1662
rect 4094 1658 4098 1662
rect 4182 1658 4186 1662
rect 4198 1658 4202 1662
rect 4230 1658 4234 1662
rect 4286 1658 4290 1662
rect 4334 1658 4338 1662
rect 4406 1659 4410 1663
rect 4470 1658 4474 1662
rect 4486 1658 4490 1662
rect 4494 1658 4498 1662
rect 4526 1658 4530 1662
rect 4590 1658 4594 1662
rect 4646 1658 4650 1662
rect 4686 1658 4690 1662
rect 4718 1658 4722 1662
rect 4758 1658 4762 1662
rect 4766 1658 4770 1662
rect 4822 1658 4826 1662
rect 4878 1658 4882 1662
rect 4894 1658 4898 1662
rect 4974 1658 4978 1662
rect 4982 1658 4986 1662
rect 5030 1658 5034 1662
rect 5062 1658 5066 1662
rect 5070 1658 5074 1662
rect 5078 1658 5082 1662
rect 5126 1658 5130 1662
rect 5182 1658 5186 1662
rect 5190 1658 5194 1662
rect 5214 1658 5218 1662
rect 5262 1658 5266 1662
rect 102 1648 106 1652
rect 134 1648 138 1652
rect 198 1648 202 1652
rect 422 1648 426 1652
rect 590 1648 594 1652
rect 622 1648 626 1652
rect 782 1648 786 1652
rect 838 1648 842 1652
rect 1110 1648 1114 1652
rect 1414 1648 1418 1652
rect 1686 1648 1690 1652
rect 1694 1648 1698 1652
rect 1710 1648 1714 1652
rect 1766 1648 1770 1652
rect 1886 1648 1890 1652
rect 1998 1648 2002 1652
rect 2094 1648 2098 1652
rect 2470 1648 2474 1652
rect 2638 1648 2642 1652
rect 2902 1648 2906 1652
rect 3110 1648 3114 1652
rect 3118 1648 3122 1652
rect 3174 1648 3178 1652
rect 3198 1648 3202 1652
rect 3390 1648 3394 1652
rect 3598 1648 3602 1652
rect 4006 1648 4010 1652
rect 4158 1648 4162 1652
rect 4278 1648 4282 1652
rect 4454 1648 4458 1652
rect 4742 1648 4746 1652
rect 4878 1648 4882 1652
rect 5046 1648 5050 1652
rect 5238 1648 5242 1652
rect 726 1638 730 1642
rect 1006 1638 1010 1642
rect 1846 1638 1850 1642
rect 2110 1638 2114 1642
rect 2574 1638 2578 1642
rect 2958 1638 2962 1642
rect 3966 1638 3970 1642
rect 758 1628 762 1632
rect 2622 1628 2626 1632
rect 318 1618 322 1622
rect 406 1618 410 1622
rect 638 1618 642 1622
rect 1014 1618 1018 1622
rect 1150 1618 1154 1622
rect 1342 1618 1346 1622
rect 2134 1618 2138 1622
rect 2246 1618 2250 1622
rect 2286 1618 2290 1622
rect 2318 1618 2322 1622
rect 2350 1618 2354 1622
rect 3678 1618 3682 1622
rect 3982 1618 3986 1622
rect 4470 1618 4474 1622
rect 4702 1618 4706 1622
rect 5230 1618 5234 1622
rect 330 1603 334 1607
rect 337 1603 341 1607
rect 1354 1603 1358 1607
rect 1361 1603 1365 1607
rect 2386 1603 2390 1607
rect 2393 1603 2397 1607
rect 3402 1603 3406 1607
rect 3409 1603 3413 1607
rect 4426 1603 4430 1607
rect 4433 1603 4437 1607
rect 190 1588 194 1592
rect 222 1588 226 1592
rect 438 1588 442 1592
rect 574 1588 578 1592
rect 622 1588 626 1592
rect 686 1588 690 1592
rect 838 1588 842 1592
rect 958 1588 962 1592
rect 1102 1588 1106 1592
rect 1126 1588 1130 1592
rect 1406 1588 1410 1592
rect 1446 1588 1450 1592
rect 1678 1588 1682 1592
rect 1694 1588 1698 1592
rect 1894 1588 1898 1592
rect 2006 1588 2010 1592
rect 2174 1588 2178 1592
rect 2278 1588 2282 1592
rect 2846 1588 2850 1592
rect 2998 1588 3002 1592
rect 3214 1588 3218 1592
rect 3230 1588 3234 1592
rect 3334 1588 3338 1592
rect 3598 1588 3602 1592
rect 3670 1588 3674 1592
rect 3742 1588 3746 1592
rect 3854 1588 3858 1592
rect 4038 1588 4042 1592
rect 4126 1588 4130 1592
rect 4190 1588 4194 1592
rect 4286 1588 4290 1592
rect 4334 1588 4338 1592
rect 5030 1588 5034 1592
rect 5094 1588 5098 1592
rect 2390 1578 2394 1582
rect 2878 1578 2882 1582
rect 94 1568 98 1572
rect 270 1568 274 1572
rect 942 1568 946 1572
rect 1086 1568 1090 1572
rect 1134 1568 1138 1572
rect 1166 1568 1170 1572
rect 2502 1568 2506 1572
rect 2958 1568 2962 1572
rect 3110 1568 3114 1572
rect 3238 1568 3242 1572
rect 4406 1568 4410 1572
rect 4702 1568 4706 1572
rect 4926 1568 4930 1572
rect 102 1558 106 1562
rect 134 1558 138 1562
rect 238 1558 242 1562
rect 254 1558 258 1562
rect 414 1558 418 1562
rect 422 1558 426 1562
rect 606 1558 610 1562
rect 638 1558 642 1562
rect 670 1558 674 1562
rect 1118 1558 1122 1562
rect 1150 1558 1154 1562
rect 1310 1558 1314 1562
rect 1390 1558 1394 1562
rect 1494 1558 1498 1562
rect 1502 1558 1506 1562
rect 1550 1558 1554 1562
rect 38 1548 42 1552
rect 118 1548 122 1552
rect 134 1548 138 1552
rect 150 1548 154 1552
rect 206 1548 210 1552
rect 222 1548 226 1552
rect 254 1548 258 1552
rect 310 1548 314 1552
rect 326 1548 330 1552
rect 342 1548 346 1552
rect 374 1548 378 1552
rect 382 1548 386 1552
rect 398 1548 402 1552
rect 438 1548 442 1552
rect 478 1548 482 1552
rect 518 1548 522 1552
rect 590 1548 594 1552
rect 598 1548 602 1552
rect 622 1548 626 1552
rect 654 1548 658 1552
rect 662 1548 666 1552
rect 702 1548 706 1552
rect 758 1548 762 1552
rect 822 1548 826 1552
rect 902 1548 906 1552
rect 982 1548 986 1552
rect 1014 1548 1018 1552
rect 1046 1548 1050 1552
rect 1054 1548 1058 1552
rect 1102 1548 1106 1552
rect 1126 1548 1130 1552
rect 1166 1548 1170 1552
rect 1182 1548 1186 1552
rect 1246 1548 1250 1552
rect 1326 1548 1330 1552
rect 1334 1548 1338 1552
rect 1358 1548 1362 1552
rect 1366 1548 1370 1552
rect 1406 1548 1410 1552
rect 1430 1548 1434 1552
rect 1454 1548 1458 1552
rect 1462 1548 1466 1552
rect 1478 1548 1482 1552
rect 1534 1548 1538 1552
rect 1574 1558 1578 1562
rect 1718 1558 1722 1562
rect 1734 1558 1738 1562
rect 1766 1558 1770 1562
rect 1782 1558 1786 1562
rect 1798 1558 1802 1562
rect 1918 1558 1922 1562
rect 1958 1558 1962 1562
rect 1990 1558 1994 1562
rect 2022 1558 2026 1562
rect 2422 1558 2426 1562
rect 1574 1548 1578 1552
rect 1622 1548 1626 1552
rect 1718 1548 1722 1552
rect 1750 1548 1754 1552
rect 1766 1548 1770 1552
rect 1782 1548 1786 1552
rect 1838 1548 1842 1552
rect 1966 1548 1970 1552
rect 2030 1548 2034 1552
rect 2046 1548 2050 1552
rect 14 1538 18 1542
rect 102 1538 106 1542
rect 126 1538 130 1542
rect 158 1538 162 1542
rect 214 1538 218 1542
rect 246 1538 250 1542
rect 278 1538 282 1542
rect 326 1538 330 1542
rect 390 1538 394 1542
rect 446 1538 450 1542
rect 510 1538 514 1542
rect 582 1538 586 1542
rect 614 1538 618 1542
rect 646 1538 650 1542
rect 718 1538 722 1542
rect 878 1538 882 1542
rect 990 1538 994 1542
rect 1014 1538 1018 1542
rect 1078 1538 1082 1542
rect 1110 1538 1114 1542
rect 1174 1538 1178 1542
rect 1206 1538 1210 1542
rect 1222 1538 1226 1542
rect 1414 1538 1418 1542
rect 1470 1538 1474 1542
rect 1518 1538 1522 1542
rect 1526 1538 1530 1542
rect 1582 1538 1586 1542
rect 1614 1538 1618 1542
rect 1622 1538 1626 1542
rect 1718 1538 1722 1542
rect 1742 1538 1746 1542
rect 1774 1538 1778 1542
rect 1846 1538 1850 1542
rect 1934 1538 1938 1542
rect 1966 1538 1970 1542
rect 1998 1538 2002 1542
rect 2078 1547 2082 1551
rect 2110 1548 2114 1552
rect 2150 1548 2154 1552
rect 2158 1548 2162 1552
rect 2182 1548 2186 1552
rect 2190 1548 2194 1552
rect 2254 1548 2258 1552
rect 2334 1548 2338 1552
rect 2350 1548 2354 1552
rect 2438 1548 2442 1552
rect 2446 1548 2450 1552
rect 2462 1558 2466 1562
rect 2486 1548 2490 1552
rect 2566 1558 2570 1562
rect 2550 1548 2554 1552
rect 2678 1558 2682 1562
rect 2822 1558 2826 1562
rect 2934 1558 2938 1562
rect 2974 1558 2978 1562
rect 3070 1558 3074 1562
rect 2582 1548 2586 1552
rect 2590 1548 2594 1552
rect 2630 1547 2634 1551
rect 2726 1547 2730 1551
rect 2806 1548 2810 1552
rect 2814 1548 2818 1552
rect 2846 1548 2850 1552
rect 2918 1548 2922 1552
rect 2942 1548 2946 1552
rect 3046 1548 3050 1552
rect 3222 1558 3226 1562
rect 3374 1558 3378 1562
rect 3518 1558 3522 1562
rect 3622 1558 3626 1562
rect 3654 1558 3658 1562
rect 4094 1558 4098 1562
rect 4166 1558 4170 1562
rect 4174 1558 4178 1562
rect 4222 1558 4226 1562
rect 4230 1558 4234 1562
rect 4382 1558 4386 1562
rect 4390 1558 4394 1562
rect 4438 1558 4442 1562
rect 4470 1558 4474 1562
rect 4550 1558 4554 1562
rect 4574 1558 4578 1562
rect 4638 1558 4642 1562
rect 4686 1558 4690 1562
rect 4822 1558 4826 1562
rect 4886 1558 4890 1562
rect 3094 1548 3098 1552
rect 3150 1548 3154 1552
rect 3230 1548 3234 1552
rect 3254 1548 3258 1552
rect 3286 1548 3290 1552
rect 3334 1548 3338 1552
rect 3430 1548 3434 1552
rect 3502 1548 3506 1552
rect 3526 1548 3530 1552
rect 3550 1548 3554 1552
rect 3574 1548 3578 1552
rect 3590 1548 3594 1552
rect 3606 1548 3610 1552
rect 3638 1548 3642 1552
rect 3686 1548 3690 1552
rect 3702 1548 3706 1552
rect 3734 1548 3738 1552
rect 3798 1548 3802 1552
rect 3838 1548 3842 1552
rect 3846 1548 3850 1552
rect 3870 1548 3874 1552
rect 3910 1548 3914 1552
rect 3982 1548 3986 1552
rect 4078 1548 4082 1552
rect 4086 1548 4090 1552
rect 4142 1548 4146 1552
rect 4150 1548 4154 1552
rect 4166 1548 4170 1552
rect 4190 1548 4194 1552
rect 4254 1548 4258 1552
rect 4286 1548 4290 1552
rect 4302 1548 4306 1552
rect 4318 1548 4322 1552
rect 4326 1548 4330 1552
rect 4350 1548 4354 1552
rect 4406 1548 4410 1552
rect 4414 1548 4418 1552
rect 4462 1548 4466 1552
rect 4494 1548 4498 1552
rect 4526 1548 4530 1552
rect 4534 1548 4538 1552
rect 4542 1548 4546 1552
rect 4550 1548 4554 1552
rect 4590 1548 4594 1552
rect 4606 1548 4610 1552
rect 4654 1548 4658 1552
rect 4662 1548 4666 1552
rect 4734 1548 4738 1552
rect 2286 1538 2290 1542
rect 2406 1538 2410 1542
rect 2430 1538 2434 1542
rect 2494 1538 2498 1542
rect 2534 1538 2538 1542
rect 2542 1538 2546 1542
rect 2598 1538 2602 1542
rect 2614 1538 2618 1542
rect 2662 1538 2666 1542
rect 2710 1538 2714 1542
rect 2798 1538 2802 1542
rect 2854 1538 2858 1542
rect 2902 1538 2906 1542
rect 2990 1538 2994 1542
rect 3014 1538 3018 1542
rect 3046 1538 3050 1542
rect 3086 1538 3090 1542
rect 3102 1538 3106 1542
rect 3190 1538 3194 1542
rect 3262 1538 3266 1542
rect 3358 1538 3362 1542
rect 3438 1538 3442 1542
rect 3494 1538 3498 1542
rect 3574 1538 3578 1542
rect 3582 1538 3586 1542
rect 3646 1538 3650 1542
rect 3678 1538 3682 1542
rect 3726 1538 3730 1542
rect 3822 1538 3826 1542
rect 3966 1538 3970 1542
rect 4054 1538 4058 1542
rect 4110 1538 4114 1542
rect 4134 1538 4138 1542
rect 4766 1547 4770 1551
rect 4806 1548 4810 1552
rect 4814 1548 4818 1552
rect 4830 1548 4834 1552
rect 4838 1548 4842 1552
rect 4846 1548 4850 1552
rect 4862 1548 4866 1552
rect 4902 1548 4906 1552
rect 4926 1548 4930 1552
rect 4974 1548 4978 1552
rect 5046 1548 5050 1552
rect 5054 1548 5058 1552
rect 5078 1548 5082 1552
rect 5142 1548 5146 1552
rect 5238 1548 5242 1552
rect 5262 1548 5266 1552
rect 4198 1538 4202 1542
rect 4206 1538 4210 1542
rect 4222 1538 4226 1542
rect 4246 1538 4250 1542
rect 4310 1538 4314 1542
rect 4366 1538 4370 1542
rect 4414 1538 4418 1542
rect 4462 1538 4466 1542
rect 4494 1538 4498 1542
rect 4526 1538 4530 1542
rect 4598 1538 4602 1542
rect 4614 1538 4618 1542
rect 4630 1538 4634 1542
rect 4662 1538 4666 1542
rect 4798 1538 4802 1542
rect 4854 1538 4858 1542
rect 4894 1538 4898 1542
rect 4910 1538 4914 1542
rect 5014 1538 5018 1542
rect 5086 1538 5090 1542
rect 5150 1538 5154 1542
rect 166 1528 170 1532
rect 310 1528 314 1532
rect 1494 1528 1498 1532
rect 2030 1528 2034 1532
rect 2790 1528 2794 1532
rect 2830 1528 2834 1532
rect 2934 1528 2938 1532
rect 2998 1528 3002 1532
rect 3038 1528 3042 1532
rect 3206 1528 3210 1532
rect 3302 1528 3306 1532
rect 3310 1528 3314 1532
rect 3558 1528 3562 1532
rect 3686 1528 3690 1532
rect 4118 1528 4122 1532
rect 4270 1528 4274 1532
rect 4502 1528 4506 1532
rect 4566 1528 4570 1532
rect 4630 1528 4634 1532
rect 4878 1528 4882 1532
rect 5038 1528 5042 1532
rect 5198 1528 5202 1532
rect 5270 1528 5274 1532
rect 174 1518 178 1522
rect 190 1518 194 1522
rect 414 1518 418 1522
rect 462 1518 466 1522
rect 574 1518 578 1522
rect 814 1518 818 1522
rect 838 1518 842 1522
rect 1030 1518 1034 1522
rect 1510 1518 1514 1522
rect 1734 1518 1738 1522
rect 1926 1518 1930 1522
rect 1958 1518 1962 1522
rect 2142 1518 2146 1522
rect 2214 1518 2218 1522
rect 2238 1518 2242 1522
rect 2414 1518 2418 1522
rect 2526 1518 2530 1522
rect 2694 1518 2698 1522
rect 2862 1518 2866 1522
rect 2974 1518 2978 1522
rect 3270 1518 3274 1522
rect 3486 1518 3490 1522
rect 3534 1518 3538 1522
rect 3718 1518 3722 1522
rect 3894 1518 3898 1522
rect 4094 1518 4098 1522
rect 4238 1518 4242 1522
rect 4382 1518 4386 1522
rect 4470 1518 4474 1522
rect 4510 1518 4514 1522
rect 4574 1518 4578 1522
rect 4622 1518 4626 1522
rect 4870 1518 4874 1522
rect 5190 1518 5194 1522
rect 5206 1518 5210 1522
rect 850 1503 854 1507
rect 857 1503 861 1507
rect 1874 1503 1878 1507
rect 1881 1503 1885 1507
rect 2890 1503 2894 1507
rect 2897 1503 2901 1507
rect 3922 1503 3926 1507
rect 3929 1503 3933 1507
rect 4938 1503 4942 1507
rect 4945 1503 4949 1507
rect 94 1488 98 1492
rect 294 1488 298 1492
rect 350 1488 354 1492
rect 478 1488 482 1492
rect 566 1488 570 1492
rect 606 1488 610 1492
rect 638 1488 642 1492
rect 734 1488 738 1492
rect 758 1488 762 1492
rect 822 1488 826 1492
rect 918 1488 922 1492
rect 1126 1488 1130 1492
rect 1390 1488 1394 1492
rect 1486 1488 1490 1492
rect 1590 1488 1594 1492
rect 1686 1488 1690 1492
rect 1798 1488 1802 1492
rect 1998 1488 2002 1492
rect 2046 1488 2050 1492
rect 2078 1488 2082 1492
rect 2118 1488 2122 1492
rect 2462 1488 2466 1492
rect 2486 1488 2490 1492
rect 2654 1488 2658 1492
rect 2710 1488 2714 1492
rect 2870 1488 2874 1492
rect 2934 1488 2938 1492
rect 3110 1488 3114 1492
rect 3294 1488 3298 1492
rect 3342 1488 3346 1492
rect 3470 1488 3474 1492
rect 3494 1488 3498 1492
rect 3686 1488 3690 1492
rect 3854 1488 3858 1492
rect 4054 1488 4058 1492
rect 4654 1488 4658 1492
rect 4862 1488 4866 1492
rect 4958 1488 4962 1492
rect 5078 1488 5082 1492
rect 198 1478 202 1482
rect 790 1478 794 1482
rect 926 1478 930 1482
rect 1294 1478 1298 1482
rect 1398 1478 1402 1482
rect 1478 1478 1482 1482
rect 1622 1478 1626 1482
rect 1694 1478 1698 1482
rect 1942 1478 1946 1482
rect 2182 1478 2186 1482
rect 2454 1478 2458 1482
rect 2558 1478 2562 1482
rect 2742 1478 2746 1482
rect 2942 1478 2946 1482
rect 3014 1478 3018 1482
rect 3326 1478 3330 1482
rect 14 1468 18 1472
rect 126 1468 130 1472
rect 142 1468 146 1472
rect 158 1468 162 1472
rect 166 1468 170 1472
rect 302 1468 306 1472
rect 374 1468 378 1472
rect 382 1468 386 1472
rect 438 1468 442 1472
rect 446 1468 450 1472
rect 502 1468 506 1472
rect 510 1468 514 1472
rect 582 1468 586 1472
rect 614 1468 618 1472
rect 654 1468 658 1472
rect 910 1468 914 1472
rect 942 1468 946 1472
rect 1094 1468 1098 1472
rect 1102 1468 1106 1472
rect 1142 1468 1146 1472
rect 1310 1468 1314 1472
rect 1326 1468 1330 1472
rect 1382 1468 1386 1472
rect 1462 1468 1466 1472
rect 1510 1468 1514 1472
rect 1566 1468 1570 1472
rect 1710 1468 1714 1472
rect 1726 1468 1730 1472
rect 1742 1468 1746 1472
rect 1782 1468 1786 1472
rect 1790 1468 1794 1472
rect 1822 1468 1826 1472
rect 1862 1468 1866 1472
rect 1918 1468 1922 1472
rect 1942 1468 1946 1472
rect 1958 1468 1962 1472
rect 2022 1468 2026 1472
rect 2054 1468 2058 1472
rect 2110 1468 2114 1472
rect 2222 1468 2226 1472
rect 2238 1468 2242 1472
rect 2270 1468 2274 1472
rect 2278 1468 2282 1472
rect 2302 1468 2306 1472
rect 2310 1468 2314 1472
rect 2350 1468 2354 1472
rect 2366 1468 2370 1472
rect 2518 1468 2522 1472
rect 2606 1468 2610 1472
rect 2702 1468 2706 1472
rect 2750 1468 2754 1472
rect 2910 1468 2914 1472
rect 2990 1468 2994 1472
rect 2998 1468 3002 1472
rect 3118 1468 3122 1472
rect 3174 1468 3178 1472
rect 3262 1468 3266 1472
rect 3526 1478 3530 1482
rect 3750 1478 3754 1482
rect 3990 1478 3994 1482
rect 4094 1478 4098 1482
rect 4238 1478 4242 1482
rect 4318 1478 4322 1482
rect 4382 1478 4386 1482
rect 4478 1478 4482 1482
rect 4822 1478 4826 1482
rect 4838 1478 4842 1482
rect 4870 1478 4874 1482
rect 5094 1478 5098 1482
rect 5118 1478 5122 1482
rect 5238 1478 5242 1482
rect 5270 1478 5274 1482
rect 3366 1468 3370 1472
rect 3478 1468 3482 1472
rect 3542 1468 3546 1472
rect 3630 1468 3634 1472
rect 3654 1468 3658 1472
rect 3678 1468 3682 1472
rect 3782 1468 3786 1472
rect 3814 1468 3818 1472
rect 3838 1468 3842 1472
rect 3862 1468 3866 1472
rect 3886 1468 3890 1472
rect 3910 1468 3914 1472
rect 3966 1468 3970 1472
rect 4030 1468 4034 1472
rect 4142 1468 4146 1472
rect 4182 1468 4186 1472
rect 4214 1468 4218 1472
rect 4270 1468 4274 1472
rect 4342 1468 4346 1472
rect 4406 1468 4410 1472
rect 4574 1468 4578 1472
rect 4622 1468 4626 1472
rect 4734 1468 4738 1472
rect 4758 1468 4762 1472
rect 4774 1468 4778 1472
rect 4782 1468 4786 1472
rect 4814 1468 4818 1472
rect 4854 1468 4858 1472
rect 4878 1468 4882 1472
rect 4934 1468 4938 1472
rect 5014 1468 5018 1472
rect 5054 1468 5058 1472
rect 5126 1468 5130 1472
rect 5198 1468 5202 1472
rect 46 1458 50 1462
rect 110 1458 114 1462
rect 118 1458 122 1462
rect 150 1458 154 1462
rect 182 1458 186 1462
rect 198 1458 202 1462
rect 238 1458 242 1462
rect 262 1458 266 1462
rect 310 1458 314 1462
rect 342 1458 346 1462
rect 366 1458 370 1462
rect 390 1458 394 1462
rect 430 1458 434 1462
rect 454 1458 458 1462
rect 494 1458 498 1462
rect 590 1458 594 1462
rect 622 1458 626 1462
rect 678 1458 682 1462
rect 750 1458 754 1462
rect 774 1458 778 1462
rect 782 1458 786 1462
rect 838 1458 842 1462
rect 846 1458 850 1462
rect 870 1458 874 1462
rect 902 1458 906 1462
rect 974 1458 978 1462
rect 1046 1458 1050 1462
rect 1054 1458 1058 1462
rect 1062 1458 1066 1462
rect 1110 1458 1114 1462
rect 1166 1458 1170 1462
rect 1246 1458 1250 1462
rect 1254 1458 1258 1462
rect 1270 1458 1274 1462
rect 1286 1458 1290 1462
rect 1318 1458 1322 1462
rect 1326 1458 1330 1462
rect 1374 1458 1378 1462
rect 1406 1458 1410 1462
rect 1438 1458 1442 1462
rect 1446 1458 1450 1462
rect 1454 1458 1458 1462
rect 1502 1458 1506 1462
rect 1526 1458 1530 1462
rect 1550 1458 1554 1462
rect 1558 1458 1562 1462
rect 1574 1458 1578 1462
rect 1630 1458 1634 1462
rect 1702 1458 1706 1462
rect 1726 1458 1730 1462
rect 1734 1458 1738 1462
rect 1774 1458 1778 1462
rect 1782 1458 1786 1462
rect 1854 1458 1858 1462
rect 1886 1458 1890 1462
rect 1910 1458 1914 1462
rect 1934 1458 1938 1462
rect 1966 1458 1970 1462
rect 1974 1458 1978 1462
rect 2006 1458 2010 1462
rect 2014 1458 2018 1462
rect 2022 1458 2026 1462
rect 2062 1458 2066 1462
rect 2110 1458 2114 1462
rect 2174 1458 2178 1462
rect 2230 1458 2234 1462
rect 2238 1458 2242 1462
rect 2262 1458 2266 1462
rect 2286 1458 2290 1462
rect 2318 1458 2322 1462
rect 2382 1459 2386 1463
rect 2470 1458 2474 1462
rect 2502 1458 2506 1462
rect 2510 1458 2514 1462
rect 2542 1458 2546 1462
rect 2590 1459 2594 1463
rect 2614 1458 2618 1462
rect 2686 1458 2690 1462
rect 2694 1458 2698 1462
rect 2726 1458 2730 1462
rect 2758 1458 2762 1462
rect 2766 1458 2770 1462
rect 2806 1459 2810 1463
rect 2830 1458 2834 1462
rect 2878 1458 2882 1462
rect 2894 1458 2898 1462
rect 2926 1458 2930 1462
rect 2950 1458 2954 1462
rect 2958 1458 2962 1462
rect 2982 1458 2986 1462
rect 2998 1458 3002 1462
rect 3062 1458 3066 1462
rect 3078 1458 3082 1462
rect 3126 1458 3130 1462
rect 3134 1458 3138 1462
rect 3166 1458 3170 1462
rect 3230 1458 3234 1462
rect 3238 1458 3242 1462
rect 3278 1458 3282 1462
rect 3310 1458 3314 1462
rect 3358 1458 3362 1462
rect 3430 1458 3434 1462
rect 3438 1458 3442 1462
rect 3478 1458 3482 1462
rect 3510 1458 3514 1462
rect 3582 1458 3586 1462
rect 3638 1458 3642 1462
rect 3726 1458 3730 1462
rect 3790 1458 3794 1462
rect 3854 1458 3858 1462
rect 3862 1458 3866 1462
rect 3958 1459 3962 1463
rect 4038 1458 4042 1462
rect 4126 1459 4130 1463
rect 4166 1458 4170 1462
rect 4174 1458 4178 1462
rect 4182 1458 4186 1462
rect 4206 1458 4210 1462
rect 4286 1459 4290 1463
rect 4366 1458 4370 1462
rect 4374 1458 4378 1462
rect 4398 1458 4402 1462
rect 4430 1458 4434 1462
rect 4438 1458 4442 1462
rect 4550 1458 4554 1462
rect 4590 1458 4594 1462
rect 4598 1458 4602 1462
rect 4702 1458 4706 1462
rect 4766 1458 4770 1462
rect 4790 1458 4794 1462
rect 4806 1458 4810 1462
rect 4822 1458 4826 1462
rect 4846 1458 4850 1462
rect 4886 1458 4890 1462
rect 4926 1458 4930 1462
rect 4942 1458 4946 1462
rect 5014 1458 5018 1462
rect 5062 1458 5066 1462
rect 5102 1458 5106 1462
rect 5134 1458 5138 1462
rect 5142 1458 5146 1462
rect 5158 1458 5162 1462
rect 5166 1458 5170 1462
rect 5190 1458 5194 1462
rect 5246 1458 5250 1462
rect 102 1448 106 1452
rect 134 1448 138 1452
rect 166 1448 170 1452
rect 350 1448 354 1452
rect 406 1448 410 1452
rect 470 1448 474 1452
rect 478 1448 482 1452
rect 638 1448 642 1452
rect 1078 1448 1082 1452
rect 1126 1448 1130 1452
rect 1230 1448 1234 1452
rect 1350 1448 1354 1452
rect 1590 1448 1594 1452
rect 1758 1448 1762 1452
rect 2046 1448 2050 1452
rect 2078 1448 2082 1452
rect 2086 1448 2090 1452
rect 2102 1448 2106 1452
rect 2214 1448 2218 1452
rect 2246 1448 2250 1452
rect 2302 1448 2306 1452
rect 2318 1448 2322 1452
rect 2334 1448 2338 1452
rect 2430 1448 2434 1452
rect 2534 1448 2538 1452
rect 2774 1448 2778 1452
rect 3150 1448 3154 1452
rect 3622 1448 3626 1452
rect 3662 1448 3666 1452
rect 3814 1448 3818 1452
rect 3854 1448 3858 1452
rect 3894 1448 3898 1452
rect 4054 1448 4058 1452
rect 4158 1448 4162 1452
rect 4190 1448 4194 1452
rect 4382 1448 4386 1452
rect 4454 1448 4458 1452
rect 4750 1448 4754 1452
rect 4902 1448 4906 1452
rect 4926 1448 4930 1452
rect 5078 1448 5082 1452
rect 5150 1448 5154 1452
rect 1006 1438 1010 1442
rect 4006 1438 4010 1442
rect 4670 1438 4674 1442
rect 886 1428 890 1432
rect 1294 1428 1298 1432
rect 1334 1428 1338 1432
rect 4790 1428 4794 1432
rect 430 1418 434 1422
rect 454 1418 458 1422
rect 1430 1418 1434 1422
rect 1534 1418 1538 1422
rect 2670 1418 2674 1422
rect 5086 1418 5090 1422
rect 5102 1418 5106 1422
rect 330 1403 334 1407
rect 337 1403 341 1407
rect 1354 1403 1358 1407
rect 1361 1403 1365 1407
rect 2386 1403 2390 1407
rect 2393 1403 2397 1407
rect 3402 1403 3406 1407
rect 3409 1403 3413 1407
rect 4426 1403 4430 1407
rect 4433 1403 4437 1407
rect 14 1388 18 1392
rect 246 1388 250 1392
rect 310 1388 314 1392
rect 494 1388 498 1392
rect 654 1388 658 1392
rect 1078 1388 1082 1392
rect 1110 1388 1114 1392
rect 1230 1388 1234 1392
rect 1350 1388 1354 1392
rect 1566 1388 1570 1392
rect 1638 1388 1642 1392
rect 1782 1388 1786 1392
rect 1814 1388 1818 1392
rect 1838 1388 1842 1392
rect 1974 1388 1978 1392
rect 2030 1388 2034 1392
rect 2302 1388 2306 1392
rect 2350 1388 2354 1392
rect 2446 1388 2450 1392
rect 2750 1388 2754 1392
rect 2982 1388 2986 1392
rect 3030 1388 3034 1392
rect 3102 1388 3106 1392
rect 3686 1388 3690 1392
rect 3958 1388 3962 1392
rect 4326 1388 4330 1392
rect 4486 1388 4490 1392
rect 4638 1388 4642 1392
rect 4702 1388 4706 1392
rect 4790 1388 4794 1392
rect 5134 1388 5138 1392
rect 750 1378 754 1382
rect 4446 1378 4450 1382
rect 4518 1378 4522 1382
rect 4822 1378 4826 1382
rect 5062 1378 5066 1382
rect 166 1368 170 1372
rect 206 1368 210 1372
rect 766 1368 770 1372
rect 790 1368 794 1372
rect 1038 1368 1042 1372
rect 1102 1368 1106 1372
rect 1318 1368 1322 1372
rect 1630 1368 1634 1372
rect 1958 1368 1962 1372
rect 2142 1368 2146 1372
rect 2158 1368 2162 1372
rect 2190 1368 2194 1372
rect 2566 1368 2570 1372
rect 3270 1368 3274 1372
rect 3454 1368 3458 1372
rect 4246 1368 4250 1372
rect 4838 1368 4842 1372
rect 4926 1368 4930 1372
rect 4950 1368 4954 1372
rect 110 1348 114 1352
rect 182 1348 186 1352
rect 190 1348 194 1352
rect 502 1358 506 1362
rect 534 1358 538 1362
rect 222 1348 226 1352
rect 262 1348 266 1352
rect 278 1348 282 1352
rect 310 1348 314 1352
rect 382 1347 386 1351
rect 518 1348 522 1352
rect 534 1348 538 1352
rect 558 1348 562 1352
rect 70 1338 74 1342
rect 86 1338 90 1342
rect 174 1338 178 1342
rect 230 1338 234 1342
rect 270 1338 274 1342
rect 398 1338 402 1342
rect 414 1338 418 1342
rect 478 1338 482 1342
rect 526 1338 530 1342
rect 590 1347 594 1351
rect 622 1348 626 1352
rect 694 1348 698 1352
rect 718 1348 722 1352
rect 766 1348 770 1352
rect 910 1358 914 1362
rect 1022 1358 1026 1362
rect 1150 1358 1154 1362
rect 1158 1358 1162 1362
rect 806 1348 810 1352
rect 870 1348 874 1352
rect 950 1348 954 1352
rect 982 1348 986 1352
rect 1046 1348 1050 1352
rect 1054 1348 1058 1352
rect 1062 1348 1066 1352
rect 1086 1348 1090 1352
rect 1134 1348 1138 1352
rect 1142 1348 1146 1352
rect 1158 1348 1162 1352
rect 1174 1348 1178 1352
rect 1198 1348 1202 1352
rect 1238 1348 1242 1352
rect 1246 1348 1250 1352
rect 1254 1348 1258 1352
rect 1598 1358 1602 1362
rect 1614 1358 1618 1362
rect 2014 1358 2018 1362
rect 2046 1358 2050 1362
rect 2174 1358 2178 1362
rect 2206 1358 2210 1362
rect 2214 1358 2218 1362
rect 2254 1358 2258 1362
rect 2406 1358 2410 1362
rect 2422 1358 2426 1362
rect 2486 1358 2490 1362
rect 2502 1358 2506 1362
rect 2518 1358 2522 1362
rect 2526 1358 2530 1362
rect 2582 1358 2586 1362
rect 2614 1358 2618 1362
rect 3054 1358 3058 1362
rect 3142 1358 3146 1362
rect 3158 1358 3162 1362
rect 3174 1358 3178 1362
rect 3302 1358 3306 1362
rect 3318 1358 3322 1362
rect 3350 1358 3354 1362
rect 3382 1358 3386 1362
rect 3414 1358 3418 1362
rect 3438 1358 3442 1362
rect 3590 1358 3594 1362
rect 3750 1358 3754 1362
rect 3782 1358 3786 1362
rect 4302 1358 4306 1362
rect 4478 1358 4482 1362
rect 4502 1358 4506 1362
rect 4590 1358 4594 1362
rect 4598 1358 4602 1362
rect 4622 1358 4626 1362
rect 4686 1358 4690 1362
rect 4742 1358 4746 1362
rect 1334 1348 1338 1352
rect 1422 1348 1426 1352
rect 558 1338 562 1342
rect 670 1338 674 1342
rect 758 1338 762 1342
rect 830 1338 834 1342
rect 846 1338 850 1342
rect 958 1338 962 1342
rect 974 1338 978 1342
rect 1006 1340 1010 1344
rect 1014 1338 1018 1342
rect 1046 1338 1050 1342
rect 1118 1338 1122 1342
rect 1126 1338 1130 1342
rect 1486 1347 1490 1351
rect 1582 1348 1586 1352
rect 1598 1348 1602 1352
rect 1614 1348 1618 1352
rect 1638 1348 1642 1352
rect 1686 1348 1690 1352
rect 1286 1338 1290 1342
rect 1310 1338 1314 1342
rect 1358 1338 1362 1342
rect 1470 1338 1474 1342
rect 1574 1338 1578 1342
rect 1718 1347 1722 1351
rect 1790 1348 1794 1352
rect 1798 1348 1802 1352
rect 1822 1348 1826 1352
rect 1894 1347 1898 1351
rect 1974 1348 1978 1352
rect 2030 1348 2034 1352
rect 2094 1348 2098 1352
rect 2150 1348 2154 1352
rect 2190 1348 2194 1352
rect 2230 1348 2234 1352
rect 2238 1348 2242 1352
rect 2286 1348 2290 1352
rect 2302 1348 2306 1352
rect 2318 1348 2322 1352
rect 2334 1348 2338 1352
rect 2342 1348 2346 1352
rect 2398 1348 2402 1352
rect 2406 1348 2410 1352
rect 2430 1348 2434 1352
rect 2462 1348 2466 1352
rect 2478 1348 2482 1352
rect 2486 1348 2490 1352
rect 2518 1348 2522 1352
rect 2542 1348 2546 1352
rect 2566 1348 2570 1352
rect 2598 1348 2602 1352
rect 2662 1348 2666 1352
rect 2670 1348 2674 1352
rect 2742 1348 2746 1352
rect 2806 1348 2810 1352
rect 2870 1347 2874 1351
rect 2958 1348 2962 1352
rect 2966 1348 2970 1352
rect 2990 1348 2994 1352
rect 3014 1348 3018 1352
rect 3038 1348 3042 1352
rect 3046 1348 3050 1352
rect 3070 1348 3074 1352
rect 3086 1348 3090 1352
rect 3126 1348 3130 1352
rect 3142 1348 3146 1352
rect 3158 1348 3162 1352
rect 1606 1338 1610 1342
rect 1662 1338 1666 1342
rect 1702 1338 1706 1342
rect 1878 1338 1882 1342
rect 1966 1338 1970 1342
rect 1998 1338 2002 1342
rect 2014 1338 2018 1342
rect 2150 1338 2154 1342
rect 2182 1338 2186 1342
rect 2238 1338 2242 1342
rect 2326 1338 2330 1342
rect 2398 1338 2402 1342
rect 2462 1338 2466 1342
rect 2494 1338 2498 1342
rect 2550 1338 2554 1342
rect 2558 1338 2562 1342
rect 2590 1338 2594 1342
rect 2614 1338 2618 1342
rect 2798 1338 2802 1342
rect 3054 1338 3058 1342
rect 3078 1338 3082 1342
rect 3118 1338 3122 1342
rect 3206 1347 3210 1351
rect 3294 1348 3298 1352
rect 3334 1348 3338 1352
rect 3366 1348 3370 1352
rect 3398 1348 3402 1352
rect 3406 1348 3410 1352
rect 3502 1348 3506 1352
rect 3582 1348 3586 1352
rect 3614 1348 3618 1352
rect 3638 1348 3642 1352
rect 3646 1348 3650 1352
rect 3654 1348 3658 1352
rect 3686 1348 3690 1352
rect 3734 1348 3738 1352
rect 3766 1348 3770 1352
rect 3790 1348 3794 1352
rect 3822 1348 3826 1352
rect 3910 1348 3914 1352
rect 4006 1348 4010 1352
rect 4014 1348 4018 1352
rect 4062 1348 4066 1352
rect 4070 1348 4074 1352
rect 4094 1348 4098 1352
rect 4134 1347 4138 1351
rect 4214 1348 4218 1352
rect 4222 1348 4226 1352
rect 4254 1348 4258 1352
rect 4278 1348 4282 1352
rect 4286 1348 4290 1352
rect 4382 1348 4386 1352
rect 4390 1348 4394 1352
rect 4454 1348 4458 1352
rect 4518 1348 4522 1352
rect 4598 1348 4602 1352
rect 4638 1348 4642 1352
rect 4654 1348 4658 1352
rect 4702 1348 4706 1352
rect 4718 1348 4722 1352
rect 4734 1348 4738 1352
rect 4758 1348 4762 1352
rect 4774 1348 4778 1352
rect 4782 1348 4786 1352
rect 4806 1348 4810 1352
rect 3150 1338 3154 1342
rect 3190 1338 3194 1342
rect 3214 1338 3218 1342
rect 3326 1338 3330 1342
rect 3358 1338 3362 1342
rect 3382 1338 3386 1342
rect 3390 1338 3394 1342
rect 3542 1338 3546 1342
rect 3606 1338 3610 1342
rect 3662 1338 3666 1342
rect 3734 1338 3738 1342
rect 3758 1338 3762 1342
rect 3790 1338 3794 1342
rect 3798 1338 3802 1342
rect 3958 1338 3962 1342
rect 4102 1338 4106 1342
rect 4118 1338 4122 1342
rect 4494 1338 4498 1342
rect 4526 1338 4530 1342
rect 4534 1338 4538 1342
rect 4574 1338 4578 1342
rect 4614 1338 4618 1342
rect 4646 1338 4650 1342
rect 4886 1347 4890 1351
rect 4926 1348 4930 1352
rect 5022 1358 5026 1362
rect 5078 1358 5082 1362
rect 5174 1358 5178 1362
rect 4990 1348 4994 1352
rect 5006 1348 5010 1352
rect 5030 1348 5034 1352
rect 5046 1348 5050 1352
rect 5062 1348 5066 1352
rect 5110 1348 5114 1352
rect 5118 1348 5122 1352
rect 5302 1358 5306 1362
rect 5190 1348 5194 1352
rect 5198 1348 5202 1352
rect 4766 1338 4770 1342
rect 4902 1338 4906 1342
rect 4918 1338 4922 1342
rect 4990 1338 4994 1342
rect 4998 1338 5002 1342
rect 5054 1338 5058 1342
rect 5102 1338 5106 1342
rect 5238 1347 5242 1351
rect 5150 1338 5154 1342
rect 5206 1338 5210 1342
rect 5222 1338 5226 1342
rect 486 1328 490 1332
rect 1198 1328 1202 1332
rect 1430 1328 1434 1332
rect 1654 1328 1658 1332
rect 1862 1328 1866 1332
rect 2078 1328 2082 1332
rect 2262 1328 2266 1332
rect 2270 1328 2274 1332
rect 2726 1328 2730 1332
rect 2902 1328 2906 1332
rect 3278 1328 3282 1332
rect 3430 1328 3434 1332
rect 3558 1328 3562 1332
rect 3590 1328 3594 1332
rect 3678 1328 3682 1332
rect 3702 1328 3706 1332
rect 3726 1328 3730 1332
rect 3814 1328 3818 1332
rect 4246 1328 4250 1332
rect 4270 1328 4274 1332
rect 4406 1328 4410 1332
rect 4470 1328 4474 1332
rect 4670 1328 4674 1332
rect 4734 1328 4738 1332
rect 5030 1328 5034 1332
rect 5086 1328 5090 1332
rect 14 1318 18 1322
rect 502 1318 506 1322
rect 990 1318 994 1322
rect 1270 1318 1274 1322
rect 2214 1318 2218 1322
rect 2622 1318 2626 1322
rect 3350 1318 3354 1322
rect 3566 1318 3570 1322
rect 3670 1318 3674 1322
rect 3750 1318 3754 1322
rect 3806 1318 3810 1322
rect 3838 1318 3842 1322
rect 3854 1318 3858 1322
rect 4262 1318 4266 1322
rect 4542 1318 4546 1322
rect 4590 1318 4594 1322
rect 5038 1318 5042 1322
rect 5094 1318 5098 1322
rect 850 1303 854 1307
rect 857 1303 861 1307
rect 1874 1303 1878 1307
rect 1881 1303 1885 1307
rect 2890 1303 2894 1307
rect 2897 1303 2901 1307
rect 3922 1303 3926 1307
rect 3929 1303 3933 1307
rect 4938 1303 4942 1307
rect 4945 1303 4949 1307
rect 430 1288 434 1292
rect 446 1288 450 1292
rect 742 1288 746 1292
rect 886 1288 890 1292
rect 926 1288 930 1292
rect 982 1288 986 1292
rect 1022 1288 1026 1292
rect 1198 1288 1202 1292
rect 1414 1288 1418 1292
rect 1526 1288 1530 1292
rect 1582 1288 1586 1292
rect 1718 1288 1722 1292
rect 1830 1288 1834 1292
rect 1966 1288 1970 1292
rect 2134 1288 2138 1292
rect 2310 1288 2314 1292
rect 2438 1288 2442 1292
rect 2534 1288 2538 1292
rect 2766 1288 2770 1292
rect 3102 1288 3106 1292
rect 3230 1288 3234 1292
rect 3302 1288 3306 1292
rect 3462 1288 3466 1292
rect 3606 1288 3610 1292
rect 3702 1288 3706 1292
rect 4062 1288 4066 1292
rect 4094 1288 4098 1292
rect 4422 1288 4426 1292
rect 4462 1288 4466 1292
rect 4478 1288 4482 1292
rect 4606 1288 4610 1292
rect 4758 1288 4762 1292
rect 4926 1288 4930 1292
rect 4950 1288 4954 1292
rect 5078 1288 5082 1292
rect 5110 1288 5114 1292
rect 5206 1288 5210 1292
rect 182 1278 186 1282
rect 190 1278 194 1282
rect 438 1278 442 1282
rect 598 1278 602 1282
rect 766 1278 770 1282
rect 798 1278 802 1282
rect 806 1278 810 1282
rect 1398 1278 1402 1282
rect 1446 1278 1450 1282
rect 1534 1278 1538 1282
rect 1838 1278 1842 1282
rect 1846 1278 1850 1282
rect 1862 1278 1866 1282
rect 2302 1278 2306 1282
rect 2406 1278 2410 1282
rect 2494 1278 2498 1282
rect 3262 1278 3266 1282
rect 14 1268 18 1272
rect 102 1268 106 1272
rect 126 1268 130 1272
rect 158 1268 162 1272
rect 206 1268 210 1272
rect 398 1268 402 1272
rect 414 1268 418 1272
rect 494 1268 498 1272
rect 662 1268 666 1272
rect 758 1268 762 1272
rect 870 1268 874 1272
rect 894 1268 898 1272
rect 910 1268 914 1272
rect 38 1258 42 1262
rect 118 1258 122 1262
rect 134 1258 138 1262
rect 150 1258 154 1262
rect 158 1258 162 1262
rect 958 1268 962 1272
rect 1038 1268 1042 1272
rect 1046 1268 1050 1272
rect 1102 1268 1106 1272
rect 1214 1268 1218 1272
rect 1302 1268 1306 1272
rect 1358 1268 1362 1272
rect 1398 1268 1402 1272
rect 1406 1268 1410 1272
rect 1558 1268 1562 1272
rect 1654 1268 1658 1272
rect 1710 1268 1714 1272
rect 1782 1268 1786 1272
rect 1822 1268 1826 1272
rect 1926 1268 1930 1272
rect 1942 1268 1946 1272
rect 1982 1268 1986 1272
rect 2014 1268 2018 1272
rect 2078 1268 2082 1272
rect 2150 1268 2154 1272
rect 2238 1268 2242 1272
rect 2294 1268 2298 1272
rect 2382 1268 2386 1272
rect 2446 1268 2450 1272
rect 2462 1268 2466 1272
rect 2542 1268 2546 1272
rect 2606 1268 2610 1272
rect 2646 1268 2650 1272
rect 2718 1268 2722 1272
rect 2734 1268 2738 1272
rect 2790 1268 2794 1272
rect 2862 1268 2866 1272
rect 2870 1268 2874 1272
rect 2910 1268 2914 1272
rect 2966 1268 2970 1272
rect 2982 1268 2986 1272
rect 3094 1268 3098 1272
rect 3254 1268 3258 1272
rect 3278 1268 3282 1272
rect 3318 1278 3322 1282
rect 3798 1278 3802 1282
rect 3806 1278 3810 1282
rect 4070 1278 4074 1282
rect 4854 1278 4858 1282
rect 5270 1278 5274 1282
rect 3374 1268 3378 1272
rect 3478 1268 3482 1272
rect 3542 1268 3546 1272
rect 3622 1268 3626 1272
rect 3710 1268 3714 1272
rect 3742 1268 3746 1272
rect 238 1258 242 1262
rect 246 1258 250 1262
rect 270 1258 274 1262
rect 278 1258 282 1262
rect 294 1258 298 1262
rect 350 1258 354 1262
rect 374 1258 378 1262
rect 414 1258 418 1262
rect 486 1258 490 1262
rect 502 1258 506 1262
rect 574 1258 578 1262
rect 702 1258 706 1262
rect 750 1258 754 1262
rect 782 1258 786 1262
rect 822 1258 826 1262
rect 846 1258 850 1262
rect 902 1258 906 1262
rect 942 1258 946 1262
rect 950 1258 954 1262
rect 966 1258 970 1262
rect 1014 1258 1018 1262
rect 1054 1258 1058 1262
rect 1086 1258 1090 1262
rect 1094 1258 1098 1262
rect 1134 1259 1138 1263
rect 1166 1258 1170 1262
rect 1238 1258 1242 1262
rect 1310 1258 1314 1262
rect 1318 1258 1322 1262
rect 1350 1258 1354 1262
rect 1358 1258 1362 1262
rect 1414 1258 1418 1262
rect 1430 1258 1434 1262
rect 1462 1258 1466 1262
rect 1470 1258 1474 1262
rect 1478 1258 1482 1262
rect 1502 1258 1506 1262
rect 1518 1258 1522 1262
rect 1542 1258 1546 1262
rect 1598 1258 1602 1262
rect 1606 1258 1610 1262
rect 1614 1258 1618 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 1694 1258 1698 1262
rect 1702 1258 1706 1262
rect 1774 1258 1778 1262
rect 1814 1258 1818 1262
rect 1846 1258 1850 1262
rect 1950 1258 1954 1262
rect 1990 1258 1994 1262
rect 2006 1258 2010 1262
rect 2022 1258 2026 1262
rect 2070 1259 2074 1263
rect 2102 1258 2106 1262
rect 2174 1258 2178 1262
rect 2198 1258 2202 1262
rect 2246 1258 2250 1262
rect 2286 1258 2290 1262
rect 2422 1258 2426 1262
rect 2454 1258 2458 1262
rect 2478 1258 2482 1262
rect 2518 1258 2522 1262
rect 2542 1258 2546 1262
rect 2558 1258 2562 1262
rect 2598 1259 2602 1263
rect 2694 1258 2698 1262
rect 2742 1258 2746 1262
rect 2774 1258 2778 1262
rect 2782 1258 2786 1262
rect 2886 1258 2890 1262
rect 2918 1258 2922 1262
rect 2950 1258 2954 1262
rect 2958 1258 2962 1262
rect 2998 1259 3002 1263
rect 3070 1258 3074 1262
rect 3150 1258 3154 1262
rect 3182 1259 3186 1263
rect 3774 1268 3778 1272
rect 3790 1268 3794 1272
rect 3814 1268 3818 1272
rect 3830 1268 3834 1272
rect 3854 1268 3858 1272
rect 3878 1268 3882 1272
rect 3958 1268 3962 1272
rect 4054 1268 4058 1272
rect 4102 1268 4106 1272
rect 4166 1268 4170 1272
rect 4254 1268 4258 1272
rect 4302 1268 4306 1272
rect 4334 1268 4338 1272
rect 4350 1268 4354 1272
rect 4366 1268 4370 1272
rect 4382 1268 4386 1272
rect 4398 1268 4402 1272
rect 4574 1268 4578 1272
rect 4622 1268 4626 1272
rect 4838 1268 4842 1272
rect 4878 1268 4882 1272
rect 4894 1268 4898 1272
rect 4910 1268 4914 1272
rect 5046 1268 5050 1272
rect 5102 1268 5106 1272
rect 5190 1268 5194 1272
rect 3214 1258 3218 1262
rect 3222 1258 3226 1262
rect 3246 1258 3250 1262
rect 3286 1258 3290 1262
rect 3294 1258 3298 1262
rect 3334 1258 3338 1262
rect 3382 1258 3386 1262
rect 3502 1258 3506 1262
rect 3510 1258 3514 1262
rect 3550 1258 3554 1262
rect 3662 1258 3666 1262
rect 3718 1258 3722 1262
rect 3758 1258 3762 1262
rect 3782 1258 3786 1262
rect 3822 1258 3826 1262
rect 3838 1258 3842 1262
rect 3894 1258 3898 1262
rect 3918 1258 3922 1262
rect 3926 1258 3930 1262
rect 3974 1259 3978 1263
rect 4078 1258 4082 1262
rect 4134 1258 4138 1262
rect 4174 1258 4178 1262
rect 4262 1258 4266 1262
rect 4286 1258 4290 1262
rect 4294 1258 4298 1262
rect 4310 1258 4314 1262
rect 4326 1258 4330 1262
rect 4342 1258 4346 1262
rect 4374 1258 4378 1262
rect 4406 1258 4410 1262
rect 4446 1258 4450 1262
rect 4510 1258 4514 1262
rect 4542 1259 4546 1263
rect 4582 1258 4586 1262
rect 4590 1258 4594 1262
rect 4630 1258 4634 1262
rect 4694 1258 4698 1262
rect 4726 1259 4730 1263
rect 4822 1259 4826 1263
rect 4870 1258 4874 1262
rect 4902 1258 4906 1262
rect 4982 1258 4986 1262
rect 5014 1259 5018 1263
rect 5054 1258 5058 1262
rect 5094 1258 5098 1262
rect 5150 1258 5154 1262
rect 5246 1258 5250 1262
rect 5270 1259 5274 1263
rect 102 1248 106 1252
rect 134 1248 138 1252
rect 254 1248 258 1252
rect 886 1248 890 1252
rect 918 1248 922 1252
rect 926 1248 930 1252
rect 982 1248 986 1252
rect 1070 1248 1074 1252
rect 1334 1248 1338 1252
rect 1678 1248 1682 1252
rect 1942 1248 1946 1252
rect 2006 1248 2010 1252
rect 2038 1248 2042 1252
rect 2246 1248 2250 1252
rect 2486 1248 2490 1252
rect 2534 1248 2538 1252
rect 2566 1248 2570 1252
rect 2718 1248 2722 1252
rect 2934 1248 2938 1252
rect 3046 1248 3050 1252
rect 3742 1248 3746 1252
rect 3766 1248 3770 1252
rect 3862 1248 3866 1252
rect 4022 1248 4026 1252
rect 4326 1248 4330 1252
rect 4358 1248 4362 1252
rect 4390 1248 4394 1252
rect 4422 1248 4426 1252
rect 4598 1248 4602 1252
rect 4606 1248 4610 1252
rect 4926 1248 4930 1252
rect 5070 1248 5074 1252
rect 5222 1248 5226 1252
rect 94 1238 98 1242
rect 174 1238 178 1242
rect 726 1238 730 1242
rect 1022 1238 1026 1242
rect 1294 1238 1298 1242
rect 2022 1238 2026 1242
rect 2230 1238 2234 1242
rect 2270 1238 2274 1242
rect 2326 1238 2330 1242
rect 4966 1238 4970 1242
rect 1494 1228 1498 1232
rect 214 1218 218 1222
rect 646 1218 650 1222
rect 814 1218 818 1222
rect 830 1218 834 1222
rect 998 1218 1002 1222
rect 1630 1218 1634 1222
rect 1894 1218 1898 1222
rect 3910 1218 3914 1222
rect 4462 1218 4466 1222
rect 4646 1218 4650 1222
rect 4662 1218 4666 1222
rect 330 1203 334 1207
rect 337 1203 341 1207
rect 1354 1203 1358 1207
rect 1361 1203 1365 1207
rect 2386 1203 2390 1207
rect 2393 1203 2397 1207
rect 3402 1203 3406 1207
rect 3409 1203 3413 1207
rect 4426 1203 4430 1207
rect 4433 1203 4437 1207
rect 638 1188 642 1192
rect 806 1188 810 1192
rect 838 1188 842 1192
rect 1014 1188 1018 1192
rect 1046 1188 1050 1192
rect 1334 1188 1338 1192
rect 1382 1188 1386 1192
rect 1502 1188 1506 1192
rect 1598 1188 1602 1192
rect 1726 1188 1730 1192
rect 1734 1188 1738 1192
rect 1758 1188 1762 1192
rect 1854 1188 1858 1192
rect 1982 1188 1986 1192
rect 2030 1188 2034 1192
rect 2126 1188 2130 1192
rect 2302 1188 2306 1192
rect 2422 1188 2426 1192
rect 2566 1188 2570 1192
rect 2950 1188 2954 1192
rect 3030 1188 3034 1192
rect 3230 1188 3234 1192
rect 3310 1188 3314 1192
rect 3550 1188 3554 1192
rect 3766 1188 3770 1192
rect 3846 1188 3850 1192
rect 4150 1188 4154 1192
rect 4334 1188 4338 1192
rect 4358 1188 4362 1192
rect 4654 1188 4658 1192
rect 4726 1188 4730 1192
rect 5214 1188 5218 1192
rect 2542 1178 2546 1182
rect 3126 1178 3130 1182
rect 4638 1178 4642 1182
rect 150 1168 154 1172
rect 230 1168 234 1172
rect 918 1168 922 1172
rect 1198 1168 1202 1172
rect 1214 1168 1218 1172
rect 1694 1168 1698 1172
rect 2094 1168 2098 1172
rect 2718 1168 2722 1172
rect 4366 1168 4370 1172
rect 4502 1168 4506 1172
rect 4526 1168 4530 1172
rect 4662 1168 4666 1172
rect 4774 1168 4778 1172
rect 4870 1168 4874 1172
rect 4886 1168 4890 1172
rect 94 1158 98 1162
rect 102 1158 106 1162
rect 134 1158 138 1162
rect 182 1158 186 1162
rect 190 1158 194 1162
rect 246 1158 250 1162
rect 422 1158 426 1162
rect 438 1158 442 1162
rect 454 1158 458 1162
rect 558 1158 562 1162
rect 718 1158 722 1162
rect 854 1158 858 1162
rect 902 1158 906 1162
rect 942 1158 946 1162
rect 982 1158 986 1162
rect 1094 1158 1098 1162
rect 1254 1158 1258 1162
rect 1294 1158 1298 1162
rect 1398 1158 1402 1162
rect 1430 1158 1434 1162
rect 1438 1158 1442 1162
rect 1454 1158 1458 1162
rect 1822 1158 1826 1162
rect 2174 1158 2178 1162
rect 2294 1158 2298 1162
rect 2454 1158 2458 1162
rect 46 1148 50 1152
rect 102 1148 106 1152
rect 118 1148 122 1152
rect 158 1148 162 1152
rect 206 1148 210 1152
rect 214 1148 218 1152
rect 246 1148 250 1152
rect 342 1148 346 1152
rect 390 1148 394 1152
rect 406 1148 410 1152
rect 422 1148 426 1152
rect 510 1148 514 1152
rect 582 1148 586 1152
rect 606 1148 610 1152
rect 614 1148 618 1152
rect 630 1148 634 1152
rect 654 1148 658 1152
rect 678 1148 682 1152
rect 718 1148 722 1152
rect 758 1148 762 1152
rect 782 1148 786 1152
rect 814 1148 818 1152
rect 822 1148 826 1152
rect 838 1148 842 1152
rect 886 1148 890 1152
rect 918 1148 922 1152
rect 966 1148 970 1152
rect 974 1148 978 1152
rect 998 1148 1002 1152
rect 1022 1148 1026 1152
rect 1030 1148 1034 1152
rect 1062 1148 1066 1152
rect 1070 1148 1074 1152
rect 1102 1148 1106 1152
rect 1150 1147 1154 1151
rect 1222 1148 1226 1152
rect 1294 1148 1298 1152
rect 1310 1148 1314 1152
rect 1318 1148 1322 1152
rect 1342 1148 1346 1152
rect 1350 1148 1354 1152
rect 1414 1148 1418 1152
rect 1454 1148 1458 1152
rect 1486 1148 1490 1152
rect 1494 1148 1498 1152
rect 1502 1148 1506 1152
rect 1526 1148 1530 1152
rect 1558 1148 1562 1152
rect 1582 1148 1586 1152
rect 1614 1148 1618 1152
rect 1654 1148 1658 1152
rect 1774 1148 1778 1152
rect 1838 1148 1842 1152
rect 1870 1148 1874 1152
rect 1918 1147 1922 1151
rect 2014 1148 2018 1152
rect 2046 1148 2050 1152
rect 2054 1148 2058 1152
rect 2070 1148 2074 1152
rect 2094 1148 2098 1152
rect 2110 1148 2114 1152
rect 2158 1148 2162 1152
rect 2174 1148 2178 1152
rect 2206 1148 2210 1152
rect 2230 1148 2234 1152
rect 2262 1148 2266 1152
rect 2278 1148 2282 1152
rect 2326 1148 2330 1152
rect 2366 1148 2370 1152
rect 2454 1148 2458 1152
rect 2478 1158 2482 1162
rect 2534 1158 2538 1162
rect 2582 1158 2586 1162
rect 2782 1158 2786 1162
rect 2846 1158 2850 1162
rect 2878 1158 2882 1162
rect 2982 1158 2986 1162
rect 3046 1158 3050 1162
rect 3070 1158 3074 1162
rect 3078 1158 3082 1162
rect 3110 1158 3114 1162
rect 3246 1158 3250 1162
rect 3302 1158 3306 1162
rect 3422 1158 3426 1162
rect 3470 1158 3474 1162
rect 3510 1158 3514 1162
rect 3526 1158 3530 1162
rect 3534 1158 3538 1162
rect 3630 1158 3634 1162
rect 3758 1158 3762 1162
rect 4030 1158 4034 1162
rect 4134 1158 4138 1162
rect 4350 1158 4354 1162
rect 4382 1158 4386 1162
rect 4542 1158 4546 1162
rect 4558 1158 4562 1162
rect 4622 1158 4626 1162
rect 4670 1158 4674 1162
rect 4678 1158 4682 1162
rect 4902 1158 4906 1162
rect 4974 1158 4978 1162
rect 5102 1158 5106 1162
rect 5118 1158 5122 1162
rect 5134 1158 5138 1162
rect 2494 1148 2498 1152
rect 2510 1148 2514 1152
rect 2566 1148 2570 1152
rect 2590 1148 2594 1152
rect 2654 1148 2658 1152
rect 2734 1148 2738 1152
rect 2766 1148 2770 1152
rect 2774 1148 2778 1152
rect 2798 1148 2802 1152
rect 2838 1148 2842 1152
rect 2854 1148 2858 1152
rect 2862 1148 2866 1152
rect 2894 1148 2898 1152
rect 2918 1148 2922 1152
rect 2966 1148 2970 1152
rect 2998 1148 3002 1152
rect 3014 1148 3018 1152
rect 3030 1148 3034 1152
rect 3094 1148 3098 1152
rect 3126 1148 3130 1152
rect 3142 1148 3146 1152
rect 3246 1148 3250 1152
rect 3262 1148 3266 1152
rect 3278 1148 3282 1152
rect 3310 1148 3314 1152
rect 3358 1148 3362 1152
rect 3366 1148 3370 1152
rect 3374 1148 3378 1152
rect 3398 1148 3402 1152
rect 3454 1148 3458 1152
rect 3510 1148 3514 1152
rect 3550 1148 3554 1152
rect 3566 1148 3570 1152
rect 3574 1148 3578 1152
rect 3718 1148 3722 1152
rect 3774 1148 3778 1152
rect 3838 1148 3842 1152
rect 3894 1148 3898 1152
rect 3910 1148 3914 1152
rect 3974 1148 3978 1152
rect 4014 1148 4018 1152
rect 4030 1148 4034 1152
rect 4070 1148 4074 1152
rect 4078 1148 4082 1152
rect 4150 1148 4154 1152
rect 4166 1148 4170 1152
rect 4182 1148 4186 1152
rect 4254 1148 4258 1152
rect 4294 1148 4298 1152
rect 14 1138 18 1142
rect 126 1138 130 1142
rect 158 1138 162 1142
rect 166 1138 170 1142
rect 214 1138 218 1142
rect 222 1138 226 1142
rect 350 1138 354 1142
rect 398 1138 402 1142
rect 414 1138 418 1142
rect 430 1138 434 1142
rect 486 1138 490 1142
rect 582 1138 586 1142
rect 670 1138 674 1142
rect 702 1138 706 1142
rect 718 1138 722 1142
rect 830 1138 834 1142
rect 878 1138 882 1142
rect 910 1138 914 1142
rect 1078 1138 1082 1142
rect 1166 1138 1170 1142
rect 1270 1138 1274 1142
rect 1302 1138 1306 1142
rect 1374 1138 1378 1142
rect 1406 1138 1410 1142
rect 1462 1138 1466 1142
rect 1486 1138 1490 1142
rect 1550 1138 1554 1142
rect 1630 1138 1634 1142
rect 1934 1138 1938 1142
rect 2102 1138 2106 1142
rect 2134 1138 2138 1142
rect 2166 1138 2170 1142
rect 2198 1138 2202 1142
rect 2270 1138 2274 1142
rect 2318 1138 2322 1142
rect 2342 1138 2346 1142
rect 2446 1138 2450 1142
rect 2502 1138 2506 1142
rect 2534 1138 2538 1142
rect 2550 1138 2554 1142
rect 2558 1138 2562 1142
rect 2614 1138 2618 1142
rect 2734 1138 2738 1142
rect 2790 1138 2794 1142
rect 2806 1138 2810 1142
rect 2814 1138 2818 1142
rect 2830 1138 2834 1142
rect 2870 1138 2874 1142
rect 2886 1138 2890 1142
rect 2902 1138 2906 1142
rect 2958 1138 2962 1142
rect 3006 1138 3010 1142
rect 3022 1138 3026 1142
rect 3054 1138 3058 1142
rect 3102 1138 3106 1142
rect 3134 1138 3138 1142
rect 3150 1138 3154 1142
rect 3174 1138 3178 1142
rect 3270 1138 3274 1142
rect 3278 1138 3282 1142
rect 3350 1138 3354 1142
rect 3446 1138 3450 1142
rect 3502 1138 3506 1142
rect 3558 1138 3562 1142
rect 3598 1138 3602 1142
rect 3654 1138 3658 1142
rect 3742 1138 3746 1142
rect 3774 1138 3778 1142
rect 3958 1138 3962 1142
rect 4006 1138 4010 1142
rect 4158 1138 4162 1142
rect 4174 1138 4178 1142
rect 4278 1138 4282 1142
rect 4358 1148 4362 1152
rect 4382 1148 4386 1152
rect 4398 1148 4402 1152
rect 4470 1148 4474 1152
rect 4542 1148 4546 1152
rect 4558 1148 4562 1152
rect 4574 1148 4578 1152
rect 4598 1148 4602 1152
rect 4614 1148 4618 1152
rect 4638 1148 4642 1152
rect 4670 1148 4674 1152
rect 4734 1148 4738 1152
rect 4742 1148 4746 1152
rect 4750 1148 4754 1152
rect 4830 1148 4834 1152
rect 4886 1148 4890 1152
rect 4894 1148 4898 1152
rect 4918 1148 4922 1152
rect 4934 1148 4938 1152
rect 4998 1148 5002 1152
rect 5038 1148 5042 1152
rect 5046 1148 5050 1152
rect 5118 1148 5122 1152
rect 5150 1148 5154 1152
rect 5166 1148 5170 1152
rect 5174 1148 5178 1152
rect 5198 1148 5202 1152
rect 5246 1148 5250 1152
rect 5254 1148 5258 1152
rect 4406 1138 4410 1142
rect 4462 1138 4466 1142
rect 4550 1138 4554 1142
rect 4590 1138 4594 1142
rect 4606 1138 4610 1142
rect 4646 1138 4650 1142
rect 4814 1138 4818 1142
rect 4838 1138 4842 1142
rect 4894 1138 4898 1142
rect 4926 1138 4930 1142
rect 4990 1138 4994 1142
rect 5126 1138 5130 1142
rect 5158 1138 5162 1142
rect 5198 1138 5202 1142
rect 5270 1138 5274 1142
rect 694 1128 698 1132
rect 774 1128 778 1132
rect 942 1128 946 1132
rect 1118 1128 1122 1132
rect 1150 1128 1154 1132
rect 1470 1128 1474 1132
rect 1534 1128 1538 1132
rect 1742 1128 1746 1132
rect 1950 1128 1954 1132
rect 2054 1128 2058 1132
rect 2070 1128 2074 1132
rect 2142 1128 2146 1132
rect 2526 1128 2530 1132
rect 2646 1128 2650 1132
rect 2814 1128 2818 1132
rect 2910 1128 2914 1132
rect 2950 1128 2954 1132
rect 3166 1128 3170 1132
rect 3326 1128 3330 1132
rect 3334 1128 3338 1132
rect 3438 1128 3442 1132
rect 3494 1128 3498 1132
rect 3622 1128 3626 1132
rect 4190 1128 4194 1132
rect 4326 1128 4330 1132
rect 4342 1128 4346 1132
rect 4590 1128 4594 1132
rect 4686 1128 4690 1132
rect 4950 1128 4954 1132
rect 5070 1128 5074 1132
rect 182 1118 186 1122
rect 190 1118 194 1122
rect 270 1118 274 1122
rect 286 1118 290 1122
rect 742 1118 746 1122
rect 902 1118 906 1122
rect 1238 1118 1242 1122
rect 1430 1118 1434 1122
rect 1734 1118 1738 1122
rect 1758 1118 1762 1122
rect 1798 1118 1802 1122
rect 1998 1118 2002 1122
rect 2214 1118 2218 1122
rect 2246 1118 2250 1122
rect 2518 1118 2522 1122
rect 3070 1118 3074 1122
rect 3078 1118 3082 1122
rect 3158 1118 3162 1122
rect 3230 1118 3234 1122
rect 3302 1118 3306 1122
rect 3318 1118 3322 1122
rect 3342 1118 3346 1122
rect 3390 1118 3394 1122
rect 3486 1118 3490 1122
rect 3630 1118 3634 1122
rect 3662 1118 3666 1122
rect 3798 1118 3802 1122
rect 3822 1118 3826 1122
rect 3990 1118 3994 1122
rect 4038 1118 4042 1122
rect 4198 1118 4202 1122
rect 4758 1118 4762 1122
rect 5006 1118 5010 1122
rect 5134 1118 5138 1122
rect 850 1103 854 1107
rect 857 1103 861 1107
rect 1874 1103 1878 1107
rect 1881 1103 1885 1107
rect 2890 1103 2894 1107
rect 2897 1103 2901 1107
rect 3922 1103 3926 1107
rect 3929 1103 3933 1107
rect 4938 1103 4942 1107
rect 4945 1103 4949 1107
rect 254 1088 258 1092
rect 366 1088 370 1092
rect 374 1088 378 1092
rect 494 1088 498 1092
rect 590 1088 594 1092
rect 670 1088 674 1092
rect 798 1088 802 1092
rect 814 1088 818 1092
rect 942 1088 946 1092
rect 958 1088 962 1092
rect 982 1088 986 1092
rect 1022 1088 1026 1092
rect 1182 1088 1186 1092
rect 1486 1088 1490 1092
rect 1654 1088 1658 1092
rect 1758 1088 1762 1092
rect 1894 1088 1898 1092
rect 1918 1088 1922 1092
rect 2102 1088 2106 1092
rect 2158 1088 2162 1092
rect 2526 1088 2530 1092
rect 2654 1088 2658 1092
rect 2878 1088 2882 1092
rect 3134 1088 3138 1092
rect 3142 1088 3146 1092
rect 3494 1088 3498 1092
rect 3574 1088 3578 1092
rect 3758 1088 3762 1092
rect 3806 1088 3810 1092
rect 3982 1088 3986 1092
rect 4038 1088 4042 1092
rect 4086 1088 4090 1092
rect 4134 1088 4138 1092
rect 4158 1088 4162 1092
rect 4246 1088 4250 1092
rect 4526 1088 4530 1092
rect 4582 1088 4586 1092
rect 4654 1088 4658 1092
rect 4750 1088 4754 1092
rect 4918 1088 4922 1092
rect 5014 1088 5018 1092
rect 5118 1088 5122 1092
rect 5150 1088 5154 1092
rect 62 1078 66 1082
rect 430 1078 434 1082
rect 526 1078 530 1082
rect 646 1078 650 1082
rect 678 1078 682 1082
rect 734 1078 738 1082
rect 1086 1078 1090 1082
rect 1318 1078 1322 1082
rect 1422 1078 1426 1082
rect 1454 1078 1458 1082
rect 1566 1078 1570 1082
rect 14 1068 18 1072
rect 118 1068 122 1072
rect 174 1068 178 1072
rect 262 1068 266 1072
rect 294 1068 298 1072
rect 326 1068 330 1072
rect 398 1068 402 1072
rect 606 1068 610 1072
rect 662 1068 666 1072
rect 702 1068 706 1072
rect 878 1068 882 1072
rect 966 1068 970 1072
rect 990 1068 994 1072
rect 998 1068 1002 1072
rect 1070 1068 1074 1072
rect 1102 1068 1106 1072
rect 1198 1068 1202 1072
rect 1366 1068 1370 1072
rect 1390 1068 1394 1072
rect 1406 1068 1410 1072
rect 1822 1078 1826 1082
rect 1950 1078 1954 1082
rect 2006 1078 2010 1082
rect 2038 1078 2042 1082
rect 2430 1078 2434 1082
rect 3038 1078 3042 1082
rect 3206 1078 3210 1082
rect 3334 1078 3338 1082
rect 3366 1078 3370 1082
rect 3430 1078 3434 1082
rect 3606 1078 3610 1082
rect 3622 1078 3626 1082
rect 3670 1078 3674 1082
rect 3718 1078 3722 1082
rect 3742 1078 3746 1082
rect 3750 1078 3754 1082
rect 4022 1078 4026 1082
rect 1502 1068 1506 1072
rect 1550 1068 1554 1072
rect 1614 1068 1618 1072
rect 1630 1068 1634 1072
rect 1750 1068 1754 1072
rect 1854 1068 1858 1072
rect 1910 1068 1914 1072
rect 1966 1068 1970 1072
rect 2134 1068 2138 1072
rect 2222 1068 2226 1072
rect 2270 1068 2274 1072
rect 2326 1068 2330 1072
rect 2382 1068 2386 1072
rect 2414 1068 2418 1072
rect 2534 1068 2538 1072
rect 2574 1068 2578 1072
rect 2662 1068 2666 1072
rect 2694 1068 2698 1072
rect 2718 1068 2722 1072
rect 2726 1068 2730 1072
rect 2766 1068 2770 1072
rect 2782 1068 2786 1072
rect 2910 1068 2914 1072
rect 3022 1068 3026 1072
rect 3070 1068 3074 1072
rect 3238 1068 3242 1072
rect 3294 1068 3298 1072
rect 3302 1068 3306 1072
rect 3502 1068 3506 1072
rect 3534 1068 3538 1072
rect 3654 1068 3658 1072
rect 3662 1068 3666 1072
rect 3694 1068 3698 1072
rect 3718 1068 3722 1072
rect 3854 1068 3858 1072
rect 3886 1068 3890 1072
rect 3902 1068 3906 1072
rect 3918 1068 3922 1072
rect 3974 1068 3978 1072
rect 4118 1078 4122 1082
rect 4150 1078 4154 1082
rect 4238 1078 4242 1082
rect 4302 1078 4306 1082
rect 4462 1078 4466 1082
rect 4550 1078 4554 1082
rect 4814 1078 4818 1082
rect 4846 1078 4850 1082
rect 5110 1078 5114 1082
rect 5270 1078 5274 1082
rect 4046 1068 4050 1072
rect 4126 1068 4130 1072
rect 4166 1068 4170 1072
rect 4182 1068 4186 1072
rect 4230 1068 4234 1072
rect 4254 1068 4258 1072
rect 4350 1068 4354 1072
rect 4366 1068 4370 1072
rect 4390 1068 4394 1072
rect 4414 1068 4418 1072
rect 4558 1068 4562 1072
rect 4606 1068 4610 1072
rect 4622 1068 4626 1072
rect 4638 1068 4642 1072
rect 4646 1068 4650 1072
rect 4678 1068 4682 1072
rect 4686 1068 4690 1072
rect 4742 1068 4746 1072
rect 4886 1068 4890 1072
rect 4966 1068 4970 1072
rect 5070 1068 5074 1072
rect 5126 1068 5130 1072
rect 5190 1068 5194 1072
rect 38 1058 42 1062
rect 118 1058 122 1062
rect 126 1058 130 1062
rect 150 1058 154 1062
rect 158 1058 162 1062
rect 190 1059 194 1063
rect 270 1058 274 1062
rect 294 1058 298 1062
rect 302 1058 306 1062
rect 334 1058 338 1062
rect 390 1058 394 1062
rect 430 1059 434 1063
rect 534 1058 538 1062
rect 598 1058 602 1062
rect 614 1058 618 1062
rect 630 1058 634 1062
rect 646 1058 650 1062
rect 742 1058 746 1062
rect 830 1058 834 1062
rect 902 1058 906 1062
rect 1006 1058 1010 1062
rect 1030 1058 1034 1062
rect 1038 1058 1042 1062
rect 1062 1058 1066 1062
rect 1118 1059 1122 1063
rect 1222 1058 1226 1062
rect 1302 1058 1306 1062
rect 1310 1058 1314 1062
rect 1334 1058 1338 1062
rect 1374 1058 1378 1062
rect 1422 1059 1426 1063
rect 1526 1058 1530 1062
rect 1606 1058 1610 1062
rect 1646 1058 1650 1062
rect 1678 1058 1682 1062
rect 1710 1058 1714 1062
rect 1718 1058 1722 1062
rect 1742 1058 1746 1062
rect 1814 1058 1818 1062
rect 1862 1058 1866 1062
rect 1902 1058 1906 1062
rect 1934 1058 1938 1062
rect 1958 1058 1962 1062
rect 1990 1058 1994 1062
rect 2038 1059 2042 1063
rect 2142 1058 2146 1062
rect 2166 1058 2170 1062
rect 2198 1058 2202 1062
rect 2262 1058 2266 1062
rect 2334 1058 2338 1062
rect 2342 1058 2346 1062
rect 2374 1058 2378 1062
rect 2406 1058 2410 1062
rect 2462 1059 2466 1063
rect 2494 1058 2498 1062
rect 2558 1058 2562 1062
rect 2598 1058 2602 1062
rect 2670 1058 2674 1062
rect 2710 1058 2714 1062
rect 2734 1058 2738 1062
rect 2774 1058 2778 1062
rect 2814 1059 2818 1063
rect 2838 1058 2842 1062
rect 2926 1058 2930 1062
rect 2942 1058 2946 1062
rect 2966 1058 2970 1062
rect 2974 1058 2978 1062
rect 2982 1058 2986 1062
rect 2990 1058 2994 1062
rect 3078 1058 3082 1062
rect 3206 1059 3210 1063
rect 3246 1058 3250 1062
rect 3254 1058 3258 1062
rect 3286 1058 3290 1062
rect 3302 1058 3306 1062
rect 3350 1058 3354 1062
rect 3382 1058 3386 1062
rect 3430 1059 3434 1063
rect 3526 1058 3530 1062
rect 3542 1058 3546 1062
rect 3574 1058 3578 1062
rect 3590 1058 3594 1062
rect 3622 1058 3626 1062
rect 3646 1058 3650 1062
rect 3670 1058 3674 1062
rect 3686 1058 3690 1062
rect 3702 1058 3706 1062
rect 3718 1058 3722 1062
rect 3726 1058 3730 1062
rect 3766 1058 3770 1062
rect 3798 1058 3802 1062
rect 3870 1059 3874 1063
rect 3958 1058 3962 1062
rect 3998 1058 4002 1062
rect 4006 1058 4010 1062
rect 4054 1058 4058 1062
rect 4094 1058 4098 1062
rect 4102 1058 4106 1062
rect 4118 1058 4122 1062
rect 4174 1058 4178 1062
rect 4206 1058 4210 1062
rect 4222 1058 4226 1062
rect 4334 1059 4338 1063
rect 4406 1058 4410 1062
rect 4486 1058 4490 1062
rect 4494 1058 4498 1062
rect 4534 1058 4538 1062
rect 4550 1058 4554 1062
rect 4566 1058 4570 1062
rect 4630 1058 4634 1062
rect 4654 1058 4658 1062
rect 4670 1058 4674 1062
rect 4694 1058 4698 1062
rect 4726 1058 4730 1062
rect 4734 1058 4738 1062
rect 4806 1058 4810 1062
rect 4862 1058 4866 1062
rect 4878 1058 4882 1062
rect 4894 1058 4898 1062
rect 4974 1058 4978 1062
rect 5078 1059 5082 1063
rect 5134 1058 5138 1062
rect 5158 1058 5162 1062
rect 5166 1058 5170 1062
rect 5190 1058 5194 1062
rect 5246 1058 5250 1062
rect 286 1048 290 1052
rect 318 1048 322 1052
rect 366 1048 370 1052
rect 374 1048 378 1052
rect 686 1048 690 1052
rect 966 1048 970 1052
rect 1022 1048 1026 1052
rect 1286 1048 1290 1052
rect 1390 1048 1394 1052
rect 1878 1048 1882 1052
rect 1982 1048 1986 1052
rect 2110 1048 2114 1052
rect 2126 1048 2130 1052
rect 2158 1048 2162 1052
rect 2358 1048 2362 1052
rect 2430 1048 2434 1052
rect 2686 1048 2690 1052
rect 2750 1048 2754 1052
rect 3270 1048 3274 1052
rect 3326 1048 3330 1052
rect 3558 1048 3562 1052
rect 3630 1048 3634 1052
rect 3918 1048 3922 1052
rect 4142 1048 4146 1052
rect 4198 1048 4202 1052
rect 4206 1048 4210 1052
rect 4382 1048 4386 1052
rect 4590 1048 4594 1052
rect 4614 1048 4618 1052
rect 4710 1048 4714 1052
rect 5150 1048 5154 1052
rect 702 1038 706 1042
rect 950 1038 954 1042
rect 1262 1038 1266 1042
rect 1566 1038 1570 1042
rect 2318 1038 2322 1042
rect 1054 1028 1058 1032
rect 254 1018 258 1022
rect 302 1018 306 1022
rect 1694 1018 1698 1022
rect 2182 1018 2186 1022
rect 2958 1018 2962 1022
rect 3782 1018 3786 1022
rect 3982 1018 3986 1022
rect 4190 1018 4194 1022
rect 5014 1018 5018 1022
rect 5206 1018 5210 1022
rect 330 1003 334 1007
rect 337 1003 341 1007
rect 1354 1003 1358 1007
rect 1361 1003 1365 1007
rect 2386 1003 2390 1007
rect 2393 1003 2397 1007
rect 3402 1003 3406 1007
rect 3409 1003 3413 1007
rect 4426 1003 4430 1007
rect 4433 1003 4437 1007
rect 222 988 226 992
rect 454 988 458 992
rect 798 988 802 992
rect 814 988 818 992
rect 998 988 1002 992
rect 1030 988 1034 992
rect 1190 988 1194 992
rect 1278 988 1282 992
rect 1614 988 1618 992
rect 1654 988 1658 992
rect 1686 988 1690 992
rect 2134 988 2138 992
rect 2310 988 2314 992
rect 2750 988 2754 992
rect 2806 988 2810 992
rect 3022 988 3026 992
rect 3134 988 3138 992
rect 3446 988 3450 992
rect 3830 988 3834 992
rect 4166 988 4170 992
rect 4214 988 4218 992
rect 4406 988 4410 992
rect 4838 988 4842 992
rect 4862 988 4866 992
rect 5150 988 5154 992
rect 5278 988 5282 992
rect 198 978 202 982
rect 566 978 570 982
rect 2110 978 2114 982
rect 4646 978 4650 982
rect 94 968 98 972
rect 134 968 138 972
rect 318 968 322 972
rect 686 968 690 972
rect 958 968 962 972
rect 1502 968 1506 972
rect 1958 968 1962 972
rect 2022 968 2026 972
rect 2038 968 2042 972
rect 2582 968 2586 972
rect 2718 968 2722 972
rect 2942 968 2946 972
rect 3174 968 3178 972
rect 3854 968 3858 972
rect 110 958 114 962
rect 38 948 42 952
rect 110 948 114 952
rect 182 958 186 962
rect 238 958 242 962
rect 302 958 306 962
rect 334 958 338 962
rect 398 958 402 962
rect 702 958 706 962
rect 150 948 154 952
rect 198 948 202 952
rect 222 948 226 952
rect 246 948 250 952
rect 262 948 266 952
rect 278 948 282 952
rect 350 948 354 952
rect 366 948 370 952
rect 398 948 402 952
rect 414 948 418 952
rect 438 948 442 952
rect 462 948 466 952
rect 470 948 474 952
rect 510 948 514 952
rect 574 948 578 952
rect 606 948 610 952
rect 654 948 658 952
rect 686 948 690 952
rect 734 947 738 951
rect 814 948 818 952
rect 838 958 842 962
rect 942 958 946 962
rect 1022 958 1026 962
rect 886 948 890 952
rect 910 948 914 952
rect 918 948 922 952
rect 958 948 962 952
rect 974 948 978 952
rect 982 948 986 952
rect 1006 948 1010 952
rect 1054 948 1058 952
rect 1078 958 1082 962
rect 1094 948 1098 952
rect 1118 948 1122 952
rect 1126 948 1130 952
rect 1142 958 1146 962
rect 1238 958 1242 962
rect 1166 948 1170 952
rect 1174 948 1178 952
rect 1198 948 1202 952
rect 1222 948 1226 952
rect 1446 958 1450 962
rect 1494 958 1498 962
rect 2054 958 2058 962
rect 2670 958 2674 962
rect 2734 958 2738 962
rect 2766 958 2770 962
rect 2790 958 2794 962
rect 1262 948 1266 952
rect 1318 948 1322 952
rect 1414 948 1418 952
rect 1422 948 1426 952
rect 1454 948 1458 952
rect 1478 948 1482 952
rect 1558 948 1562 952
rect 1598 948 1602 952
rect 1638 948 1642 952
rect 1662 948 1666 952
rect 1670 948 1674 952
rect 1678 948 1682 952
rect 1702 948 1706 952
rect 1750 948 1754 952
rect 1806 948 1810 952
rect 1910 948 1914 952
rect 1966 948 1970 952
rect 2014 948 2018 952
rect 2038 948 2042 952
rect 2070 948 2074 952
rect 2086 948 2090 952
rect 2094 948 2098 952
rect 2118 948 2122 952
rect 2198 948 2202 952
rect 2262 948 2266 952
rect 2286 948 2290 952
rect 2302 948 2306 952
rect 2326 948 2330 952
rect 2334 948 2338 952
rect 2430 948 2434 952
rect 2462 948 2466 952
rect 2518 948 2522 952
rect 2598 948 2602 952
rect 2606 948 2610 952
rect 2630 948 2634 952
rect 2638 948 2642 952
rect 2646 948 2650 952
rect 2686 948 2690 952
rect 2702 948 2706 952
rect 2718 948 2722 952
rect 2750 948 2754 952
rect 2806 948 2810 952
rect 2830 958 2834 962
rect 2918 958 2922 962
rect 2870 948 2874 952
rect 2910 948 2914 952
rect 2966 948 2970 952
rect 3070 948 3074 952
rect 3094 948 3098 952
rect 102 938 106 942
rect 158 938 162 942
rect 206 938 210 942
rect 214 938 218 942
rect 270 938 274 942
rect 278 938 282 942
rect 310 938 314 942
rect 358 938 362 942
rect 422 938 426 942
rect 486 938 490 942
rect 526 938 530 942
rect 582 938 586 942
rect 718 938 722 942
rect 806 938 810 942
rect 870 938 874 942
rect 926 938 930 942
rect 966 938 970 942
rect 1038 938 1042 942
rect 1046 938 1050 942
rect 1102 938 1106 942
rect 1110 938 1114 942
rect 1158 938 1162 942
rect 1214 938 1218 942
rect 1246 938 1250 942
rect 1270 938 1274 942
rect 1334 938 1338 942
rect 1374 938 1378 942
rect 1430 938 1434 942
rect 1566 938 1570 942
rect 1734 938 1738 942
rect 1742 938 1746 942
rect 1902 938 1906 942
rect 1974 938 1978 942
rect 1982 938 1986 942
rect 2046 938 2050 942
rect 2078 938 2082 942
rect 2230 938 2234 942
rect 2246 938 2250 942
rect 2270 938 2274 942
rect 2406 938 2410 942
rect 2438 938 2442 942
rect 2454 938 2458 942
rect 2494 938 2498 942
rect 3246 947 3250 951
rect 3286 948 3290 952
rect 3310 948 3314 952
rect 3318 948 3322 952
rect 3358 948 3362 952
rect 3454 948 3458 952
rect 3462 948 3466 952
rect 3494 948 3498 952
rect 3510 948 3514 952
rect 3542 948 3546 952
rect 3590 948 3594 952
rect 3622 948 3626 952
rect 3662 948 3666 952
rect 3734 948 3738 952
rect 3742 948 3746 952
rect 3758 958 3762 962
rect 3782 958 3786 962
rect 4198 958 4202 962
rect 4206 958 4210 962
rect 4222 958 4226 962
rect 4262 958 4266 962
rect 4390 958 4394 962
rect 4438 958 4442 962
rect 4638 958 4642 962
rect 4758 958 4762 962
rect 4806 958 4810 962
rect 4910 958 4914 962
rect 5270 958 5274 962
rect 3774 948 3778 952
rect 3798 948 3802 952
rect 3830 948 3834 952
rect 3886 948 3890 952
rect 3950 948 3954 952
rect 4014 948 4018 952
rect 4038 948 4042 952
rect 4078 948 4082 952
rect 4110 948 4114 952
rect 4134 948 4138 952
rect 4182 948 4186 952
rect 4198 948 4202 952
rect 4246 948 4250 952
rect 4262 948 4266 952
rect 4278 948 4282 952
rect 4334 948 4338 952
rect 4406 948 4410 952
rect 4454 948 4458 952
rect 4470 948 4474 952
rect 4510 948 4514 952
rect 2646 938 2650 942
rect 2694 938 2698 942
rect 2710 938 2714 942
rect 2742 938 2746 942
rect 2774 938 2778 942
rect 2790 938 2794 942
rect 2854 938 2858 942
rect 2894 938 2898 942
rect 3006 938 3010 942
rect 3150 938 3154 942
rect 3262 938 3266 942
rect 3278 938 3282 942
rect 3334 938 3338 942
rect 3438 938 3442 942
rect 3470 938 3474 942
rect 3486 938 3490 942
rect 3614 938 3618 942
rect 3638 938 3642 942
rect 3726 938 3730 942
rect 3774 938 3778 942
rect 3806 938 3810 942
rect 3918 938 3922 942
rect 3990 938 3994 942
rect 4086 938 4090 942
rect 4182 938 4186 942
rect 4222 938 4226 942
rect 4254 938 4258 942
rect 4286 938 4290 942
rect 4302 938 4306 942
rect 4374 938 4378 942
rect 4542 947 4546 951
rect 4574 948 4578 952
rect 4622 948 4626 952
rect 4630 948 4634 952
rect 4702 948 4706 952
rect 4782 948 4786 952
rect 4830 948 4834 952
rect 4838 948 4842 952
rect 4862 948 4866 952
rect 4886 948 4890 952
rect 4934 948 4938 952
rect 5006 948 5010 952
rect 5110 948 5114 952
rect 5198 948 5202 952
rect 5246 948 5250 952
rect 4462 938 4466 942
rect 4526 938 4530 942
rect 4614 938 4618 942
rect 4694 938 4698 942
rect 4766 938 4770 942
rect 4830 938 4834 942
rect 4926 938 4930 942
rect 5038 938 5042 942
rect 5134 938 5138 942
rect 5206 938 5210 942
rect 5286 938 5290 942
rect 30 928 34 932
rect 166 928 170 932
rect 374 928 378 932
rect 382 928 386 932
rect 590 928 594 932
rect 622 928 626 932
rect 662 928 666 932
rect 766 928 770 932
rect 902 928 906 932
rect 926 928 930 932
rect 1702 928 1706 932
rect 1718 928 1722 932
rect 1998 928 2002 932
rect 2246 928 2250 932
rect 2270 928 2274 932
rect 2478 928 2482 932
rect 2886 928 2890 932
rect 3134 928 3138 932
rect 3510 928 3514 932
rect 3534 928 3538 932
rect 3574 928 3578 932
rect 3814 928 3818 932
rect 4094 928 4098 932
rect 4134 928 4138 932
rect 4150 928 4154 932
rect 4486 928 4490 932
rect 4494 928 4498 932
rect 4510 928 4514 932
rect 4590 928 4594 932
rect 4654 928 4658 932
rect 4798 928 4802 932
rect 4854 928 4858 932
rect 4878 928 4882 932
rect 4902 928 4906 932
rect 4950 928 4954 932
rect 5262 928 5266 932
rect 174 918 178 922
rect 302 918 306 922
rect 398 918 402 922
rect 638 918 642 922
rect 1070 918 1074 922
rect 1494 918 1498 922
rect 1614 918 1618 922
rect 1758 918 1762 922
rect 2054 918 2058 922
rect 2350 918 2354 922
rect 2790 918 2794 922
rect 3526 918 3530 922
rect 3558 918 3562 922
rect 3606 918 3610 922
rect 3718 918 3722 922
rect 3838 918 3842 922
rect 3966 918 3970 922
rect 4070 918 4074 922
rect 4230 918 4234 922
rect 4478 918 4482 922
rect 4750 918 4754 922
rect 4806 918 4810 922
rect 5054 918 5058 922
rect 5254 918 5258 922
rect 850 903 854 907
rect 857 903 861 907
rect 1874 903 1878 907
rect 1881 903 1885 907
rect 2890 903 2894 907
rect 2897 903 2901 907
rect 3922 903 3926 907
rect 3929 903 3933 907
rect 4938 903 4942 907
rect 4945 903 4949 907
rect 94 888 98 892
rect 214 888 218 892
rect 222 888 226 892
rect 486 888 490 892
rect 558 888 562 892
rect 686 888 690 892
rect 814 888 818 892
rect 934 888 938 892
rect 1038 888 1042 892
rect 1198 888 1202 892
rect 1622 888 1626 892
rect 1726 888 1730 892
rect 1822 888 1826 892
rect 1990 888 1994 892
rect 2174 888 2178 892
rect 2374 888 2378 892
rect 2510 888 2514 892
rect 2526 888 2530 892
rect 2638 888 2642 892
rect 2766 888 2770 892
rect 2846 888 2850 892
rect 2982 888 2986 892
rect 3046 888 3050 892
rect 3086 888 3090 892
rect 3254 888 3258 892
rect 3374 888 3378 892
rect 3446 888 3450 892
rect 3550 888 3554 892
rect 3670 888 3674 892
rect 3718 888 3722 892
rect 3814 888 3818 892
rect 3886 888 3890 892
rect 3998 888 4002 892
rect 4238 888 4242 892
rect 4334 888 4338 892
rect 4374 888 4378 892
rect 4510 888 4514 892
rect 4582 888 4586 892
rect 4670 888 4674 892
rect 4702 888 4706 892
rect 4830 888 4834 892
rect 4838 888 4842 892
rect 5038 888 5042 892
rect 5062 888 5066 892
rect 30 878 34 882
rect 150 878 154 882
rect 382 878 386 882
rect 598 878 602 882
rect 718 878 722 882
rect 918 878 922 882
rect 1406 878 1410 882
rect 1646 878 1650 882
rect 110 868 114 872
rect 158 868 162 872
rect 190 868 194 872
rect 246 868 250 872
rect 262 868 266 872
rect 446 868 450 872
rect 582 868 586 872
rect 606 868 610 872
rect 662 868 666 872
rect 678 868 682 872
rect 822 868 826 872
rect 894 868 898 872
rect 942 868 946 872
rect 958 868 962 872
rect 1046 868 1050 872
rect 1102 868 1106 872
rect 1118 868 1122 872
rect 1150 868 1154 872
rect 1206 868 1210 872
rect 1238 868 1242 872
rect 1262 868 1266 872
rect 1270 868 1274 872
rect 1302 868 1306 872
rect 1334 868 1338 872
rect 1422 868 1426 872
rect 1470 868 1474 872
rect 1486 868 1490 872
rect 1542 868 1546 872
rect 1918 878 1922 882
rect 2054 878 2058 882
rect 2518 878 2522 882
rect 2694 878 2698 882
rect 2726 878 2730 882
rect 1670 868 1674 872
rect 1686 868 1690 872
rect 1718 868 1722 872
rect 1782 868 1786 872
rect 1806 866 1810 870
rect 1814 868 1818 872
rect 1902 868 1906 872
rect 1926 868 1930 872
rect 1958 868 1962 872
rect 1974 868 1978 872
rect 2182 868 2186 872
rect 2214 868 2218 872
rect 2342 868 2346 872
rect 2414 868 2418 872
rect 2430 868 2434 872
rect 2534 868 2538 872
rect 2542 868 2546 872
rect 2598 868 2602 872
rect 2646 868 2650 872
rect 2774 868 2778 872
rect 3094 878 3098 882
rect 3406 878 3410 882
rect 3454 878 3458 882
rect 3494 878 3498 882
rect 3750 878 3754 882
rect 2822 868 2826 872
rect 38 858 42 862
rect 62 858 66 862
rect 102 858 106 862
rect 118 858 122 862
rect 134 858 138 862
rect 166 858 170 862
rect 198 858 202 862
rect 238 858 242 862
rect 302 858 306 862
rect 398 858 402 862
rect 422 858 426 862
rect 462 858 466 862
rect 470 858 474 862
rect 494 858 498 862
rect 518 858 522 862
rect 542 858 546 862
rect 550 858 554 862
rect 574 858 578 862
rect 614 858 618 862
rect 654 858 658 862
rect 670 858 674 862
rect 702 858 706 862
rect 758 858 762 862
rect 782 858 786 862
rect 822 858 826 862
rect 886 858 890 862
rect 902 858 906 862
rect 982 858 986 862
rect 1054 858 1058 862
rect 1094 858 1098 862
rect 1142 858 1146 862
rect 1214 858 1218 862
rect 1254 858 1258 862
rect 1326 858 1330 862
rect 1454 858 1458 862
rect 1462 858 1466 862
rect 1478 858 1482 862
rect 1502 858 1506 862
rect 1566 858 1570 862
rect 1630 858 1634 862
rect 1654 858 1658 862
rect 1678 858 1682 862
rect 1686 858 1690 862
rect 1726 858 1730 862
rect 1742 858 1746 862
rect 1854 858 1858 862
rect 1886 859 1890 863
rect 1950 858 1954 862
rect 1982 858 1986 862
rect 2046 858 2050 862
rect 2086 858 2090 862
rect 2118 858 2122 862
rect 2158 858 2162 862
rect 2190 858 2194 862
rect 2206 858 2210 862
rect 2222 858 2226 862
rect 2270 859 2274 863
rect 2302 858 2306 862
rect 2374 858 2378 862
rect 2406 858 2410 862
rect 2454 858 2458 862
rect 2550 858 2554 862
rect 2558 858 2562 862
rect 2582 858 2586 862
rect 2590 858 2594 862
rect 2606 858 2610 862
rect 2654 858 2658 862
rect 2710 858 2714 862
rect 2798 858 2802 862
rect 2806 858 2810 862
rect 2830 858 2834 862
rect 2862 858 2866 862
rect 2934 858 2938 862
rect 2942 858 2946 862
rect 2998 858 3002 862
rect 3038 868 3042 872
rect 3070 868 3074 872
rect 3134 868 3138 872
rect 3270 868 3274 872
rect 3366 868 3370 872
rect 3438 868 3442 872
rect 3462 868 3466 872
rect 3478 868 3482 872
rect 3494 868 3498 872
rect 3542 868 3546 872
rect 3630 868 3634 872
rect 3646 868 3650 872
rect 3710 868 3714 872
rect 3798 868 3802 872
rect 3830 878 3834 882
rect 4094 878 4098 882
rect 4302 878 4306 882
rect 4550 878 4554 882
rect 4734 878 4738 882
rect 4934 878 4938 882
rect 3878 868 3882 872
rect 3910 868 3914 872
rect 3958 868 3962 872
rect 4038 868 4042 872
rect 4078 868 4082 872
rect 4110 868 4114 872
rect 4158 868 4162 872
rect 4214 868 4218 872
rect 4302 868 4306 872
rect 4342 868 4346 872
rect 4454 868 4458 872
rect 4470 868 4474 872
rect 4486 868 4490 872
rect 4502 868 4506 872
rect 4542 868 4546 872
rect 4694 868 4698 872
rect 4766 868 4770 872
rect 4918 868 4922 872
rect 4974 868 4978 872
rect 5014 868 5018 872
rect 5054 868 5058 872
rect 5078 878 5082 882
rect 5150 878 5154 882
rect 5238 878 5242 882
rect 5198 868 5202 872
rect 3022 858 3026 862
rect 3030 858 3034 862
rect 3062 858 3066 862
rect 3078 858 3082 862
rect 3102 858 3106 862
rect 3110 858 3114 862
rect 3142 858 3146 862
rect 3174 859 3178 863
rect 3206 858 3210 862
rect 3310 858 3314 862
rect 3350 858 3354 862
rect 3358 858 3362 862
rect 3390 858 3394 862
rect 3430 858 3434 862
rect 3470 858 3474 862
rect 3542 858 3546 862
rect 3590 858 3594 862
rect 3606 858 3610 862
rect 3654 858 3658 862
rect 3678 858 3682 862
rect 3718 858 3722 862
rect 3734 858 3738 862
rect 3766 858 3770 862
rect 3790 858 3794 862
rect 3806 858 3810 862
rect 3846 858 3850 862
rect 3870 858 3874 862
rect 3902 858 3906 862
rect 3926 858 3930 862
rect 3950 858 3954 862
rect 3966 858 3970 862
rect 4062 859 4066 863
rect 4142 858 4146 862
rect 4150 858 4154 862
rect 4166 858 4170 862
rect 4198 858 4202 862
rect 4206 858 4210 862
rect 4222 858 4226 862
rect 4230 858 4234 862
rect 4254 858 4258 862
rect 4286 858 4290 862
rect 4318 858 4322 862
rect 4358 858 4362 862
rect 4366 858 4370 862
rect 4390 858 4394 862
rect 4398 858 4402 862
rect 4430 858 4434 862
rect 4462 858 4466 862
rect 4478 858 4482 862
rect 4494 858 4498 862
rect 4526 858 4530 862
rect 4598 858 4602 862
rect 4606 858 4610 862
rect 4614 858 4618 862
rect 4638 858 4642 862
rect 4654 858 4658 862
rect 4678 858 4682 862
rect 4718 858 4722 862
rect 4774 858 4778 862
rect 4902 859 4906 863
rect 4998 858 5002 862
rect 5006 858 5010 862
rect 5022 858 5026 862
rect 5046 858 5050 862
rect 5094 858 5098 862
rect 5102 858 5106 862
rect 5134 858 5138 862
rect 5158 858 5162 862
rect 5166 858 5170 862
rect 5190 858 5194 862
rect 5238 858 5242 862
rect 5246 858 5250 862
rect 182 848 186 852
rect 214 848 218 852
rect 222 848 226 852
rect 558 848 562 852
rect 630 848 634 852
rect 862 848 866 852
rect 1078 848 1082 852
rect 1230 848 1234 852
rect 1286 848 1290 852
rect 1494 848 1498 852
rect 1710 848 1714 852
rect 1758 848 1762 852
rect 2174 848 2178 852
rect 2206 848 2210 852
rect 2222 848 2226 852
rect 2390 848 2394 852
rect 2622 848 2626 852
rect 2758 848 2762 852
rect 2982 848 2986 852
rect 3014 848 3018 852
rect 3046 848 3050 852
rect 3486 848 3490 852
rect 3518 848 3522 852
rect 3670 848 3674 852
rect 3854 848 3858 852
rect 3870 848 3874 852
rect 3886 848 3890 852
rect 3934 848 3938 852
rect 4182 848 4186 852
rect 4270 848 4274 852
rect 4286 848 4290 852
rect 5038 848 5042 852
rect 326 838 330 842
rect 830 838 834 842
rect 926 838 930 842
rect 1606 838 1610 842
rect 2238 838 2242 842
rect 2334 838 2338 842
rect 2494 838 2498 842
rect 2974 838 2978 842
rect 3334 838 3338 842
rect 3790 838 3794 842
rect 910 828 914 832
rect 166 818 170 822
rect 350 818 354 822
rect 534 818 538 822
rect 654 818 658 822
rect 1054 818 1058 822
rect 1278 818 1282 822
rect 1518 818 1522 822
rect 1694 818 1698 822
rect 2102 818 2106 822
rect 2134 818 2138 822
rect 3694 818 3698 822
rect 3982 818 3986 822
rect 4414 818 4418 822
rect 4630 818 4634 822
rect 4830 818 4834 822
rect 5126 818 5130 822
rect 330 803 334 807
rect 337 803 341 807
rect 1354 803 1358 807
rect 1361 803 1365 807
rect 2386 803 2390 807
rect 2393 803 2397 807
rect 3402 803 3406 807
rect 3409 803 3413 807
rect 4426 803 4430 807
rect 4433 803 4437 807
rect 502 788 506 792
rect 606 788 610 792
rect 614 788 618 792
rect 750 788 754 792
rect 846 788 850 792
rect 942 788 946 792
rect 974 788 978 792
rect 1134 788 1138 792
rect 1222 788 1226 792
rect 1246 788 1250 792
rect 1390 788 1394 792
rect 1590 788 1594 792
rect 1806 788 1810 792
rect 1838 788 1842 792
rect 2278 788 2282 792
rect 2358 788 2362 792
rect 2446 788 2450 792
rect 2598 788 2602 792
rect 2926 788 2930 792
rect 2958 788 2962 792
rect 3702 788 3706 792
rect 4198 788 4202 792
rect 4390 788 4394 792
rect 4494 788 4498 792
rect 4662 788 4666 792
rect 4966 788 4970 792
rect 5262 788 5266 792
rect 5278 788 5282 792
rect 3318 778 3322 782
rect 3574 778 3578 782
rect 5166 778 5170 782
rect 1118 768 1122 772
rect 1886 768 1890 772
rect 2222 768 2226 772
rect 2566 768 2570 772
rect 2878 768 2882 772
rect 2918 768 2922 772
rect 3094 768 3098 772
rect 3590 768 3594 772
rect 3918 768 3922 772
rect 4294 768 4298 772
rect 4806 768 4810 772
rect 4926 768 4930 772
rect 5126 768 5130 772
rect 206 758 210 762
rect 510 758 514 762
rect 734 758 738 762
rect 958 758 962 762
rect 30 748 34 752
rect 150 748 154 752
rect 206 748 210 752
rect 222 748 226 752
rect 270 748 274 752
rect 350 748 354 752
rect 366 748 370 752
rect 374 748 378 752
rect 414 748 418 752
rect 446 748 450 752
rect 470 748 474 752
rect 486 748 490 752
rect 542 747 546 751
rect 566 748 570 752
rect 646 748 650 752
rect 654 748 658 752
rect 710 748 714 752
rect 750 748 754 752
rect 766 748 770 752
rect 798 748 802 752
rect 822 748 826 752
rect 830 748 834 752
rect 854 748 858 752
rect 982 748 986 752
rect 998 748 1002 752
rect 1006 748 1010 752
rect 1022 758 1026 762
rect 1142 758 1146 762
rect 1206 758 1210 762
rect 1286 758 1290 762
rect 1326 758 1330 762
rect 1742 758 1746 762
rect 1070 747 1074 751
rect 1166 748 1170 752
rect 1190 748 1194 752
rect 1198 748 1202 752
rect 1222 748 1226 752
rect 1238 748 1242 752
rect 1270 748 1274 752
rect 1294 748 1298 752
rect 1342 748 1346 752
rect 1366 748 1370 752
rect 1398 748 1402 752
rect 1406 748 1410 752
rect 1414 748 1418 752
rect 1422 748 1426 752
rect 1534 748 1538 752
rect 1574 748 1578 752
rect 1606 748 1610 752
rect 1614 748 1618 752
rect 1654 748 1658 752
rect 1726 748 1730 752
rect 2302 758 2306 762
rect 2318 758 2322 762
rect 2342 758 2346 762
rect 1766 748 1770 752
rect 1782 748 1786 752
rect 1822 748 1826 752
rect 1838 748 1842 752
rect 1886 748 1890 752
rect 1926 748 1930 752
rect 1958 747 1962 751
rect 1990 748 1994 752
rect 2038 748 2042 752
rect 2046 748 2050 752
rect 2070 748 2074 752
rect 2094 748 2098 752
rect 2110 748 2114 752
rect 2158 747 2162 751
rect 2230 748 2234 752
rect 2262 748 2266 752
rect 2278 748 2282 752
rect 2286 748 2290 752
rect 2302 748 2306 752
rect 2326 748 2330 752
rect 2382 748 2386 752
rect 2398 748 2402 752
rect 2422 748 2426 752
rect 2430 748 2434 752
rect 2446 748 2450 752
rect 2470 758 2474 762
rect 2638 758 2642 762
rect 2862 758 2866 762
rect 2934 758 2938 762
rect 2990 758 2994 762
rect 3022 758 3026 762
rect 3078 758 3082 762
rect 3438 758 3442 762
rect 2542 748 2546 752
rect 2614 748 2618 752
rect 2630 748 2634 752
rect 2638 748 2642 752
rect 2654 748 2658 752
rect 6 738 10 742
rect 38 738 42 742
rect 102 738 106 742
rect 118 738 122 742
rect 230 738 234 742
rect 262 738 266 742
rect 422 738 426 742
rect 486 738 490 742
rect 526 738 530 742
rect 710 738 714 742
rect 758 738 762 742
rect 774 738 778 742
rect 886 738 890 742
rect 982 738 986 742
rect 990 738 994 742
rect 1038 738 1042 742
rect 1054 738 1058 742
rect 1230 738 1234 742
rect 1262 738 1266 742
rect 1454 738 1458 742
rect 1486 738 1490 742
rect 1630 738 1634 742
rect 1718 738 1722 742
rect 1750 738 1754 742
rect 1782 738 1786 742
rect 1790 738 1794 742
rect 1814 738 1818 742
rect 1846 738 1850 742
rect 1854 738 1858 742
rect 1998 738 2002 742
rect 2070 738 2074 742
rect 2086 738 2090 742
rect 2142 738 2146 742
rect 2246 738 2250 742
rect 2254 738 2258 742
rect 2286 738 2290 742
rect 2734 747 2738 751
rect 2782 748 2786 752
rect 2814 748 2818 752
rect 2822 748 2826 752
rect 2838 748 2842 752
rect 2854 748 2858 752
rect 2902 748 2906 752
rect 2926 748 2930 752
rect 2950 748 2954 752
rect 2974 748 2978 752
rect 2982 748 2986 752
rect 3038 748 3042 752
rect 3062 748 3066 752
rect 3166 747 3170 751
rect 3206 748 3210 752
rect 3214 748 3218 752
rect 3230 748 3234 752
rect 3238 748 3242 752
rect 3310 748 3314 752
rect 3350 748 3354 752
rect 3382 747 3386 751
rect 3438 748 3442 752
rect 3462 758 3466 762
rect 3798 758 3802 762
rect 3974 758 3978 762
rect 4030 758 4034 762
rect 4038 758 4042 762
rect 4054 758 4058 762
rect 4070 758 4074 762
rect 4166 758 4170 762
rect 4414 758 4418 762
rect 4598 758 4602 762
rect 4950 758 4954 762
rect 3478 748 3482 752
rect 3494 748 3498 752
rect 3534 748 3538 752
rect 3566 748 3570 752
rect 3606 748 3610 752
rect 3614 748 3618 752
rect 3678 748 3682 752
rect 3694 748 3698 752
rect 3734 748 3738 752
rect 3766 747 3770 751
rect 3814 748 3818 752
rect 3862 748 3866 752
rect 3950 748 3954 752
rect 3958 748 3962 752
rect 3966 748 3970 752
rect 3990 748 3994 752
rect 3998 748 4002 752
rect 4014 748 4018 752
rect 4062 748 4066 752
rect 4086 748 4090 752
rect 4102 748 4106 752
rect 4110 748 4114 752
rect 4174 748 4178 752
rect 4182 748 4186 752
rect 4238 748 4242 752
rect 4334 748 4338 752
rect 4350 748 4354 752
rect 4390 748 4394 752
rect 4430 748 4434 752
rect 4454 748 4458 752
rect 4462 748 4466 752
rect 2366 738 2370 742
rect 2438 738 2442 742
rect 2486 738 2490 742
rect 2502 738 2506 742
rect 2622 738 2626 742
rect 2662 738 2666 742
rect 2726 738 2730 742
rect 2790 738 2794 742
rect 2854 738 2858 742
rect 2886 738 2890 742
rect 3014 738 3018 742
rect 3046 738 3050 742
rect 3054 738 3058 742
rect 3182 738 3186 742
rect 3246 738 3250 742
rect 3422 738 3426 742
rect 3430 738 3434 742
rect 3494 738 3498 742
rect 3558 738 3562 742
rect 3670 738 3674 742
rect 3798 738 3802 742
rect 3822 738 3826 742
rect 3870 738 3874 742
rect 3942 738 3946 742
rect 3998 738 4002 742
rect 4558 747 4562 751
rect 4718 748 4722 752
rect 4774 748 4778 752
rect 4806 748 4810 752
rect 4822 748 4826 752
rect 4870 748 4874 752
rect 4966 748 4970 752
rect 4982 748 4986 752
rect 5014 748 5018 752
rect 5022 748 5026 752
rect 5038 758 5042 762
rect 5054 748 5058 752
rect 5070 748 5074 752
rect 5110 748 5114 752
rect 5150 758 5154 762
rect 5158 748 5162 752
rect 5222 748 5226 752
rect 4062 738 4066 742
rect 4094 738 4098 742
rect 4142 738 4146 742
rect 4190 738 4194 742
rect 4278 738 4282 742
rect 4422 738 4426 742
rect 4446 738 4450 742
rect 4654 738 4658 742
rect 4758 738 4762 742
rect 4790 738 4794 742
rect 4798 738 4802 742
rect 4830 738 4834 742
rect 4870 738 4874 742
rect 5006 738 5010 742
rect 5062 738 5066 742
rect 5094 738 5098 742
rect 5158 738 5162 742
rect 5246 738 5250 742
rect 462 728 466 732
rect 470 728 474 732
rect 726 728 730 732
rect 814 728 818 732
rect 1142 728 1146 732
rect 1238 728 1242 732
rect 1254 728 1258 732
rect 1310 728 1314 732
rect 1542 728 1546 732
rect 1806 728 1810 732
rect 1854 728 1858 732
rect 2006 728 2010 732
rect 2022 728 2026 732
rect 2126 728 2130 732
rect 2246 728 2250 732
rect 2326 728 2330 732
rect 2606 728 2610 732
rect 2702 728 2706 732
rect 2766 728 2770 732
rect 2830 728 2834 732
rect 2990 728 2994 732
rect 3078 728 3082 732
rect 3510 728 3514 732
rect 3518 728 3522 732
rect 3550 728 3554 732
rect 3974 728 3978 732
rect 4158 728 4162 732
rect 4406 728 4410 732
rect 4510 728 4514 732
rect 4558 728 4562 732
rect 4790 728 4794 732
rect 4998 728 5002 732
rect 5270 728 5274 732
rect 5286 728 5290 732
rect 198 718 202 722
rect 382 718 386 722
rect 430 718 434 722
rect 782 718 786 722
rect 1174 718 1178 722
rect 1286 718 1290 722
rect 1302 718 1306 722
rect 1710 718 1714 722
rect 2406 718 2410 722
rect 3502 718 3506 722
rect 4030 718 4034 722
rect 4070 718 4074 722
rect 4478 718 4482 722
rect 5086 718 5090 722
rect 850 703 854 707
rect 857 703 861 707
rect 1874 703 1878 707
rect 1881 703 1885 707
rect 2890 703 2894 707
rect 2897 703 2901 707
rect 3922 703 3926 707
rect 3929 703 3933 707
rect 4938 703 4942 707
rect 4945 703 4949 707
rect 174 688 178 692
rect 214 688 218 692
rect 486 688 490 692
rect 494 688 498 692
rect 614 688 618 692
rect 638 688 642 692
rect 718 688 722 692
rect 734 688 738 692
rect 838 688 842 692
rect 942 688 946 692
rect 958 688 962 692
rect 1078 688 1082 692
rect 1182 688 1186 692
rect 1350 688 1354 692
rect 1462 688 1466 692
rect 1502 688 1506 692
rect 1606 688 1610 692
rect 1806 688 1810 692
rect 1966 688 1970 692
rect 2062 688 2066 692
rect 2238 688 2242 692
rect 2270 688 2274 692
rect 2454 688 2458 692
rect 2510 688 2514 692
rect 2838 688 2842 692
rect 2886 688 2890 692
rect 3078 688 3082 692
rect 3206 688 3210 692
rect 3334 688 3338 692
rect 3486 688 3490 692
rect 3814 688 3818 692
rect 3886 688 3890 692
rect 4094 688 4098 692
rect 4118 688 4122 692
rect 4214 688 4218 692
rect 4334 688 4338 692
rect 4438 688 4442 692
rect 4574 688 4578 692
rect 4654 688 4658 692
rect 4694 688 4698 692
rect 4878 688 4882 692
rect 4942 688 4946 692
rect 4982 688 4986 692
rect 5198 688 5202 692
rect 62 678 66 682
rect 134 678 138 682
rect 182 678 186 682
rect 222 678 226 682
rect 670 678 674 682
rect 678 678 682 682
rect 878 678 882 682
rect 1070 678 1074 682
rect 1430 678 1434 682
rect 1510 678 1514 682
rect 1542 678 1546 682
rect 1678 678 1682 682
rect 1686 678 1690 682
rect 1758 678 1762 682
rect 1846 678 1850 682
rect 2142 678 2146 682
rect 2318 678 2322 682
rect 2502 678 2506 682
rect 2574 678 2578 682
rect 70 668 74 672
rect 126 668 130 672
rect 206 668 210 672
rect 230 668 234 672
rect 262 668 266 672
rect 294 668 298 672
rect 366 668 370 672
rect 390 668 394 672
rect 518 668 522 672
rect 534 668 538 672
rect 630 668 634 672
rect 726 668 730 672
rect 758 668 762 672
rect 886 668 890 672
rect 974 668 978 672
rect 1062 668 1066 672
rect 1190 668 1194 672
rect 1286 668 1290 672
rect 1486 668 1490 672
rect 1638 668 1642 672
rect 1646 668 1650 672
rect 1670 668 1674 672
rect 1774 668 1778 672
rect 1902 668 1906 672
rect 1958 668 1962 672
rect 2046 668 2050 672
rect 2086 668 2090 672
rect 2678 678 2682 682
rect 2878 678 2882 682
rect 3150 678 3154 682
rect 3270 678 3274 682
rect 2190 668 2194 672
rect 2230 668 2234 672
rect 2262 668 2266 672
rect 2294 668 2298 672
rect 2366 668 2370 672
rect 2422 668 2426 672
rect 2438 668 2442 672
rect 2446 668 2450 672
rect 2606 668 2610 672
rect 2630 668 2634 672
rect 2646 668 2650 672
rect 2686 668 2690 672
rect 14 658 18 662
rect 38 658 42 662
rect 46 658 50 662
rect 62 658 66 662
rect 78 658 82 662
rect 118 658 122 662
rect 158 658 162 662
rect 198 658 202 662
rect 238 658 242 662
rect 270 658 274 662
rect 302 658 306 662
rect 358 658 362 662
rect 390 658 394 662
rect 430 658 434 662
rect 446 658 450 662
rect 510 658 514 662
rect 558 658 562 662
rect 622 658 626 662
rect 654 658 658 662
rect 702 658 706 662
rect 782 658 786 662
rect 862 658 866 662
rect 1006 658 1010 662
rect 1014 658 1018 662
rect 1046 658 1050 662
rect 1054 658 1058 662
rect 1118 658 1122 662
rect 1142 659 1146 663
rect 1206 658 1210 662
rect 1214 658 1218 662
rect 1230 658 1234 662
rect 1238 658 1242 662
rect 1270 659 1274 663
rect 1374 658 1378 662
rect 1382 658 1386 662
rect 1446 658 1450 662
rect 1494 658 1498 662
rect 1558 658 1562 662
rect 1574 658 1578 662
rect 1622 658 1626 662
rect 1630 658 1634 662
rect 1662 658 1666 662
rect 1718 658 1722 662
rect 1782 658 1786 662
rect 1822 658 1826 662
rect 1854 658 1858 662
rect 1910 658 1914 662
rect 1950 658 1954 662
rect 2022 658 2026 662
rect 2078 658 2082 662
rect 2166 658 2170 662
rect 2222 658 2226 662
rect 2254 658 2258 662
rect 2294 658 2298 662
rect 2358 658 2362 662
rect 2430 658 2434 662
rect 2454 658 2458 662
rect 2470 658 2474 662
rect 2486 658 2490 662
rect 2574 659 2578 663
rect 2726 668 2730 672
rect 2814 668 2818 672
rect 2622 658 2626 662
rect 2654 658 2658 662
rect 2662 658 2666 662
rect 2694 658 2698 662
rect 2710 658 2714 662
rect 2742 659 2746 663
rect 2870 668 2874 672
rect 2918 668 2922 672
rect 2926 668 2930 672
rect 2958 668 2962 672
rect 3014 668 3018 672
rect 3110 668 3114 672
rect 3142 668 3146 672
rect 3190 668 3194 672
rect 3454 678 3458 682
rect 3526 678 3530 682
rect 3558 678 3562 682
rect 4102 678 4106 682
rect 4110 678 4114 682
rect 4222 678 4226 682
rect 4318 678 4322 682
rect 4510 678 4514 682
rect 4542 678 4546 682
rect 4854 678 4858 682
rect 4990 678 4994 682
rect 4998 678 5002 682
rect 3390 668 3394 672
rect 3414 668 3418 672
rect 3430 668 3434 672
rect 3446 668 3450 672
rect 3454 668 3458 672
rect 3534 668 3538 672
rect 3646 668 3650 672
rect 3686 668 3690 672
rect 3718 668 3722 672
rect 3846 668 3850 672
rect 3870 668 3874 672
rect 3926 668 3930 672
rect 3974 668 3978 672
rect 3990 668 3994 672
rect 4022 668 4026 672
rect 4054 668 4058 672
rect 4086 668 4090 672
rect 4126 668 4130 672
rect 4142 668 4146 672
rect 4198 668 4202 672
rect 4230 668 4234 672
rect 4294 668 4298 672
rect 4390 668 4394 672
rect 4398 668 4402 672
rect 4582 668 4586 672
rect 2822 658 2826 662
rect 2846 658 2850 662
rect 2862 658 2866 662
rect 2902 658 2906 662
rect 2910 658 2914 662
rect 2966 658 2970 662
rect 3022 658 3026 662
rect 3110 658 3114 662
rect 3118 658 3122 662
rect 3134 658 3138 662
rect 3166 658 3170 662
rect 3182 658 3186 662
rect 3198 658 3202 662
rect 3262 658 3266 662
rect 3302 658 3306 662
rect 3358 658 3362 662
rect 3366 658 3370 662
rect 3406 658 3410 662
rect 3438 658 3442 662
rect 3478 658 3482 662
rect 3502 658 3506 662
rect 3510 658 3514 662
rect 3542 658 3546 662
rect 3622 658 3626 662
rect 3678 658 3682 662
rect 3694 658 3698 662
rect 3710 658 3714 662
rect 3758 658 3762 662
rect 3782 658 3786 662
rect 3862 658 3866 662
rect 3958 659 3962 663
rect 3998 658 4002 662
rect 4030 658 4034 662
rect 4054 658 4058 662
rect 4086 658 4090 662
rect 4134 658 4138 662
rect 4150 658 4154 662
rect 4190 658 4194 662
rect 4206 658 4210 662
rect 4302 658 4306 662
rect 4398 658 4402 662
rect 4414 658 4418 662
rect 4478 658 4482 662
rect 4494 658 4498 662
rect 4558 658 4562 662
rect 4590 658 4594 662
rect 4598 658 4602 662
rect 4614 658 4618 662
rect 4630 668 4634 672
rect 4662 668 4666 672
rect 4670 668 4674 672
rect 4758 668 4762 672
rect 4910 668 4914 672
rect 4958 668 4962 672
rect 5006 668 5010 672
rect 5062 668 5066 672
rect 5150 668 5154 672
rect 5166 668 5170 672
rect 5246 668 5250 672
rect 4630 658 4634 662
rect 4638 658 4642 662
rect 4654 658 4658 662
rect 4678 658 4682 662
rect 4702 658 4706 662
rect 4710 658 4714 662
rect 4742 658 4746 662
rect 4790 658 4794 662
rect 4806 658 4810 662
rect 4894 658 4898 662
rect 4902 658 4906 662
rect 4918 658 4922 662
rect 4966 658 4970 662
rect 5014 658 5018 662
rect 5046 658 5050 662
rect 5054 658 5058 662
rect 5118 658 5122 662
rect 5166 658 5170 662
rect 5182 658 5186 662
rect 5254 658 5258 662
rect 102 648 106 652
rect 174 648 178 652
rect 254 648 258 652
rect 374 648 378 652
rect 494 648 498 652
rect 718 648 722 652
rect 742 648 746 652
rect 1470 648 1474 652
rect 1614 648 1618 652
rect 1646 648 1650 652
rect 1702 648 1706 652
rect 1798 648 1802 652
rect 1806 648 1810 652
rect 1926 648 1930 652
rect 1950 648 1954 652
rect 2062 648 2066 652
rect 2126 648 2130 652
rect 2206 648 2210 652
rect 2238 648 2242 652
rect 2270 648 2274 652
rect 2414 648 2418 652
rect 2710 648 2714 652
rect 2838 648 2842 652
rect 2846 648 2850 652
rect 2950 648 2954 652
rect 2966 648 2970 652
rect 2982 648 2986 652
rect 3102 648 3106 652
rect 3118 648 3122 652
rect 3662 648 3666 652
rect 3678 648 3682 652
rect 3694 648 3698 652
rect 3838 648 3842 652
rect 4014 648 4018 652
rect 4030 648 4034 652
rect 4078 648 4082 652
rect 4166 648 4170 652
rect 4422 648 4426 652
rect 4598 648 4602 652
rect 4694 648 4698 652
rect 4942 648 4946 652
rect 4982 648 4986 652
rect 5030 648 5034 652
rect 270 638 274 642
rect 286 638 290 642
rect 334 638 338 642
rect 958 638 962 642
rect 1174 638 1178 642
rect 2222 638 2226 642
rect 3566 638 3570 642
rect 4310 638 4314 642
rect 5070 638 5074 642
rect 30 618 34 622
rect 78 618 82 622
rect 190 618 194 622
rect 238 618 242 622
rect 358 618 362 622
rect 862 618 866 622
rect 990 618 994 622
rect 1038 618 1042 622
rect 1398 618 1402 622
rect 1742 618 1746 622
rect 1766 618 1770 622
rect 1782 618 1786 622
rect 2094 618 2098 622
rect 2670 618 2674 622
rect 2934 618 2938 622
rect 3302 618 3306 622
rect 3486 618 3490 622
rect 3550 618 3554 622
rect 3998 618 4002 622
rect 4094 618 4098 622
rect 4190 618 4194 622
rect 4214 618 4218 622
rect 4334 618 4338 622
rect 4726 618 4730 622
rect 330 603 334 607
rect 337 603 341 607
rect 1354 603 1358 607
rect 1361 603 1365 607
rect 2386 603 2390 607
rect 2393 603 2397 607
rect 3402 603 3406 607
rect 3409 603 3413 607
rect 4426 603 4430 607
rect 4433 603 4437 607
rect 94 588 98 592
rect 190 588 194 592
rect 462 588 466 592
rect 494 588 498 592
rect 542 588 546 592
rect 646 588 650 592
rect 662 588 666 592
rect 806 588 810 592
rect 910 588 914 592
rect 1054 588 1058 592
rect 1174 588 1178 592
rect 1278 588 1282 592
rect 1494 588 1498 592
rect 1814 588 1818 592
rect 1838 588 1842 592
rect 2006 588 2010 592
rect 2038 588 2042 592
rect 2110 588 2114 592
rect 2406 588 2410 592
rect 2454 588 2458 592
rect 2494 588 2498 592
rect 2862 588 2866 592
rect 3078 588 3082 592
rect 3182 588 3186 592
rect 3518 588 3522 592
rect 3582 588 3586 592
rect 3614 588 3618 592
rect 3630 588 3634 592
rect 4054 588 4058 592
rect 4302 588 4306 592
rect 4622 588 4626 592
rect 4750 588 4754 592
rect 4870 588 4874 592
rect 4934 588 4938 592
rect 5006 588 5010 592
rect 5038 588 5042 592
rect 5102 588 5106 592
rect 766 578 770 582
rect 1678 578 1682 582
rect 2662 578 2666 582
rect 3854 578 3858 582
rect 870 568 874 572
rect 894 568 898 572
rect 1606 568 1610 572
rect 1782 568 1786 572
rect 1950 568 1954 572
rect 2182 568 2186 572
rect 2198 568 2202 572
rect 2438 568 2442 572
rect 2510 568 2514 572
rect 2902 568 2906 572
rect 3998 568 4002 572
rect 4206 568 4210 572
rect 4222 568 4226 572
rect 5206 568 5210 572
rect 534 558 538 562
rect 670 558 674 562
rect 822 558 826 562
rect 854 558 858 562
rect 926 558 930 562
rect 1046 558 1050 562
rect 1294 558 1298 562
rect 1326 558 1330 562
rect 1350 558 1354 562
rect 1398 558 1402 562
rect 30 547 34 551
rect 126 547 130 551
rect 230 548 234 552
rect 310 548 314 552
rect 318 548 322 552
rect 342 548 346 552
rect 350 548 354 552
rect 398 547 402 551
rect 494 548 498 552
rect 582 547 586 551
rect 710 548 714 552
rect 734 548 738 552
rect 790 548 794 552
rect 806 548 810 552
rect 838 548 842 552
rect 846 548 850 552
rect 902 548 906 552
rect 950 548 954 552
rect 982 548 986 552
rect 1014 548 1018 552
rect 1022 548 1026 552
rect 1094 548 1098 552
rect 1150 548 1154 552
rect 1230 548 1234 552
rect 1278 548 1282 552
rect 1310 548 1314 552
rect 1334 548 1338 552
rect 1366 548 1370 552
rect 1382 548 1386 552
rect 1390 548 1394 552
rect 1430 547 1434 551
rect 1510 548 1514 552
rect 1534 558 1538 562
rect 1590 558 1594 562
rect 1622 558 1626 562
rect 1654 558 1658 562
rect 1550 548 1554 552
rect 1574 548 1578 552
rect 1606 548 1610 552
rect 1622 548 1626 552
rect 1638 548 1642 552
rect 1862 558 1866 562
rect 1966 558 1970 562
rect 1990 558 1994 562
rect 2022 558 2026 562
rect 2054 558 2058 562
rect 2142 558 2146 562
rect 1678 548 1682 552
rect 110 538 114 542
rect 206 538 210 542
rect 238 538 242 542
rect 310 538 314 542
rect 382 538 386 542
rect 518 538 522 542
rect 566 538 570 542
rect 654 538 658 542
rect 798 538 802 542
rect 830 538 834 542
rect 894 538 898 542
rect 902 538 906 542
rect 974 538 978 542
rect 1030 538 1034 542
rect 1230 538 1234 542
rect 1270 538 1274 542
rect 1302 538 1306 542
rect 1334 538 1338 542
rect 1374 538 1378 542
rect 1502 538 1506 542
rect 1558 538 1562 542
rect 1566 538 1570 542
rect 1598 538 1602 542
rect 1718 547 1722 551
rect 1822 548 1826 552
rect 1838 548 1842 552
rect 1902 548 1906 552
rect 1926 548 1930 552
rect 1982 548 1986 552
rect 2022 548 2026 552
rect 2038 548 2042 552
rect 2070 548 2074 552
rect 2086 548 2090 552
rect 2118 548 2122 552
rect 2302 558 2306 562
rect 2478 558 2482 562
rect 3038 558 3042 562
rect 2174 548 2178 552
rect 2238 548 2242 552
rect 2278 548 2282 552
rect 2302 548 2306 552
rect 1686 538 1690 542
rect 1806 538 1810 542
rect 1830 538 1834 542
rect 1894 538 1898 542
rect 1934 538 1938 542
rect 2014 538 2018 542
rect 2046 538 2050 542
rect 2078 538 2082 542
rect 2094 538 2098 542
rect 2110 538 2114 542
rect 2158 538 2162 542
rect 2174 538 2178 542
rect 2262 538 2266 542
rect 2278 538 2282 542
rect 2334 547 2338 551
rect 2366 548 2370 552
rect 2438 548 2442 552
rect 2446 548 2450 552
rect 2502 548 2506 552
rect 2574 547 2578 551
rect 2622 548 2626 552
rect 2654 548 2658 552
rect 2726 547 2730 551
rect 2758 548 2762 552
rect 2774 548 2778 552
rect 2806 548 2810 552
rect 2822 548 2826 552
rect 2846 548 2850 552
rect 2854 548 2858 552
rect 2886 548 2890 552
rect 2982 548 2986 552
rect 3558 558 3562 562
rect 3566 558 3570 562
rect 3694 558 3698 562
rect 3886 558 3890 562
rect 3958 558 3962 562
rect 4998 558 5002 562
rect 5086 558 5090 562
rect 3062 548 3066 552
rect 3134 548 3138 552
rect 3182 548 3186 552
rect 3230 548 3234 552
rect 3294 548 3298 552
rect 3310 548 3314 552
rect 3374 548 3378 552
rect 3454 548 3458 552
rect 3502 548 3506 552
rect 3526 548 3530 552
rect 3534 548 3538 552
rect 3590 548 3594 552
rect 3598 548 3602 552
rect 3654 548 3658 552
rect 3662 548 3666 552
rect 3702 548 3706 552
rect 3790 547 3794 551
rect 3870 548 3874 552
rect 3878 548 3882 552
rect 3886 548 3890 552
rect 3902 548 3906 552
rect 3950 548 3954 552
rect 3974 548 3978 552
rect 3998 548 4002 552
rect 4014 548 4018 552
rect 4030 548 4034 552
rect 4110 548 4114 552
rect 4166 548 4170 552
rect 4198 548 4202 552
rect 4246 548 4250 552
rect 4334 548 4338 552
rect 4342 548 4346 552
rect 4470 548 4474 552
rect 4510 548 4514 552
rect 4566 548 4570 552
rect 4590 548 4594 552
rect 4598 548 4602 552
rect 4678 548 4682 552
rect 4718 548 4722 552
rect 4806 548 4810 552
rect 4934 548 4938 552
rect 4982 548 4986 552
rect 5030 548 5034 552
rect 5062 548 5066 552
rect 5102 548 5106 552
rect 5150 548 5154 552
rect 5158 548 5162 552
rect 5190 558 5194 562
rect 5246 548 5250 552
rect 5270 548 5274 552
rect 2318 538 2322 542
rect 2446 538 2450 542
rect 2502 538 2506 542
rect 2558 538 2562 542
rect 2606 538 2610 542
rect 2630 538 2634 542
rect 2646 538 2650 542
rect 2742 538 2746 542
rect 2766 538 2770 542
rect 2894 538 2898 542
rect 3006 538 3010 542
rect 3022 538 3026 542
rect 3038 538 3042 542
rect 3070 538 3074 542
rect 3126 538 3130 542
rect 3174 538 3178 542
rect 3222 538 3226 542
rect 3238 538 3242 542
rect 3462 538 3466 542
rect 3534 538 3538 542
rect 3590 538 3594 542
rect 3646 538 3650 542
rect 3686 538 3690 542
rect 3718 538 3722 542
rect 3782 538 3786 542
rect 3822 538 3826 542
rect 3918 538 3922 542
rect 3950 538 3954 542
rect 3966 538 3970 542
rect 3982 538 3986 542
rect 3990 538 3994 542
rect 4022 538 4026 542
rect 4134 538 4138 542
rect 4190 538 4194 542
rect 4286 538 4290 542
rect 4478 538 4482 542
rect 4518 538 4522 542
rect 4526 538 4530 542
rect 4702 538 4706 542
rect 30 528 34 532
rect 62 528 66 532
rect 550 528 554 532
rect 934 528 938 532
rect 1046 528 1050 532
rect 1118 528 1122 532
rect 1150 528 1154 532
rect 1430 528 1434 532
rect 1718 528 1722 532
rect 1790 528 1794 532
rect 1806 528 1810 532
rect 1878 528 1882 532
rect 1910 528 1914 532
rect 1950 528 1954 532
rect 2110 528 2114 532
rect 2470 528 2474 532
rect 2790 528 2794 532
rect 2838 528 2842 532
rect 2862 528 2866 532
rect 3206 528 3210 532
rect 3366 528 3370 532
rect 3486 528 3490 532
rect 3502 528 3506 532
rect 3630 528 3634 532
rect 3934 528 3938 532
rect 4030 528 4034 532
rect 4046 528 4050 532
rect 4150 528 4154 532
rect 4182 528 4186 532
rect 4446 528 4450 532
rect 4542 528 4546 532
rect 4926 538 4930 542
rect 4974 538 4978 542
rect 5022 538 5026 542
rect 5054 538 5058 542
rect 5062 538 5066 542
rect 5086 538 5090 542
rect 5094 538 5098 542
rect 5142 538 5146 542
rect 5158 538 5162 542
rect 5190 538 5194 542
rect 5206 538 5210 542
rect 4798 528 4802 532
rect 4830 528 4834 532
rect 4958 528 4962 532
rect 5006 528 5010 532
rect 5038 528 5042 532
rect 5126 528 5130 532
rect 782 518 786 522
rect 966 518 970 522
rect 998 518 1002 522
rect 1526 518 1530 522
rect 1590 518 1594 522
rect 1886 518 1890 522
rect 1918 518 1922 522
rect 2054 518 2058 522
rect 3078 518 3082 522
rect 3326 518 3330 522
rect 3430 518 3434 522
rect 3470 518 3474 522
rect 3558 518 3562 522
rect 3726 518 3730 522
rect 4574 518 4578 522
rect 4606 518 4610 522
rect 4734 518 4738 522
rect 4998 518 5002 522
rect 850 503 854 507
rect 857 503 861 507
rect 1874 503 1878 507
rect 1881 503 1885 507
rect 2890 503 2894 507
rect 2897 503 2901 507
rect 3922 503 3926 507
rect 3929 503 3933 507
rect 4938 503 4942 507
rect 4945 503 4949 507
rect 190 488 194 492
rect 302 488 306 492
rect 326 488 330 492
rect 646 488 650 492
rect 662 488 666 492
rect 694 488 698 492
rect 766 488 770 492
rect 846 488 850 492
rect 1006 488 1010 492
rect 1262 488 1266 492
rect 1294 488 1298 492
rect 1470 488 1474 492
rect 1566 488 1570 492
rect 1662 488 1666 492
rect 1670 488 1674 492
rect 2166 488 2170 492
rect 2182 488 2186 492
rect 2462 488 2466 492
rect 2574 488 2578 492
rect 2726 488 2730 492
rect 2966 488 2970 492
rect 3150 488 3154 492
rect 3782 488 3786 492
rect 3806 488 3810 492
rect 4046 488 4050 492
rect 4438 488 4442 492
rect 4630 488 4634 492
rect 4654 488 4658 492
rect 4686 488 4690 492
rect 4766 488 4770 492
rect 4774 488 4778 492
rect 5038 488 5042 492
rect 5158 488 5162 492
rect 5166 488 5170 492
rect 5270 488 5274 492
rect 30 478 34 482
rect 238 478 242 482
rect 318 468 322 472
rect 342 478 346 482
rect 502 478 506 482
rect 702 478 706 482
rect 1150 478 1154 482
rect 1214 478 1218 482
rect 1358 478 1362 482
rect 1534 478 1538 482
rect 1734 478 1738 482
rect 1750 478 1754 482
rect 1774 478 1778 482
rect 382 468 386 472
rect 446 468 450 472
rect 542 468 546 472
rect 566 468 570 472
rect 670 468 674 472
rect 686 468 690 472
rect 702 468 706 472
rect 774 468 778 472
rect 894 468 898 472
rect 982 468 986 472
rect 1110 468 1114 472
rect 1126 468 1130 472
rect 1270 468 1274 472
rect 46 458 50 462
rect 62 458 66 462
rect 118 458 122 462
rect 126 458 130 462
rect 150 458 154 462
rect 166 458 170 462
rect 174 458 178 462
rect 198 458 202 462
rect 246 458 250 462
rect 310 458 314 462
rect 374 458 378 462
rect 454 458 458 462
rect 486 458 490 462
rect 494 458 498 462
rect 518 458 522 462
rect 534 458 538 462
rect 550 458 554 462
rect 582 459 586 463
rect 678 458 682 462
rect 718 458 722 462
rect 742 458 746 462
rect 750 458 754 462
rect 774 458 778 462
rect 814 458 818 462
rect 822 458 826 462
rect 910 459 914 463
rect 942 458 946 462
rect 950 458 954 462
rect 1038 458 1042 462
rect 1062 458 1066 462
rect 1102 458 1106 462
rect 1134 458 1138 462
rect 1182 459 1186 463
rect 1214 458 1218 462
rect 1270 458 1274 462
rect 1334 468 1338 472
rect 1422 468 1426 472
rect 1430 468 1434 472
rect 1486 468 1490 472
rect 1582 468 1586 472
rect 1694 468 1698 472
rect 1726 468 1730 472
rect 1862 468 1866 472
rect 1870 468 1874 472
rect 1902 478 1906 482
rect 2030 478 2034 482
rect 2078 478 2082 482
rect 1918 468 1922 472
rect 1942 468 1946 472
rect 1958 468 1962 472
rect 1974 468 1978 472
rect 1990 468 1994 472
rect 1998 468 2002 472
rect 2014 468 2018 472
rect 2078 468 2082 472
rect 2094 468 2098 472
rect 2110 468 2114 472
rect 2174 468 2178 472
rect 2262 468 2266 472
rect 2278 468 2282 472
rect 2334 468 2338 472
rect 2366 468 2370 472
rect 2374 468 2378 472
rect 2390 468 2394 472
rect 2422 468 2426 472
rect 2974 478 2978 482
rect 3526 478 3530 482
rect 3542 478 3546 482
rect 3790 478 3794 482
rect 2558 468 2562 472
rect 2670 468 2674 472
rect 2694 468 2698 472
rect 2710 468 2714 472
rect 2846 468 2850 472
rect 2878 468 2882 472
rect 2958 468 2962 472
rect 2982 468 2986 472
rect 2998 468 3002 472
rect 3094 468 3098 472
rect 3158 468 3162 472
rect 3174 468 3178 472
rect 3214 468 3218 472
rect 3278 468 3282 472
rect 3310 468 3314 472
rect 3318 468 3322 472
rect 3350 468 3354 472
rect 3382 468 3386 472
rect 3526 468 3530 472
rect 3542 468 3546 472
rect 3606 468 3610 472
rect 3710 468 3714 472
rect 3742 468 3746 472
rect 3766 468 3770 472
rect 3790 468 3794 472
rect 3830 478 3834 482
rect 3854 478 3858 482
rect 4006 478 4010 482
rect 3902 468 3906 472
rect 3926 468 3930 472
rect 3982 468 3986 472
rect 4174 478 4178 482
rect 4334 478 4338 482
rect 4406 478 4410 482
rect 4590 478 4594 482
rect 4622 478 4626 482
rect 4894 478 4898 482
rect 5126 478 5130 482
rect 5262 478 5266 482
rect 4030 468 4034 472
rect 4126 468 4130 472
rect 4142 468 4146 472
rect 4190 468 4194 472
rect 4230 468 4234 472
rect 4254 468 4258 472
rect 4374 468 4378 472
rect 4454 468 4458 472
rect 4518 468 4522 472
rect 4638 468 4642 472
rect 4678 468 4682 472
rect 4702 468 4706 472
rect 4710 468 4714 472
rect 4742 468 4746 472
rect 4830 468 4834 472
rect 4870 468 4874 472
rect 4926 468 4930 472
rect 4958 468 4962 472
rect 5046 468 5050 472
rect 5078 468 5082 472
rect 1302 458 1306 462
rect 1310 458 1314 462
rect 1406 459 1410 463
rect 1526 458 1530 462
rect 1598 459 1602 463
rect 1630 458 1634 462
rect 1734 458 1738 462
rect 1790 458 1794 462
rect 1822 459 1826 463
rect 1854 458 1858 462
rect 1918 458 1922 462
rect 1934 458 1938 462
rect 1966 458 1970 462
rect 1982 458 1986 462
rect 1998 458 2002 462
rect 2054 458 2058 462
rect 2086 458 2090 462
rect 2102 458 2106 462
rect 2118 458 2122 462
rect 2142 458 2146 462
rect 2166 458 2170 462
rect 2246 459 2250 463
rect 2286 458 2290 462
rect 2294 458 2298 462
rect 2326 458 2330 462
rect 2358 458 2362 462
rect 2398 458 2402 462
rect 2414 458 2418 462
rect 2430 458 2434 462
rect 2534 458 2538 462
rect 2606 458 2610 462
rect 2638 459 2642 463
rect 2686 458 2690 462
rect 2718 458 2722 462
rect 2766 458 2770 462
rect 2782 458 2786 462
rect 2838 458 2842 462
rect 2870 458 2874 462
rect 2902 458 2906 462
rect 2910 458 2914 462
rect 2950 458 2954 462
rect 2990 458 2994 462
rect 3014 458 3018 462
rect 3022 458 3026 462
rect 3054 458 3058 462
rect 3102 458 3106 462
rect 3166 458 3170 462
rect 3206 458 3210 462
rect 3254 458 3258 462
rect 3270 458 3274 462
rect 3302 458 3306 462
rect 3326 458 3330 462
rect 3358 458 3362 462
rect 3422 458 3426 462
rect 3462 458 3466 462
rect 3486 458 3490 462
rect 3558 458 3562 462
rect 3598 458 3602 462
rect 3646 458 3650 462
rect 3662 458 3666 462
rect 3710 458 3714 462
rect 3758 458 3762 462
rect 3774 458 3778 462
rect 3822 458 3826 462
rect 3926 458 3930 462
rect 3934 458 3938 462
rect 3982 458 3986 462
rect 3990 458 3994 462
rect 4022 458 4026 462
rect 4038 458 4042 462
rect 4102 458 4106 462
rect 4166 458 4170 462
rect 4182 458 4186 462
rect 4198 458 4202 462
rect 4206 458 4210 462
rect 4270 458 4274 462
rect 4302 459 4306 463
rect 4350 458 4354 462
rect 4366 458 4370 462
rect 4382 458 4386 462
rect 4390 458 4394 462
rect 4414 458 4418 462
rect 4470 458 4474 462
rect 4502 458 4506 462
rect 4510 458 4514 462
rect 4574 458 4578 462
rect 4646 458 4650 462
rect 4670 458 4674 462
rect 4742 458 4746 462
rect 4750 458 4754 462
rect 4806 458 4810 462
rect 4838 459 4842 463
rect 5246 468 5250 472
rect 5278 468 5282 472
rect 4878 458 4882 462
rect 4918 458 4922 462
rect 4998 458 5002 462
rect 5054 458 5058 462
rect 5078 458 5082 462
rect 5086 458 5090 462
rect 5102 458 5106 462
rect 5110 458 5114 462
rect 5134 458 5138 462
rect 5198 458 5202 462
rect 5222 458 5226 462
rect 5286 458 5290 462
rect 1294 448 1298 452
rect 1670 448 1674 452
rect 1702 448 1706 452
rect 1950 448 1954 452
rect 2022 448 2026 452
rect 2070 448 2074 452
rect 2134 448 2138 452
rect 2310 448 2314 452
rect 2342 448 2346 452
rect 2414 448 2418 452
rect 2430 448 2434 452
rect 2454 448 2458 452
rect 2822 448 2826 452
rect 2838 448 2842 452
rect 2854 448 2858 452
rect 2870 448 2874 452
rect 3006 448 3010 452
rect 3190 448 3194 452
rect 3270 448 3274 452
rect 3286 448 3290 452
rect 3342 448 3346 452
rect 3358 448 3362 452
rect 3374 448 3378 452
rect 3558 448 3562 452
rect 3734 448 3738 452
rect 3878 448 3882 452
rect 3950 448 3954 452
rect 4206 448 4210 452
rect 4438 448 4442 452
rect 4486 448 4490 452
rect 4526 448 4530 452
rect 4686 448 4690 452
rect 4766 448 4770 452
rect 4790 448 4794 452
rect 4902 448 4906 452
rect 5070 448 5074 452
rect 5102 448 5106 452
rect 5158 448 5162 452
rect 654 438 658 442
rect 758 438 762 442
rect 1230 438 1234 442
rect 2446 438 2450 442
rect 2478 438 2482 442
rect 3254 438 3258 442
rect 3518 438 3522 442
rect 3582 438 3586 442
rect 3702 438 3706 442
rect 4654 438 4658 442
rect 3534 428 3538 432
rect 134 418 138 422
rect 478 418 482 422
rect 806 418 810 422
rect 2358 418 2362 422
rect 2926 418 2930 422
rect 3038 418 3042 422
rect 3302 418 3306 422
rect 3326 418 3330 422
rect 3390 418 3394 422
rect 3974 418 3978 422
rect 330 403 334 407
rect 337 403 341 407
rect 1354 403 1358 407
rect 1361 403 1365 407
rect 2386 403 2390 407
rect 2393 403 2397 407
rect 3402 403 3406 407
rect 3409 403 3413 407
rect 4426 403 4430 407
rect 4433 403 4437 407
rect 62 388 66 392
rect 182 388 186 392
rect 198 388 202 392
rect 550 388 554 392
rect 646 388 650 392
rect 742 388 746 392
rect 766 388 770 392
rect 934 388 938 392
rect 958 388 962 392
rect 1566 388 1570 392
rect 1766 388 1770 392
rect 1878 388 1882 392
rect 2206 388 2210 392
rect 2278 388 2282 392
rect 2590 388 2594 392
rect 2814 388 2818 392
rect 2990 388 2994 392
rect 3014 388 3018 392
rect 3062 388 3066 392
rect 3334 388 3338 392
rect 3534 388 3538 392
rect 3638 388 3642 392
rect 3670 388 3674 392
rect 3726 388 3730 392
rect 3790 388 3794 392
rect 3822 388 3826 392
rect 3926 388 3930 392
rect 4542 388 4546 392
rect 4662 388 4666 392
rect 4958 388 4962 392
rect 5142 388 5146 392
rect 5182 388 5186 392
rect 5238 388 5242 392
rect 5278 388 5282 392
rect 5294 388 5298 392
rect 750 378 754 382
rect 2710 378 2714 382
rect 3550 378 3554 382
rect 4038 378 4042 382
rect 1374 368 1378 372
rect 1478 368 1482 372
rect 1790 368 1794 372
rect 3094 368 3098 372
rect 4166 368 4170 372
rect 4350 368 4354 372
rect 206 358 210 362
rect 910 358 914 362
rect 126 348 130 352
rect 206 348 210 352
rect 254 348 258 352
rect 310 348 314 352
rect 326 348 330 352
rect 350 348 354 352
rect 398 348 402 352
rect 406 348 410 352
rect 454 348 458 352
rect 6 338 10 342
rect 70 338 74 342
rect 86 338 90 342
rect 190 338 194 342
rect 294 338 298 342
rect 358 338 362 342
rect 486 347 490 351
rect 582 347 586 351
rect 702 348 706 352
rect 710 348 714 352
rect 814 348 818 352
rect 838 348 842 352
rect 1270 358 1274 362
rect 942 348 946 352
rect 998 348 1002 352
rect 1006 348 1010 352
rect 1118 348 1122 352
rect 1198 348 1202 352
rect 1206 348 1210 352
rect 1230 348 1234 352
rect 1238 348 1242 352
rect 1254 348 1258 352
rect 1334 358 1338 362
rect 1350 358 1354 362
rect 1510 358 1514 362
rect 1590 358 1594 362
rect 1606 358 1610 362
rect 1638 358 1642 362
rect 1318 348 1322 352
rect 1334 348 1338 352
rect 1342 348 1346 352
rect 1414 347 1418 351
rect 1518 348 1522 352
rect 1534 348 1538 352
rect 1550 348 1554 352
rect 1582 348 1586 352
rect 1590 348 1594 352
rect 1622 348 1626 352
rect 1774 358 1778 362
rect 1822 358 1826 362
rect 1854 358 1858 362
rect 1934 358 1938 362
rect 2086 358 2090 362
rect 2246 358 2250 362
rect 2390 358 2394 362
rect 3054 358 3058 362
rect 3654 358 3658 362
rect 3710 358 3714 362
rect 3766 358 3770 362
rect 3806 358 3810 362
rect 3862 358 3866 362
rect 3878 358 3882 362
rect 1654 348 1658 352
rect 1662 348 1666 352
rect 1702 347 1706 351
rect 1798 348 1802 352
rect 1822 348 1826 352
rect 1830 348 1834 352
rect 1902 348 1906 352
rect 1918 348 1922 352
rect 1934 348 1938 352
rect 566 338 570 342
rect 662 338 666 342
rect 894 338 898 342
rect 942 338 946 342
rect 1014 338 1018 342
rect 1094 338 1098 342
rect 1198 338 1202 342
rect 1246 338 1250 342
rect 1302 338 1306 342
rect 1310 338 1314 342
rect 1342 338 1346 342
rect 1398 338 1402 342
rect 1422 338 1426 342
rect 1486 338 1490 342
rect 1542 338 1546 342
rect 1574 338 1578 342
rect 1582 338 1586 342
rect 1614 338 1618 342
rect 1670 338 1674 342
rect 1686 338 1690 342
rect 1718 338 1722 342
rect 1790 338 1794 342
rect 1798 338 1802 342
rect 1830 338 1834 342
rect 1878 338 1882 342
rect 1894 338 1898 342
rect 1910 338 1914 342
rect 1966 347 1970 351
rect 2038 348 2042 352
rect 2070 348 2074 352
rect 2110 348 2114 352
rect 2150 348 2154 352
rect 2174 348 2178 352
rect 2182 348 2186 352
rect 2214 348 2218 352
rect 2310 348 2314 352
rect 2342 347 2346 351
rect 2398 348 2402 352
rect 2406 348 2410 352
rect 2422 348 2426 352
rect 2430 348 2434 352
rect 2454 348 2458 352
rect 2462 348 2466 352
rect 2542 348 2546 352
rect 2614 348 2618 352
rect 2646 348 2650 352
rect 2670 348 2674 352
rect 2702 348 2706 352
rect 2758 348 2762 352
rect 2926 348 2930 352
rect 3006 348 3010 352
rect 3038 348 3042 352
rect 3054 348 3058 352
rect 3134 348 3138 352
rect 3174 348 3178 352
rect 3206 348 3210 352
rect 3214 348 3218 352
rect 3230 348 3234 352
rect 3294 348 3298 352
rect 3366 348 3370 352
rect 3390 348 3394 352
rect 3470 347 3474 351
rect 3550 348 3554 352
rect 3566 348 3570 352
rect 3606 348 3610 352
rect 3622 348 3626 352
rect 3646 348 3650 352
rect 3670 348 3674 352
rect 3694 348 3698 352
rect 3710 348 3714 352
rect 3726 348 3730 352
rect 3742 348 3746 352
rect 3758 348 3762 352
rect 3782 348 3786 352
rect 3830 348 3834 352
rect 3838 348 3842 352
rect 3894 348 3898 352
rect 3918 348 3922 352
rect 3982 348 3986 352
rect 1950 338 1954 342
rect 2062 338 2066 342
rect 2134 338 2138 342
rect 2190 338 2194 342
rect 2254 338 2258 342
rect 2270 338 2274 342
rect 2414 338 2418 342
rect 2462 338 2466 342
rect 2566 338 2570 342
rect 2598 338 2602 342
rect 2638 338 2642 342
rect 2678 338 2682 342
rect 2694 338 2698 342
rect 2766 338 2770 342
rect 2870 338 2874 342
rect 2902 338 2906 342
rect 3030 338 3034 342
rect 3158 338 3162 342
rect 3542 338 3546 342
rect 3574 338 3578 342
rect 3582 338 3586 342
rect 3678 338 3682 342
rect 3686 338 3690 342
rect 4102 347 4106 351
rect 4142 348 4146 352
rect 4150 348 4154 352
rect 4246 358 4250 362
rect 4526 358 4530 362
rect 4678 358 4682 362
rect 4974 358 4978 362
rect 5158 358 5162 362
rect 5166 358 5170 362
rect 5222 358 5226 362
rect 4182 348 4186 352
rect 4198 348 4202 352
rect 4206 348 4210 352
rect 4238 348 4242 352
rect 4286 347 4290 351
rect 4358 348 4362 352
rect 4390 348 4394 352
rect 4406 348 4410 352
rect 4454 347 4458 351
rect 4542 348 4546 352
rect 4606 348 4610 352
rect 4662 348 4666 352
rect 4686 348 4690 352
rect 4718 348 4722 352
rect 4750 348 4754 352
rect 4814 348 4818 352
rect 4878 348 4882 352
rect 4894 348 4898 352
rect 4910 348 4914 352
rect 4942 348 4946 352
rect 4982 348 4986 352
rect 5006 348 5010 352
rect 5014 348 5018 352
rect 5030 348 5034 352
rect 5078 348 5082 352
rect 5142 348 5146 352
rect 5182 348 5186 352
rect 5198 348 5202 352
rect 5238 348 5242 352
rect 5254 348 5258 352
rect 5286 348 5290 352
rect 3718 338 3722 342
rect 3750 338 3754 342
rect 3774 338 3778 342
rect 3974 338 3978 342
rect 4022 338 4026 342
rect 4134 338 4138 342
rect 4190 338 4194 342
rect 4230 338 4234 342
rect 4270 338 4274 342
rect 4294 338 4298 342
rect 4398 338 4402 342
rect 4462 338 4466 342
rect 310 328 314 332
rect 382 328 386 332
rect 438 328 442 332
rect 486 328 490 332
rect 758 328 762 332
rect 950 328 954 332
rect 1510 328 1514 332
rect 1518 328 1522 332
rect 1878 328 1882 332
rect 2038 328 2042 332
rect 2054 328 2058 332
rect 2094 328 2098 332
rect 2158 328 2162 332
rect 2206 328 2210 332
rect 2582 328 2586 332
rect 2654 328 2658 332
rect 2998 328 3002 332
rect 3022 328 3026 332
rect 3198 328 3202 332
rect 3302 328 3306 332
rect 3582 328 3586 332
rect 3598 328 3602 332
rect 3774 328 3778 332
rect 3814 328 3818 332
rect 3838 328 3842 332
rect 3854 328 3858 332
rect 4102 328 4106 332
rect 4254 328 4258 332
rect 4374 328 4378 332
rect 4566 338 4570 342
rect 4638 338 4642 342
rect 4654 338 4658 342
rect 4694 338 4698 342
rect 4886 338 4890 342
rect 4950 338 4954 342
rect 4990 338 4994 342
rect 5070 338 5074 342
rect 5118 338 5122 342
rect 5134 338 5138 342
rect 5190 338 5194 342
rect 5246 338 5250 342
rect 5262 338 5266 342
rect 4710 328 4714 332
rect 4806 328 4810 332
rect 4942 328 4946 332
rect 5214 328 5218 332
rect 5278 328 5282 332
rect 5302 328 5306 332
rect 366 318 370 322
rect 422 318 426 322
rect 646 318 650 322
rect 982 318 986 322
rect 1070 318 1074 322
rect 1278 318 1282 322
rect 2030 318 2034 322
rect 2086 318 2090 322
rect 2126 318 2130 322
rect 2230 318 2234 322
rect 2590 318 2594 322
rect 2630 318 2634 322
rect 2982 318 2986 322
rect 3902 318 3906 322
rect 4518 318 4522 322
rect 4702 318 4706 322
rect 4734 318 4738 322
rect 4766 318 4770 322
rect 4870 318 4874 322
rect 5206 318 5210 322
rect 850 303 854 307
rect 857 303 861 307
rect 1874 303 1878 307
rect 1881 303 1885 307
rect 2890 303 2894 307
rect 2897 303 2901 307
rect 3922 303 3926 307
rect 3929 303 3933 307
rect 4938 303 4942 307
rect 4945 303 4949 307
rect 38 288 42 292
rect 206 288 210 292
rect 398 288 402 292
rect 470 288 474 292
rect 742 288 746 292
rect 886 288 890 292
rect 982 288 986 292
rect 1270 288 1274 292
rect 1438 288 1442 292
rect 1534 288 1538 292
rect 1718 288 1722 292
rect 1798 288 1802 292
rect 1862 288 1866 292
rect 1974 288 1978 292
rect 2126 288 2130 292
rect 2142 288 2146 292
rect 2166 288 2170 292
rect 2246 288 2250 292
rect 2270 288 2274 292
rect 2318 288 2322 292
rect 2470 288 2474 292
rect 2582 288 2586 292
rect 2718 288 2722 292
rect 2854 288 2858 292
rect 3054 288 3058 292
rect 3438 288 3442 292
rect 3614 288 3618 292
rect 3646 288 3650 292
rect 3654 288 3658 292
rect 3718 288 3722 292
rect 3742 288 3746 292
rect 3910 288 3914 292
rect 4062 288 4066 292
rect 4350 288 4354 292
rect 4526 288 4530 292
rect 4606 288 4610 292
rect 4718 288 4722 292
rect 4750 288 4754 292
rect 4982 288 4986 292
rect 5014 288 5018 292
rect 5134 288 5138 292
rect 5158 288 5162 292
rect 5182 288 5186 292
rect 5206 288 5210 292
rect 5238 288 5242 292
rect 5278 288 5282 292
rect 22 278 26 282
rect 110 278 114 282
rect 238 278 242 282
rect 502 278 506 282
rect 566 278 570 282
rect 878 278 882 282
rect 1046 278 1050 282
rect 1126 278 1130 282
rect 1206 278 1210 282
rect 1294 278 1298 282
rect 70 268 74 272
rect 150 268 154 272
rect 222 268 226 272
rect 294 268 298 272
rect 318 268 322 272
rect 366 268 370 272
rect 454 268 458 272
rect 518 268 522 272
rect 662 268 666 272
rect 678 268 682 272
rect 766 268 770 272
rect 822 268 826 272
rect 1086 268 1090 272
rect 1102 268 1106 272
rect 1374 278 1378 282
rect 1590 278 1594 282
rect 1622 278 1626 282
rect 1726 278 1730 282
rect 1734 278 1738 282
rect 1774 278 1778 282
rect 1998 278 2002 282
rect 1318 268 1322 272
rect 1454 268 1458 272
rect 1542 268 1546 272
rect 1582 268 1586 272
rect 1638 268 1642 272
rect 1686 268 1690 272
rect 1742 268 1746 272
rect 1774 268 1778 272
rect 1790 268 1794 272
rect 1838 268 1842 272
rect 1926 268 1930 272
rect 1958 268 1962 272
rect 2158 278 2162 282
rect 2254 278 2258 282
rect 2278 278 2282 282
rect 2638 278 2642 282
rect 2646 278 2650 282
rect 2846 278 2850 282
rect 2886 278 2890 282
rect 2926 278 2930 282
rect 2958 278 2962 282
rect 3158 278 3162 282
rect 3486 278 3490 282
rect 3710 278 3714 282
rect 3726 278 3730 282
rect 3974 278 3978 282
rect 4022 278 4026 282
rect 2022 268 2026 272
rect 2190 268 2194 272
rect 2238 268 2242 272
rect 2302 268 2306 272
rect 2366 268 2370 272
rect 2430 268 2434 272
rect 2478 268 2482 272
rect 2518 268 2522 272
rect 2598 268 2602 272
rect 2678 268 2682 272
rect 2710 268 2714 272
rect 2782 268 2786 272
rect 2822 268 2826 272
rect 2838 268 2842 272
rect 2862 268 2866 272
rect 2918 268 2922 272
rect 2958 268 2962 272
rect 3062 268 3066 272
rect 3118 268 3122 272
rect 3206 268 3210 272
rect 3222 268 3226 272
rect 3254 268 3258 272
rect 3286 268 3290 272
rect 3342 268 3346 272
rect 3382 268 3386 272
rect 3518 268 3522 272
rect 3622 268 3626 272
rect 3670 268 3674 272
rect 3678 268 3682 272
rect 3710 268 3714 272
rect 3750 268 3754 272
rect 3790 268 3794 272
rect 3822 268 3826 272
rect 3830 268 3834 272
rect 3886 268 3890 272
rect 4358 278 4362 282
rect 4430 278 4434 282
rect 4534 278 4538 282
rect 4566 278 4570 282
rect 4630 278 4634 282
rect 4710 278 4714 282
rect 4758 278 4762 282
rect 4974 278 4978 282
rect 5006 278 5010 282
rect 5038 278 5042 282
rect 5070 278 5074 282
rect 5166 278 5170 282
rect 5174 278 5178 282
rect 5214 278 5218 282
rect 5270 278 5274 282
rect 5286 278 5290 282
rect 4046 268 4050 272
rect 4102 268 4106 272
rect 4126 268 4130 272
rect 4142 268 4146 272
rect 4182 268 4186 272
rect 4190 268 4194 272
rect 4206 268 4210 272
rect 4230 268 4234 272
rect 4366 268 4370 272
rect 4382 268 4386 272
rect 4398 268 4402 272
rect 4414 268 4418 272
rect 4518 268 4522 272
rect 4542 268 4546 272
rect 4646 268 4650 272
rect 4710 268 4714 272
rect 4734 268 4738 272
rect 4766 268 4770 272
rect 4782 268 4786 272
rect 4830 268 4834 272
rect 4838 268 4842 272
rect 4926 268 4930 272
rect 4990 268 4994 272
rect 5150 268 5154 272
rect 5198 268 5202 272
rect 5230 268 5234 272
rect 6 258 10 262
rect 54 258 58 262
rect 62 258 66 262
rect 94 258 98 262
rect 142 259 146 263
rect 214 258 218 262
rect 254 258 258 262
rect 278 258 282 262
rect 302 258 306 262
rect 342 258 346 262
rect 414 258 418 262
rect 438 258 442 262
rect 446 258 450 262
rect 454 258 458 262
rect 486 258 490 262
rect 558 258 562 262
rect 606 258 610 262
rect 614 258 618 262
rect 638 258 642 262
rect 686 258 690 262
rect 798 258 802 262
rect 806 258 810 262
rect 814 258 818 262
rect 862 258 866 262
rect 926 258 930 262
rect 950 259 954 263
rect 1038 258 1042 262
rect 1078 258 1082 262
rect 1110 258 1114 262
rect 1142 258 1146 262
rect 1166 258 1170 262
rect 1174 258 1178 262
rect 1214 258 1218 262
rect 1278 258 1282 262
rect 1310 258 1314 262
rect 1326 258 1330 262
rect 1374 259 1378 263
rect 1478 258 1482 262
rect 1566 258 1570 262
rect 1574 258 1578 262
rect 1606 258 1610 262
rect 1662 258 1666 262
rect 1750 258 1754 262
rect 1782 258 1786 262
rect 1854 258 1858 262
rect 1918 258 1922 262
rect 1982 258 1986 262
rect 2014 258 2018 262
rect 2030 258 2034 262
rect 2062 259 2066 263
rect 2094 258 2098 262
rect 2134 258 2138 262
rect 2174 258 2178 262
rect 2182 258 2186 262
rect 2214 258 2218 262
rect 2222 258 2226 262
rect 2230 258 2234 262
rect 2262 258 2266 262
rect 2286 258 2290 262
rect 2382 259 2386 263
rect 2430 258 2434 262
rect 2486 258 2490 262
rect 2526 258 2530 262
rect 2598 258 2602 262
rect 2622 258 2626 262
rect 2630 258 2634 262
rect 2670 258 2674 262
rect 2702 258 2706 262
rect 2774 258 2778 262
rect 2830 258 2834 262
rect 2910 258 2914 262
rect 2942 258 2946 262
rect 2990 259 2994 263
rect 3022 258 3026 262
rect 3070 258 3074 262
rect 3110 258 3114 262
rect 3182 258 3186 262
rect 3230 258 3234 262
rect 3262 258 3266 262
rect 3294 258 3298 262
rect 3334 258 3338 262
rect 3374 259 3378 263
rect 3462 258 3466 262
rect 3470 258 3474 262
rect 3494 258 3498 262
rect 3534 259 3538 263
rect 3622 258 3626 262
rect 3670 258 3674 262
rect 3726 258 3730 262
rect 3758 258 3762 262
rect 3798 258 3802 262
rect 3814 258 3818 262
rect 3838 258 3842 262
rect 3886 258 3890 262
rect 3966 258 3970 262
rect 4006 258 4010 262
rect 4038 258 4042 262
rect 4054 258 4058 262
rect 4102 258 4106 262
rect 4174 258 4178 262
rect 4198 258 4202 262
rect 4246 259 4250 263
rect 4278 258 4282 262
rect 4318 258 4322 262
rect 4334 258 4338 262
rect 4374 258 4378 262
rect 4406 258 4410 262
rect 4494 258 4498 262
rect 4502 258 4506 262
rect 4510 258 4514 262
rect 4558 258 4562 262
rect 4590 258 4594 262
rect 4678 259 4682 263
rect 4726 258 4730 262
rect 4734 258 4738 262
rect 4774 258 4778 262
rect 4790 258 4794 262
rect 4806 258 4810 262
rect 4910 258 4914 262
rect 4998 258 5002 262
rect 5022 258 5026 262
rect 5070 259 5074 263
rect 5142 258 5146 262
rect 5190 258 5194 262
rect 5222 258 5226 262
rect 5254 258 5258 262
rect 1814 248 1818 252
rect 2454 248 2458 252
rect 2646 248 2650 252
rect 2670 248 2674 252
rect 2686 248 2690 252
rect 2702 248 2706 252
rect 2814 248 2818 252
rect 3110 248 3114 252
rect 3246 248 3250 252
rect 3262 248 3266 252
rect 3310 248 3314 252
rect 3334 248 3338 252
rect 3646 248 3650 252
rect 3702 248 3706 252
rect 3766 248 3770 252
rect 3782 248 3786 252
rect 3798 248 3802 252
rect 3854 248 3858 252
rect 3878 248 3882 252
rect 4158 248 4162 252
rect 4174 248 4178 252
rect 4214 248 4218 252
rect 4390 248 4394 252
rect 4422 248 4426 252
rect 4558 248 4562 252
rect 4606 248 4610 252
rect 4790 248 4794 252
rect 902 238 906 242
rect 1518 238 1522 242
rect 1974 238 1978 242
rect 3086 238 3090 242
rect 3126 238 3130 242
rect 3278 238 3282 242
rect 3654 238 3658 242
rect 3926 238 3930 242
rect 86 218 90 222
rect 238 218 242 222
rect 270 218 274 222
rect 430 218 434 222
rect 598 218 602 222
rect 630 218 634 222
rect 854 218 858 222
rect 1150 218 1154 222
rect 3230 218 3234 222
rect 3814 218 3818 222
rect 4478 218 4482 222
rect 5030 218 5034 222
rect 330 203 334 207
rect 337 203 341 207
rect 1354 203 1358 207
rect 1361 203 1365 207
rect 2386 203 2390 207
rect 2393 203 2397 207
rect 3402 203 3406 207
rect 3409 203 3413 207
rect 4426 203 4430 207
rect 4433 203 4437 207
rect 166 188 170 192
rect 262 188 266 192
rect 390 188 394 192
rect 534 188 538 192
rect 566 188 570 192
rect 606 188 610 192
rect 718 188 722 192
rect 918 188 922 192
rect 1102 188 1106 192
rect 1214 188 1218 192
rect 1334 188 1338 192
rect 1534 188 1538 192
rect 2006 188 2010 192
rect 2246 188 2250 192
rect 2518 188 2522 192
rect 3222 188 3226 192
rect 3398 188 3402 192
rect 3542 188 3546 192
rect 3566 188 3570 192
rect 3654 188 3658 192
rect 3742 188 3746 192
rect 3854 188 3858 192
rect 4046 188 4050 192
rect 4206 188 4210 192
rect 4222 188 4226 192
rect 4382 188 4386 192
rect 4582 188 4586 192
rect 4966 188 4970 192
rect 5006 188 5010 192
rect 5078 188 5082 192
rect 5246 188 5250 192
rect 5278 188 5282 192
rect 2398 178 2402 182
rect 5230 178 5234 182
rect 150 168 154 172
rect 342 168 346 172
rect 1454 168 1458 172
rect 2750 168 2754 172
rect 3382 168 3386 172
rect 4366 168 4370 172
rect 4774 168 4778 172
rect 4790 168 4794 172
rect 734 158 738 162
rect 1518 158 1522 162
rect 3582 158 3586 162
rect 3678 158 3682 162
rect 3838 158 3842 162
rect 4054 158 4058 162
rect 102 147 106 151
rect 206 148 210 152
rect 294 147 298 151
rect 318 148 322 152
rect 398 148 402 152
rect 430 148 434 152
rect 518 148 522 152
rect 542 148 546 152
rect 574 148 578 152
rect 670 148 674 152
rect 718 148 722 152
rect 854 147 858 151
rect 886 148 890 152
rect 958 148 962 152
rect 1038 148 1042 152
rect 1046 148 1050 152
rect 1070 148 1074 152
rect 1078 148 1082 152
rect 1102 148 1106 152
rect 1150 148 1154 152
rect 1222 148 1226 152
rect 1254 148 1258 152
rect 1398 148 1402 152
rect 1462 148 1466 152
rect 1494 148 1498 152
rect 1534 148 1538 152
rect 1582 148 1586 152
rect 1662 148 1666 152
rect 1670 148 1674 152
rect 1694 148 1698 152
rect 1702 148 1706 152
rect 1774 147 1778 151
rect 1806 148 1810 152
rect 1822 148 1826 152
rect 1830 148 1834 152
rect 1846 148 1850 152
rect 1886 148 1890 152
rect 1942 147 1946 151
rect 1974 148 1978 152
rect 2014 148 2018 152
rect 2030 148 2034 152
rect 2038 148 2042 152
rect 2062 148 2066 152
rect 2094 148 2098 152
rect 2102 148 2106 152
rect 2126 148 2130 152
rect 2134 148 2138 152
rect 2190 148 2194 152
rect 2198 148 2202 152
rect 2254 148 2258 152
rect 2270 148 2274 152
rect 2278 148 2282 152
rect 2310 148 2314 152
rect 2334 148 2338 152
rect 2374 148 2378 152
rect 2566 148 2570 152
rect 2630 148 2634 152
rect 2646 148 2650 152
rect 2654 148 2658 152
rect 2678 148 2682 152
rect 2742 148 2746 152
rect 2782 148 2786 152
rect 2814 147 2818 151
rect 2846 148 2850 152
rect 2862 148 2866 152
rect 2894 148 2898 152
rect 2942 148 2946 152
rect 2982 148 2986 152
rect 3006 148 3010 152
rect 3046 148 3050 152
rect 3062 148 3066 152
rect 3070 148 3074 152
rect 3086 148 3090 152
rect 3094 148 3098 152
rect 3110 148 3114 152
rect 3134 148 3138 152
rect 3158 148 3162 152
rect 3302 148 3306 152
rect 3334 147 3338 151
rect 3422 148 3426 152
rect 3470 148 3474 152
rect 3478 148 3482 152
rect 3510 148 3514 152
rect 3550 148 3554 152
rect 3566 148 3570 152
rect 3606 148 3610 152
rect 3638 148 3642 152
rect 3654 148 3658 152
rect 3694 148 3698 152
rect 3702 148 3706 152
rect 3734 148 3738 152
rect 6 138 10 142
rect 86 138 90 142
rect 182 138 186 142
rect 230 138 234 142
rect 278 138 282 142
rect 406 138 410 142
rect 454 138 458 142
rect 550 138 554 142
rect 678 138 682 142
rect 710 138 714 142
rect 742 138 746 142
rect 1038 138 1042 142
rect 1118 138 1122 142
rect 1230 138 1234 142
rect 1278 138 1282 142
rect 1374 138 1378 142
rect 1470 138 1474 142
rect 1542 138 1546 142
rect 1662 138 1666 142
rect 1790 138 1794 142
rect 1894 138 1898 142
rect 1910 138 1914 142
rect 1926 138 1930 142
rect 2078 138 2082 142
rect 2094 138 2098 142
rect 2358 138 2362 142
rect 2462 138 2466 142
rect 2526 138 2530 142
rect 2542 138 2546 142
rect 2702 138 2706 142
rect 2830 138 2834 142
rect 2854 138 2858 142
rect 2934 138 2938 142
rect 3118 138 3122 142
rect 3166 138 3170 142
rect 3238 138 3242 142
rect 3318 138 3322 142
rect 3430 138 3434 142
rect 3486 138 3490 142
rect 3806 147 3810 151
rect 3854 148 3858 152
rect 3870 148 3874 152
rect 3918 148 3922 152
rect 3974 148 3978 152
rect 3998 148 4002 152
rect 4078 148 4082 152
rect 4102 148 4106 152
rect 4110 148 4114 152
rect 4150 148 4154 152
rect 4302 148 4306 152
rect 4414 148 4418 152
rect 4446 147 4450 151
rect 4518 147 4522 151
rect 4550 148 4554 152
rect 4590 148 4594 152
rect 4638 148 4642 152
rect 4710 148 4714 152
rect 4734 148 4738 152
rect 4750 148 4754 152
rect 4766 148 4770 152
rect 4814 148 4818 152
rect 4894 147 4898 151
rect 4926 148 4930 152
rect 4990 148 4994 152
rect 5014 148 5018 152
rect 5022 148 5026 152
rect 5030 148 5034 152
rect 5038 148 5042 152
rect 5062 148 5066 152
rect 5118 148 5122 152
rect 5134 148 5138 152
rect 5246 148 5250 152
rect 5270 148 5274 152
rect 3630 138 3634 142
rect 3646 138 3650 142
rect 3678 138 3682 142
rect 3822 138 3826 142
rect 3862 138 3866 142
rect 3870 138 3874 142
rect 4070 138 4074 142
rect 4126 138 4130 142
rect 4278 138 4282 142
rect 4310 138 4314 142
rect 4462 138 4466 142
rect 4486 138 4490 142
rect 4598 138 4602 142
rect 4646 138 4650 142
rect 4758 138 4762 142
rect 5070 138 5074 142
rect 5158 138 5162 142
rect 5174 138 5178 142
rect 446 128 450 132
rect 526 128 530 132
rect 590 128 594 132
rect 598 128 602 132
rect 950 128 954 132
rect 1086 128 1090 132
rect 1270 128 1274 132
rect 1478 128 1482 132
rect 1510 128 1514 132
rect 1574 128 1578 132
rect 1806 128 1810 132
rect 1910 128 1914 132
rect 1942 128 1946 132
rect 1974 128 1978 132
rect 2014 128 2018 132
rect 2254 128 2258 132
rect 2318 128 2322 132
rect 2662 128 2666 132
rect 2726 128 2730 132
rect 2878 128 2882 132
rect 2918 128 2922 132
rect 3142 128 3146 132
rect 3454 128 3458 132
rect 3526 128 3530 132
rect 3534 128 3538 132
rect 3590 128 3594 132
rect 3622 128 3626 132
rect 3678 128 3682 132
rect 3902 128 3906 132
rect 3966 128 3970 132
rect 4038 128 4042 132
rect 4054 128 4058 132
rect 4174 128 4178 132
rect 4286 128 4290 132
rect 4622 128 4626 132
rect 4718 128 4722 132
rect 5262 128 5266 132
rect 5286 128 5290 132
rect 62 118 66 122
rect 414 118 418 122
rect 614 118 618 122
rect 798 118 802 122
rect 1238 118 1242 122
rect 1710 118 1714 122
rect 2054 118 2058 122
rect 2286 118 2290 122
rect 2350 118 2354 122
rect 2710 118 2714 122
rect 2926 118 2930 122
rect 3438 118 3442 122
rect 3494 118 3498 122
rect 3710 118 3714 122
rect 3886 118 3890 122
rect 4030 118 4034 122
rect 4046 118 4050 122
rect 4294 118 4298 122
rect 4606 118 4610 122
rect 4958 118 4962 122
rect 850 103 854 107
rect 857 103 861 107
rect 1874 103 1878 107
rect 1881 103 1885 107
rect 2890 103 2894 107
rect 2897 103 2901 107
rect 3922 103 3926 107
rect 3929 103 3933 107
rect 4938 103 4942 107
rect 4945 103 4949 107
rect 6 88 10 92
rect 310 88 314 92
rect 422 88 426 92
rect 518 88 522 92
rect 702 88 706 92
rect 718 88 722 92
rect 830 88 834 92
rect 1006 88 1010 92
rect 1318 88 1322 92
rect 1342 88 1346 92
rect 1622 88 1626 92
rect 1646 88 1650 92
rect 1686 88 1690 92
rect 1870 88 1874 92
rect 1902 88 1906 92
rect 2006 88 2010 92
rect 2102 88 2106 92
rect 2366 88 2370 92
rect 2782 88 2786 92
rect 2878 88 2882 92
rect 2894 88 2898 92
rect 3014 88 3018 92
rect 3110 88 3114 92
rect 3118 88 3122 92
rect 3358 88 3362 92
rect 3470 88 3474 92
rect 3478 88 3482 92
rect 3718 88 3722 92
rect 3870 88 3874 92
rect 3894 88 3898 92
rect 3950 88 3954 92
rect 4062 88 4066 92
rect 4110 88 4114 92
rect 4238 88 4242 92
rect 4254 88 4258 92
rect 4366 88 4370 92
rect 4406 88 4410 92
rect 4654 88 4658 92
rect 4766 88 4770 92
rect 4806 88 4810 92
rect 4814 88 4818 92
rect 4830 88 4834 92
rect 4942 88 4946 92
rect 5094 88 5098 92
rect 102 78 106 82
rect 214 78 218 82
rect 454 78 458 82
rect 550 78 554 82
rect 654 78 658 82
rect 710 78 714 82
rect 838 78 842 82
rect 846 78 850 82
rect 1030 78 1034 82
rect 1062 78 1066 82
rect 1198 78 1202 82
rect 1254 78 1258 82
rect 1350 78 1354 82
rect 1422 78 1426 82
rect 62 68 66 72
rect 86 68 90 72
rect 126 68 130 72
rect 174 68 178 72
rect 190 68 194 72
rect 230 68 234 72
rect 278 68 282 72
rect 342 68 346 72
rect 694 68 698 72
rect 798 68 802 72
rect 822 68 826 72
rect 902 68 906 72
rect 926 68 930 72
rect 950 68 954 72
rect 1022 68 1026 72
rect 1078 68 1082 72
rect 1334 68 1338 72
rect 1486 68 1490 72
rect 1574 68 1578 72
rect 1638 68 1642 72
rect 1662 78 1666 82
rect 1910 78 1914 82
rect 1942 78 1946 82
rect 2190 78 2194 82
rect 2478 78 2482 82
rect 2510 78 2514 82
rect 2614 78 2618 82
rect 2910 78 2914 82
rect 3230 78 3234 82
rect 1790 68 1794 72
rect 2046 68 2050 72
rect 2374 68 2378 72
rect 2550 68 2554 72
rect 2566 68 2570 72
rect 2734 68 2738 72
rect 2830 68 2834 72
rect 2958 68 2962 72
rect 3030 68 3034 72
rect 3198 68 3202 72
rect 3622 78 3626 82
rect 3774 78 3778 82
rect 3942 78 3946 82
rect 4142 78 4146 82
rect 4246 78 4250 82
rect 4390 78 4394 82
rect 3254 68 3258 72
rect 3310 68 3314 72
rect 3422 68 3426 72
rect 3558 68 3562 72
rect 3582 68 3586 72
rect 3734 68 3738 72
rect 3886 68 3890 72
rect 4030 68 4034 72
rect 4094 68 4098 72
rect 4262 68 4266 72
rect 4286 68 4290 72
rect 4542 78 4546 82
rect 4798 78 4802 82
rect 4822 78 4826 82
rect 4414 68 4418 72
rect 4478 68 4482 72
rect 4590 68 4594 72
rect 4646 68 4650 72
rect 4750 68 4754 72
rect 4790 68 4794 72
rect 4910 68 4914 72
rect 5022 68 5026 72
rect 5038 68 5042 72
rect 5110 68 5114 72
rect 5214 68 5218 72
rect 5278 68 5282 72
rect 70 59 74 63
rect 118 58 122 62
rect 126 58 130 62
rect 150 58 154 62
rect 158 58 162 62
rect 166 58 170 62
rect 198 58 202 62
rect 246 59 250 63
rect 366 58 370 62
rect 462 58 466 62
rect 558 58 562 62
rect 638 58 642 62
rect 646 58 650 62
rect 670 58 674 62
rect 686 58 690 62
rect 782 59 786 63
rect 814 58 818 62
rect 878 58 882 62
rect 910 58 914 62
rect 966 58 970 62
rect 1014 58 1018 62
rect 1046 58 1050 62
rect 1110 58 1114 62
rect 1166 58 1170 62
rect 1182 58 1186 62
rect 1190 58 1194 62
rect 1214 58 1218 62
rect 1254 59 1258 63
rect 1326 58 1330 62
rect 1358 58 1362 62
rect 1382 58 1386 62
rect 1406 58 1410 62
rect 1494 58 1498 62
rect 1566 58 1570 62
rect 1630 58 1634 62
rect 1678 58 1682 62
rect 1750 59 1754 63
rect 1814 58 1818 62
rect 1894 58 1898 62
rect 1950 58 1954 62
rect 2062 58 2066 62
rect 2118 58 2122 62
rect 2142 58 2146 62
rect 2150 58 2154 62
rect 2166 58 2170 62
rect 2230 58 2234 62
rect 2302 58 2306 62
rect 2326 58 2330 62
rect 2414 58 2418 62
rect 2438 58 2442 62
rect 2478 58 2482 62
rect 2494 58 2498 62
rect 2502 58 2506 62
rect 2542 58 2546 62
rect 2574 58 2578 62
rect 2654 58 2658 62
rect 2726 58 2730 62
rect 2822 58 2826 62
rect 2886 58 2890 62
rect 2958 58 2962 62
rect 3054 58 3058 62
rect 3182 59 3186 63
rect 3214 58 3218 62
rect 3230 58 3234 62
rect 3262 58 3266 62
rect 3302 58 3306 62
rect 3414 58 3418 62
rect 3542 59 3546 63
rect 3574 58 3578 62
rect 3606 58 3610 62
rect 3622 58 3626 62
rect 3654 59 3658 63
rect 3686 58 3690 62
rect 3726 58 3730 62
rect 3758 58 3762 62
rect 3806 59 3810 63
rect 3838 58 3842 62
rect 3878 58 3882 62
rect 3910 58 3914 62
rect 4014 59 4018 63
rect 4046 58 4050 62
rect 4078 58 4082 62
rect 4086 58 4090 62
rect 4094 58 4098 62
rect 4126 58 4130 62
rect 4182 58 4186 62
rect 4206 58 4210 62
rect 4270 58 4274 62
rect 4326 58 4330 62
rect 4334 58 4338 62
rect 4374 58 4378 62
rect 4422 58 4426 62
rect 4446 58 4450 62
rect 4454 58 4458 62
rect 4550 58 4554 62
rect 4606 58 4610 62
rect 4614 58 4618 62
rect 4718 58 4722 62
rect 4782 58 4786 62
rect 4894 59 4898 63
rect 5006 59 5010 63
rect 5182 58 5186 62
rect 5230 59 5234 63
rect 622 48 626 52
rect 886 48 890 52
rect 1398 48 1402 52
rect 2126 48 2130 52
rect 3598 48 3602 52
rect 3750 48 3754 52
rect 4766 48 4770 52
rect 5166 48 5170 52
rect 5198 38 5202 42
rect 330 3 334 7
rect 337 3 341 7
rect 1354 3 1358 7
rect 1361 3 1365 7
rect 2386 3 2390 7
rect 2393 3 2397 7
rect 3402 3 3406 7
rect 3409 3 3413 7
rect 4426 3 4430 7
rect 4433 3 4437 7
<< metal2 >>
rect 310 5128 314 5132
rect 526 5131 530 5132
rect 958 5131 962 5132
rect 518 5128 530 5131
rect 950 5128 962 5131
rect 1094 5128 1098 5132
rect 1190 5131 1194 5132
rect 1430 5131 1434 5132
rect 1454 5131 1458 5132
rect 1550 5131 1554 5132
rect 1190 5128 1201 5131
rect 1430 5128 1441 5131
rect 1454 5128 1465 5131
rect 310 5102 313 5128
rect 518 5092 521 5128
rect 848 5103 850 5107
rect 854 5103 857 5107
rect 861 5103 864 5107
rect 950 5092 953 5128
rect 650 5088 654 5091
rect 810 5088 814 5091
rect 290 5078 294 5081
rect 306 5078 310 5081
rect 322 5078 326 5081
rect 386 5078 390 5081
rect 10 4988 14 4991
rect 38 4952 41 5068
rect 50 5058 54 5061
rect 102 4962 105 5038
rect 38 4862 41 4948
rect 70 4942 73 4947
rect 102 4932 105 4958
rect 110 4952 113 5078
rect 150 5072 153 5078
rect 174 5072 177 5078
rect 510 5072 513 5088
rect 702 5082 705 5088
rect 322 5068 326 5071
rect 118 5062 121 5068
rect 190 5062 193 5068
rect 146 5058 150 5061
rect 170 5058 174 5061
rect 210 5059 214 5062
rect 158 5052 161 5058
rect 122 5048 126 5051
rect 158 4992 161 5048
rect 222 4992 225 5018
rect 278 4972 281 4978
rect 294 4971 297 5048
rect 328 5003 330 5007
rect 334 5003 337 5007
rect 341 5003 344 5007
rect 290 4968 297 4971
rect 138 4948 142 4951
rect 118 4942 121 4948
rect 126 4912 129 4938
rect 134 4922 137 4928
rect 70 4863 73 4898
rect 106 4878 110 4881
rect 118 4872 121 4878
rect 126 4872 129 4908
rect 150 4862 153 4958
rect 158 4952 161 4958
rect 166 4922 169 4968
rect 186 4948 190 4951
rect 210 4948 214 4951
rect 222 4942 225 4968
rect 286 4962 289 4968
rect 258 4958 262 4961
rect 350 4961 353 5058
rect 374 5002 377 5058
rect 382 5052 385 5068
rect 342 4958 353 4961
rect 390 4962 393 5018
rect 406 5012 409 5068
rect 446 5062 449 5068
rect 466 5058 470 5061
rect 438 5042 441 5058
rect 454 5042 457 5048
rect 242 4948 246 4951
rect 270 4942 273 4958
rect 278 4952 281 4958
rect 242 4938 246 4941
rect 166 4882 169 4888
rect 182 4872 185 4928
rect 190 4922 193 4938
rect 210 4928 214 4931
rect 190 4892 193 4898
rect 38 4852 41 4858
rect 102 4832 105 4858
rect 134 4852 137 4858
rect 150 4852 153 4858
rect 174 4852 177 4858
rect 162 4848 166 4851
rect 6 4742 9 4818
rect 62 4742 65 4768
rect 82 4758 86 4761
rect 102 4752 105 4818
rect 110 4792 113 4818
rect 118 4752 121 4828
rect 126 4762 129 4768
rect 82 4738 86 4741
rect 6 4732 9 4738
rect 34 4718 38 4721
rect 54 4712 57 4738
rect 62 4722 65 4738
rect 86 4722 89 4728
rect 38 4672 41 4698
rect 14 4562 17 4568
rect 22 4532 25 4538
rect 22 4492 25 4528
rect 30 4512 33 4538
rect 38 4531 41 4668
rect 46 4662 49 4668
rect 94 4662 97 4688
rect 102 4662 105 4668
rect 94 4648 102 4651
rect 94 4592 97 4648
rect 110 4602 113 4718
rect 126 4681 129 4748
rect 134 4692 137 4818
rect 150 4792 153 4838
rect 142 4762 145 4768
rect 162 4748 166 4751
rect 142 4722 145 4748
rect 154 4738 158 4741
rect 158 4682 161 4728
rect 126 4678 134 4681
rect 122 4668 126 4671
rect 150 4632 153 4658
rect 158 4622 161 4678
rect 182 4642 185 4868
rect 198 4861 201 4918
rect 198 4858 206 4861
rect 214 4822 217 4848
rect 190 4762 193 4768
rect 206 4762 209 4778
rect 222 4772 225 4938
rect 230 4862 233 4928
rect 246 4872 249 4898
rect 254 4872 257 4928
rect 294 4862 297 4958
rect 326 4952 329 4958
rect 310 4942 313 4948
rect 302 4882 305 4938
rect 310 4892 313 4938
rect 342 4932 345 4958
rect 370 4948 374 4951
rect 414 4951 417 5018
rect 454 4982 457 5038
rect 462 5032 465 5048
rect 470 5022 473 5038
rect 486 5022 489 5048
rect 494 5032 497 5058
rect 502 5052 505 5058
rect 534 5012 537 5058
rect 542 5052 545 5078
rect 558 5072 561 5078
rect 562 5058 566 5061
rect 582 5042 585 5058
rect 590 5042 593 5058
rect 598 5042 601 5048
rect 606 5032 609 5048
rect 622 5042 625 5068
rect 482 4968 486 4971
rect 426 4958 430 4961
rect 458 4958 462 4961
rect 470 4952 473 4958
rect 494 4952 497 4998
rect 502 4992 505 5008
rect 534 4992 537 5008
rect 378 4948 385 4951
rect 414 4948 422 4951
rect 350 4942 353 4948
rect 362 4938 366 4941
rect 382 4932 385 4948
rect 446 4942 449 4948
rect 394 4938 398 4941
rect 458 4938 462 4941
rect 414 4932 417 4938
rect 342 4882 345 4928
rect 358 4922 361 4928
rect 470 4922 473 4928
rect 310 4862 313 4868
rect 310 4852 313 4858
rect 318 4852 321 4858
rect 254 4842 257 4848
rect 230 4762 233 4768
rect 194 4748 198 4751
rect 230 4742 233 4748
rect 262 4742 265 4747
rect 90 4568 94 4571
rect 110 4562 113 4588
rect 182 4582 185 4618
rect 190 4592 193 4738
rect 214 4732 217 4738
rect 206 4682 209 4718
rect 222 4692 225 4708
rect 238 4692 241 4718
rect 246 4702 249 4738
rect 210 4668 214 4671
rect 198 4662 201 4668
rect 214 4652 217 4658
rect 258 4648 262 4651
rect 230 4642 233 4648
rect 214 4638 222 4641
rect 130 4568 134 4571
rect 154 4568 158 4571
rect 178 4568 182 4571
rect 198 4562 201 4638
rect 214 4592 217 4638
rect 226 4568 230 4571
rect 250 4568 254 4571
rect 262 4562 265 4578
rect 50 4558 54 4561
rect 98 4558 102 4561
rect 54 4552 57 4558
rect 70 4542 73 4558
rect 50 4538 54 4541
rect 38 4528 49 4531
rect 30 4472 33 4508
rect 6 4452 9 4468
rect 6 4362 9 4438
rect 22 4372 25 4448
rect 38 4392 41 4458
rect 6 4302 9 4358
rect 22 4352 25 4368
rect 22 4292 25 4338
rect 30 4332 33 4338
rect 10 4288 14 4291
rect 46 4272 49 4528
rect 62 4482 65 4518
rect 54 4452 57 4478
rect 62 4462 65 4468
rect 78 4462 81 4518
rect 86 4452 89 4548
rect 94 4492 97 4548
rect 110 4512 113 4558
rect 166 4552 169 4558
rect 270 4552 273 4848
rect 342 4842 345 4858
rect 282 4838 286 4841
rect 330 4838 334 4841
rect 278 4782 281 4818
rect 318 4772 321 4818
rect 328 4803 330 4807
rect 334 4803 337 4807
rect 341 4803 344 4807
rect 330 4788 334 4791
rect 318 4672 321 4698
rect 290 4668 294 4671
rect 278 4652 281 4658
rect 334 4652 337 4659
rect 342 4622 345 4738
rect 350 4632 353 4918
rect 390 4882 393 4898
rect 406 4882 409 4918
rect 430 4912 433 4918
rect 430 4882 433 4908
rect 374 4862 377 4878
rect 390 4872 393 4878
rect 454 4872 457 4878
rect 358 4852 361 4858
rect 422 4852 425 4868
rect 462 4862 465 4898
rect 502 4892 505 4978
rect 534 4972 537 4978
rect 518 4952 521 4958
rect 534 4932 537 4948
rect 542 4942 545 5018
rect 574 4961 577 5018
rect 566 4958 577 4961
rect 614 5002 617 5018
rect 566 4942 569 4958
rect 602 4948 606 4951
rect 574 4942 577 4948
rect 614 4942 617 4998
rect 622 4962 625 4968
rect 630 4951 633 5078
rect 694 5072 697 5078
rect 750 5072 753 5088
rect 818 5078 822 5081
rect 798 5072 801 5078
rect 910 5072 913 5078
rect 650 5068 654 5071
rect 714 5068 718 5071
rect 850 5068 854 5071
rect 658 5058 662 5061
rect 662 4992 665 5028
rect 626 4948 633 4951
rect 554 4938 558 4941
rect 606 4932 609 4938
rect 514 4928 518 4931
rect 546 4928 550 4931
rect 534 4892 537 4928
rect 566 4892 569 4908
rect 582 4902 585 4918
rect 630 4892 633 4948
rect 638 4942 641 4958
rect 694 4952 697 5068
rect 726 5062 729 5068
rect 726 5021 729 5058
rect 742 5052 745 5068
rect 778 5058 782 5061
rect 734 5032 737 5038
rect 726 5018 737 5021
rect 734 4992 737 5018
rect 742 4972 745 5028
rect 738 4968 742 4971
rect 646 4922 649 4938
rect 694 4921 697 4938
rect 686 4918 697 4921
rect 578 4878 582 4881
rect 642 4878 646 4881
rect 542 4872 545 4878
rect 498 4868 505 4871
rect 410 4848 414 4851
rect 318 4592 321 4618
rect 328 4603 330 4607
rect 334 4603 337 4607
rect 341 4603 344 4607
rect 302 4568 310 4571
rect 294 4562 297 4568
rect 302 4551 305 4568
rect 322 4558 326 4561
rect 350 4552 353 4628
rect 358 4582 361 4848
rect 366 4762 369 4818
rect 374 4792 377 4848
rect 398 4842 401 4848
rect 430 4841 433 4858
rect 478 4852 481 4868
rect 486 4852 489 4858
rect 502 4852 505 4868
rect 510 4862 513 4868
rect 522 4858 526 4861
rect 422 4838 433 4841
rect 442 4838 446 4841
rect 386 4768 390 4771
rect 398 4762 401 4798
rect 422 4792 425 4838
rect 434 4818 438 4821
rect 462 4782 465 4818
rect 486 4782 489 4848
rect 502 4792 505 4848
rect 518 4792 521 4838
rect 526 4812 529 4848
rect 550 4782 553 4858
rect 558 4822 561 4868
rect 574 4842 577 4868
rect 622 4862 625 4868
rect 638 4862 641 4868
rect 582 4792 585 4858
rect 606 4852 609 4858
rect 642 4848 646 4851
rect 606 4802 609 4848
rect 430 4778 438 4781
rect 418 4768 422 4771
rect 430 4762 433 4778
rect 426 4748 430 4751
rect 390 4742 393 4748
rect 438 4722 441 4738
rect 366 4692 369 4718
rect 438 4692 441 4718
rect 366 4672 369 4678
rect 422 4662 425 4678
rect 406 4652 409 4658
rect 402 4638 406 4641
rect 394 4618 398 4621
rect 446 4602 449 4718
rect 462 4712 465 4748
rect 470 4742 473 4758
rect 486 4742 489 4748
rect 518 4742 521 4748
rect 506 4738 510 4741
rect 494 4702 497 4738
rect 534 4692 537 4758
rect 502 4672 505 4678
rect 486 4662 489 4668
rect 526 4662 529 4688
rect 542 4662 545 4748
rect 550 4742 553 4758
rect 566 4742 569 4778
rect 582 4772 585 4788
rect 590 4752 593 4798
rect 606 4752 609 4778
rect 614 4762 617 4818
rect 654 4792 657 4828
rect 662 4792 665 4858
rect 670 4822 673 4918
rect 678 4862 681 4878
rect 622 4782 625 4788
rect 646 4782 649 4788
rect 662 4762 665 4768
rect 598 4742 601 4748
rect 570 4738 574 4741
rect 558 4732 561 4738
rect 590 4732 593 4738
rect 626 4728 630 4731
rect 638 4712 641 4738
rect 594 4688 598 4691
rect 606 4682 609 4698
rect 606 4672 609 4678
rect 638 4672 641 4708
rect 474 4648 478 4651
rect 594 4648 598 4651
rect 582 4612 585 4618
rect 470 4562 473 4568
rect 446 4552 449 4558
rect 298 4548 305 4551
rect 422 4548 441 4551
rect 126 4532 129 4548
rect 142 4522 145 4538
rect 158 4492 161 4538
rect 142 4482 145 4488
rect 166 4472 169 4478
rect 182 4472 185 4478
rect 98 4458 102 4461
rect 118 4452 121 4458
rect 78 4392 81 4418
rect 102 4372 105 4438
rect 110 4392 113 4428
rect 126 4412 129 4468
rect 170 4458 174 4461
rect 190 4422 193 4548
rect 206 4482 209 4528
rect 214 4512 217 4548
rect 234 4538 238 4541
rect 230 4522 233 4538
rect 246 4532 249 4548
rect 214 4482 217 4488
rect 190 4392 193 4408
rect 214 4392 217 4468
rect 226 4458 230 4461
rect 246 4392 249 4508
rect 270 4472 273 4538
rect 278 4532 281 4548
rect 310 4492 313 4548
rect 374 4542 377 4548
rect 406 4542 409 4548
rect 370 4528 377 4531
rect 358 4482 361 4518
rect 290 4468 294 4471
rect 262 4452 265 4468
rect 330 4458 334 4461
rect 78 4362 81 4368
rect 142 4362 145 4388
rect 94 4342 97 4348
rect 102 4342 105 4358
rect 118 4302 121 4358
rect 126 4342 129 4358
rect 134 4302 137 4340
rect 142 4282 145 4358
rect 174 4352 177 4378
rect 198 4362 201 4378
rect 202 4348 206 4351
rect 158 4342 161 4348
rect 154 4328 158 4331
rect 102 4272 105 4278
rect 62 4262 65 4268
rect 14 4192 17 4248
rect 86 4241 89 4268
rect 102 4252 105 4258
rect 118 4252 121 4258
rect 86 4238 97 4241
rect 22 4162 25 4168
rect 78 4142 81 4198
rect 6 4092 9 4138
rect 62 4062 65 4118
rect 86 4112 89 4158
rect 94 4142 97 4238
rect 102 4192 105 4238
rect 142 4202 145 4278
rect 150 4272 153 4328
rect 166 4292 169 4298
rect 174 4278 177 4348
rect 214 4342 217 4378
rect 214 4312 217 4338
rect 230 4332 233 4388
rect 250 4368 254 4371
rect 270 4362 273 4448
rect 278 4432 281 4458
rect 310 4452 313 4458
rect 278 4392 281 4418
rect 302 4372 305 4438
rect 318 4381 321 4448
rect 342 4432 345 4478
rect 358 4462 361 4468
rect 366 4462 369 4498
rect 374 4462 377 4528
rect 382 4492 385 4538
rect 422 4532 425 4548
rect 438 4542 441 4548
rect 510 4542 513 4558
rect 526 4552 529 4598
rect 466 4538 470 4541
rect 506 4538 510 4541
rect 430 4532 433 4538
rect 402 4528 406 4531
rect 442 4528 446 4531
rect 462 4522 465 4528
rect 390 4502 393 4518
rect 328 4403 330 4407
rect 334 4403 337 4407
rect 341 4403 344 4407
rect 366 4382 369 4458
rect 374 4422 377 4458
rect 318 4378 329 4381
rect 282 4368 286 4371
rect 318 4362 321 4368
rect 210 4278 214 4281
rect 222 4272 225 4278
rect 150 4242 153 4268
rect 226 4258 230 4261
rect 214 4192 217 4218
rect 222 4192 225 4248
rect 238 4241 241 4358
rect 270 4352 273 4358
rect 250 4348 254 4351
rect 278 4292 281 4348
rect 302 4342 305 4348
rect 310 4272 313 4278
rect 250 4268 254 4271
rect 246 4252 249 4258
rect 302 4252 305 4268
rect 318 4252 321 4258
rect 238 4238 249 4241
rect 110 4142 113 4148
rect 134 4142 137 4148
rect 70 4062 73 4108
rect 94 4101 97 4138
rect 118 4132 121 4138
rect 142 4132 145 4178
rect 154 4168 158 4171
rect 174 4152 177 4178
rect 230 4172 233 4228
rect 214 4152 217 4158
rect 222 4152 225 4168
rect 162 4148 166 4151
rect 166 4142 169 4148
rect 134 4112 137 4118
rect 86 4098 97 4101
rect 86 4072 89 4098
rect 134 4092 137 4098
rect 166 4092 169 4118
rect 182 4072 185 4138
rect 202 4128 206 4131
rect 202 4088 206 4091
rect 202 4078 206 4081
rect 230 4072 233 4078
rect 154 4068 158 4071
rect 6 3962 9 3968
rect 22 3952 25 3988
rect 38 3952 41 3958
rect 6 3922 9 3928
rect 14 3792 17 3868
rect 38 3842 41 3948
rect 46 3892 49 4028
rect 62 3992 65 4008
rect 62 3942 65 3948
rect 70 3942 73 4058
rect 86 4002 89 4068
rect 102 4052 105 4068
rect 198 4062 201 4068
rect 210 4058 217 4061
rect 154 4048 158 4051
rect 86 3952 89 3978
rect 74 3938 78 3941
rect 54 3932 57 3938
rect 62 3922 65 3928
rect 54 3882 57 3898
rect 62 3872 65 3908
rect 86 3872 89 3938
rect 94 3892 97 4038
rect 102 3992 105 4038
rect 126 3952 129 3958
rect 134 3951 137 3998
rect 174 3982 177 3998
rect 146 3958 150 3961
rect 134 3948 145 3951
rect 6 3672 9 3738
rect 14 3682 17 3748
rect 22 3692 25 3838
rect 46 3792 49 3858
rect 70 3832 73 3868
rect 78 3842 81 3858
rect 110 3852 113 3928
rect 126 3872 129 3878
rect 122 3858 126 3861
rect 102 3832 105 3848
rect 110 3831 113 3848
rect 134 3842 137 3848
rect 122 3838 126 3841
rect 106 3828 113 3831
rect 30 3762 33 3778
rect 58 3768 62 3771
rect 38 3762 41 3768
rect 30 3682 33 3758
rect 50 3748 54 3751
rect 14 3672 17 3678
rect 38 3672 41 3698
rect 62 3682 65 3698
rect 70 3692 73 3808
rect 78 3772 81 3778
rect 90 3768 97 3771
rect 106 3768 110 3771
rect 82 3758 86 3761
rect 82 3748 86 3751
rect 94 3692 97 3768
rect 106 3748 110 3751
rect 106 3738 110 3741
rect 6 3662 9 3668
rect 14 3652 17 3668
rect 38 3662 41 3668
rect 58 3658 62 3661
rect 78 3652 81 3658
rect 86 3652 89 3658
rect 10 3518 14 3521
rect 54 3472 57 3648
rect 102 3582 105 3668
rect 110 3652 113 3668
rect 118 3662 121 3778
rect 126 3762 129 3768
rect 134 3762 137 3838
rect 142 3792 145 3948
rect 158 3942 161 3948
rect 166 3892 169 3948
rect 174 3942 177 3978
rect 182 3902 185 3928
rect 182 3892 185 3898
rect 150 3852 153 3888
rect 158 3872 161 3878
rect 174 3872 177 3888
rect 190 3882 193 4038
rect 206 3982 209 3988
rect 198 3962 201 3968
rect 214 3941 217 4058
rect 230 3992 233 4018
rect 238 4002 241 4218
rect 246 4162 249 4238
rect 326 4232 329 4378
rect 390 4372 393 4478
rect 414 4462 417 4518
rect 494 4492 497 4518
rect 510 4482 513 4538
rect 518 4532 521 4538
rect 438 4472 441 4478
rect 450 4468 454 4471
rect 494 4462 497 4468
rect 434 4458 438 4461
rect 482 4458 486 4461
rect 398 4452 401 4458
rect 406 4442 409 4458
rect 426 4448 433 4451
rect 466 4448 470 4451
rect 406 4432 409 4438
rect 378 4358 382 4361
rect 342 4352 345 4358
rect 358 4352 361 4358
rect 370 4348 374 4351
rect 394 4348 398 4351
rect 334 4342 337 4348
rect 406 4342 409 4348
rect 414 4342 417 4398
rect 430 4392 433 4448
rect 494 4402 497 4458
rect 494 4362 497 4378
rect 466 4348 470 4351
rect 350 4292 353 4338
rect 366 4332 369 4338
rect 462 4322 465 4338
rect 470 4332 473 4338
rect 490 4328 494 4331
rect 510 4322 513 4478
rect 518 4471 521 4528
rect 526 4512 529 4548
rect 534 4542 537 4598
rect 582 4572 585 4578
rect 566 4552 569 4558
rect 542 4542 545 4548
rect 550 4542 553 4548
rect 578 4538 582 4541
rect 518 4468 529 4471
rect 526 4462 529 4468
rect 518 4452 521 4458
rect 526 4452 529 4458
rect 534 4442 537 4448
rect 526 4391 529 4418
rect 518 4388 529 4391
rect 518 4352 521 4388
rect 526 4372 529 4378
rect 534 4342 537 4428
rect 522 4338 529 4341
rect 382 4282 385 4318
rect 494 4312 497 4318
rect 410 4278 414 4281
rect 374 4272 377 4278
rect 362 4268 366 4271
rect 370 4258 374 4261
rect 246 4152 249 4158
rect 254 4072 257 4138
rect 262 4132 265 4178
rect 286 4152 289 4158
rect 294 4152 297 4228
rect 328 4203 330 4207
rect 334 4203 337 4207
rect 341 4203 344 4207
rect 358 4192 361 4248
rect 382 4242 385 4248
rect 390 4212 393 4268
rect 402 4228 406 4231
rect 286 4142 289 4148
rect 310 4142 313 4148
rect 278 4132 281 4138
rect 326 4132 329 4168
rect 270 4092 273 4128
rect 286 4062 289 4068
rect 306 4058 310 4061
rect 274 4048 281 4051
rect 254 4042 257 4048
rect 222 3972 225 3978
rect 234 3958 238 3961
rect 254 3952 257 4008
rect 270 3992 273 4038
rect 278 3992 281 4048
rect 286 4002 289 4058
rect 318 4052 321 4098
rect 342 4092 345 4148
rect 350 4132 353 4138
rect 366 4072 369 4188
rect 390 4182 393 4208
rect 374 4152 377 4158
rect 414 4152 417 4268
rect 422 4262 425 4278
rect 430 4272 433 4278
rect 450 4268 454 4271
rect 422 4242 425 4258
rect 390 4142 393 4148
rect 382 4092 385 4118
rect 390 4082 393 4088
rect 358 4062 361 4068
rect 342 4052 345 4058
rect 374 4052 377 4058
rect 294 4038 302 4041
rect 294 3992 297 4038
rect 310 4032 313 4038
rect 398 4022 401 4078
rect 414 4072 417 4078
rect 422 4062 425 4238
rect 430 4172 433 4268
rect 462 4262 465 4278
rect 486 4272 489 4298
rect 526 4292 529 4338
rect 534 4292 537 4338
rect 542 4332 545 4528
rect 590 4522 593 4568
rect 598 4552 601 4578
rect 606 4562 609 4658
rect 614 4652 617 4668
rect 626 4658 630 4661
rect 614 4632 617 4638
rect 622 4632 625 4638
rect 614 4572 617 4628
rect 622 4592 625 4608
rect 638 4592 641 4668
rect 646 4652 649 4718
rect 662 4702 665 4758
rect 670 4752 673 4818
rect 670 4692 673 4738
rect 654 4582 657 4658
rect 678 4652 681 4748
rect 686 4692 689 4918
rect 702 4912 705 4958
rect 718 4922 721 4938
rect 694 4882 697 4888
rect 694 4852 697 4868
rect 702 4842 705 4858
rect 702 4742 705 4838
rect 694 4712 697 4728
rect 710 4682 713 4788
rect 726 4722 729 4958
rect 734 4932 737 4948
rect 734 4872 737 4928
rect 750 4912 753 5058
rect 830 5052 833 5058
rect 838 5052 841 5068
rect 874 5058 878 5061
rect 786 5048 790 5051
rect 758 5042 761 5048
rect 822 5042 825 5048
rect 862 4982 865 5048
rect 894 5002 897 5068
rect 774 4942 777 4978
rect 834 4968 838 4971
rect 882 4968 886 4971
rect 846 4962 849 4968
rect 894 4962 897 4978
rect 902 4962 905 4968
rect 794 4958 801 4961
rect 790 4942 793 4948
rect 762 4938 766 4941
rect 782 4932 785 4938
rect 758 4892 761 4928
rect 766 4882 769 4908
rect 782 4892 785 4918
rect 798 4892 801 4958
rect 814 4942 817 4958
rect 830 4952 833 4958
rect 918 4952 921 5048
rect 926 5022 929 5068
rect 1054 5062 1057 5068
rect 934 5022 937 5048
rect 942 5032 945 5048
rect 1038 5032 1041 5059
rect 1070 5052 1073 5058
rect 1094 5052 1097 5128
rect 1126 5082 1129 5088
rect 1134 5072 1137 5088
rect 1118 5062 1121 5068
rect 1182 5062 1185 5068
rect 1190 5062 1193 5068
rect 1078 5042 1081 5048
rect 1094 5042 1097 5048
rect 934 4962 937 5018
rect 942 5012 945 5028
rect 838 4948 846 4951
rect 826 4938 830 4941
rect 838 4932 841 4948
rect 818 4878 822 4881
rect 734 4762 737 4838
rect 734 4732 737 4748
rect 742 4742 745 4858
rect 766 4832 769 4878
rect 774 4862 777 4868
rect 806 4862 809 4868
rect 794 4858 798 4861
rect 774 4792 777 4828
rect 754 4758 758 4761
rect 750 4732 753 4738
rect 734 4682 737 4718
rect 782 4711 785 4858
rect 810 4848 814 4851
rect 838 4832 841 4928
rect 848 4903 850 4907
rect 854 4903 857 4907
rect 861 4903 864 4907
rect 870 4892 873 4938
rect 918 4882 921 4938
rect 934 4932 937 4938
rect 926 4922 929 4928
rect 942 4892 945 4998
rect 958 4982 961 4988
rect 950 4962 953 4968
rect 950 4902 953 4918
rect 922 4878 926 4881
rect 802 4778 806 4781
rect 814 4772 817 4808
rect 814 4762 817 4768
rect 830 4752 833 4768
rect 846 4762 849 4848
rect 854 4762 857 4868
rect 862 4862 865 4878
rect 950 4862 953 4868
rect 874 4858 878 4861
rect 890 4858 894 4861
rect 862 4832 865 4858
rect 886 4842 889 4858
rect 874 4818 878 4821
rect 926 4792 929 4858
rect 914 4768 918 4771
rect 846 4752 849 4758
rect 950 4752 953 4788
rect 958 4782 961 4798
rect 798 4742 801 4748
rect 814 4742 817 4748
rect 854 4742 857 4748
rect 826 4738 830 4741
rect 918 4742 921 4748
rect 790 4722 793 4738
rect 822 4722 825 4738
rect 886 4732 889 4740
rect 898 4738 902 4741
rect 906 4728 913 4731
rect 858 4718 862 4721
rect 778 4708 785 4711
rect 738 4668 742 4671
rect 762 4668 766 4671
rect 774 4662 777 4708
rect 848 4703 850 4707
rect 854 4703 857 4707
rect 861 4703 864 4707
rect 822 4682 825 4688
rect 886 4682 889 4688
rect 874 4678 878 4681
rect 826 4668 830 4671
rect 690 4658 694 4661
rect 754 4658 758 4661
rect 718 4652 721 4658
rect 662 4632 665 4638
rect 610 4558 614 4561
rect 670 4552 673 4618
rect 678 4552 681 4568
rect 686 4552 689 4638
rect 694 4632 697 4638
rect 702 4622 705 4628
rect 742 4562 745 4568
rect 618 4538 625 4541
rect 602 4518 609 4521
rect 566 4502 569 4518
rect 574 4472 577 4488
rect 590 4482 593 4498
rect 598 4482 601 4508
rect 582 4472 585 4478
rect 554 4468 558 4471
rect 550 4422 553 4458
rect 582 4452 585 4458
rect 562 4448 566 4451
rect 550 4392 553 4398
rect 570 4358 574 4361
rect 510 4281 513 4288
rect 510 4278 518 4281
rect 542 4272 545 4328
rect 530 4268 534 4271
rect 478 4262 481 4268
rect 490 4258 494 4261
rect 438 4252 441 4258
rect 550 4252 553 4318
rect 558 4312 561 4348
rect 582 4342 585 4358
rect 598 4352 601 4478
rect 606 4402 609 4518
rect 614 4452 617 4458
rect 622 4382 625 4538
rect 638 4522 641 4548
rect 662 4532 665 4538
rect 630 4502 633 4518
rect 630 4462 633 4488
rect 638 4472 641 4508
rect 670 4472 673 4488
rect 638 4452 641 4468
rect 650 4458 654 4461
rect 678 4452 681 4498
rect 646 4432 649 4448
rect 686 4442 689 4548
rect 702 4532 705 4558
rect 710 4542 713 4548
rect 758 4542 761 4628
rect 766 4552 769 4618
rect 694 4522 697 4528
rect 702 4472 705 4528
rect 766 4472 769 4548
rect 774 4472 777 4658
rect 790 4552 793 4648
rect 798 4562 801 4668
rect 822 4642 825 4648
rect 806 4552 809 4558
rect 782 4532 785 4548
rect 782 4482 785 4518
rect 722 4468 726 4471
rect 774 4462 777 4468
rect 790 4462 793 4548
rect 814 4542 817 4548
rect 830 4542 833 4658
rect 842 4638 846 4641
rect 854 4632 857 4648
rect 858 4538 862 4541
rect 798 4492 801 4518
rect 806 4482 809 4538
rect 802 4468 806 4471
rect 698 4458 702 4461
rect 706 4448 710 4451
rect 718 4442 721 4458
rect 766 4452 769 4458
rect 814 4452 817 4538
rect 822 4522 825 4528
rect 830 4512 833 4518
rect 826 4468 830 4471
rect 822 4452 825 4458
rect 662 4362 665 4418
rect 686 4392 689 4438
rect 702 4372 705 4398
rect 610 4358 614 4361
rect 610 4348 614 4351
rect 566 4332 569 4338
rect 590 4312 593 4338
rect 598 4322 601 4338
rect 622 4332 625 4358
rect 638 4352 641 4358
rect 646 4352 649 4358
rect 662 4352 665 4358
rect 702 4352 705 4368
rect 478 4222 481 4248
rect 470 4192 473 4198
rect 494 4192 497 4208
rect 534 4192 537 4248
rect 550 4192 553 4208
rect 558 4192 561 4308
rect 598 4292 601 4318
rect 570 4278 574 4281
rect 582 4278 590 4281
rect 566 4242 569 4268
rect 566 4192 569 4228
rect 582 4212 585 4278
rect 606 4272 609 4278
rect 590 4262 593 4268
rect 630 4262 633 4318
rect 646 4282 649 4318
rect 662 4302 665 4348
rect 726 4342 729 4398
rect 742 4362 745 4418
rect 750 4362 753 4428
rect 682 4338 686 4341
rect 670 4331 673 4338
rect 670 4328 681 4331
rect 690 4328 694 4331
rect 714 4328 718 4331
rect 662 4272 665 4288
rect 670 4262 673 4268
rect 678 4262 681 4328
rect 734 4322 737 4348
rect 766 4341 769 4448
rect 830 4442 833 4458
rect 806 4362 809 4368
rect 778 4348 782 4351
rect 766 4338 777 4341
rect 754 4318 758 4321
rect 686 4272 689 4298
rect 694 4272 697 4278
rect 702 4272 705 4278
rect 710 4272 713 4318
rect 766 4312 769 4318
rect 722 4288 726 4291
rect 610 4258 614 4261
rect 682 4258 686 4261
rect 626 4238 630 4241
rect 702 4182 705 4268
rect 714 4258 718 4261
rect 710 4222 713 4258
rect 726 4251 729 4268
rect 734 4262 737 4288
rect 742 4272 745 4278
rect 754 4268 758 4271
rect 722 4248 729 4251
rect 602 4168 606 4171
rect 650 4168 654 4171
rect 478 4162 481 4168
rect 506 4158 510 4161
rect 478 4142 481 4158
rect 438 4102 441 4128
rect 462 4082 465 4088
rect 414 4042 417 4048
rect 422 4041 425 4048
rect 430 4041 433 4058
rect 422 4038 433 4041
rect 438 4042 441 4068
rect 478 4062 481 4068
rect 458 4058 462 4061
rect 470 4042 473 4048
rect 486 4042 489 4058
rect 328 4003 330 4007
rect 334 4003 337 4007
rect 341 4003 344 4007
rect 318 3992 321 3998
rect 406 3992 409 4018
rect 430 3992 433 4038
rect 454 4032 457 4038
rect 226 3948 230 3951
rect 214 3938 225 3941
rect 198 3932 201 3938
rect 222 3922 225 3938
rect 222 3892 225 3918
rect 254 3892 257 3938
rect 278 3892 281 3958
rect 286 3942 289 3968
rect 298 3958 302 3961
rect 314 3958 318 3961
rect 302 3952 305 3958
rect 230 3872 233 3878
rect 194 3868 198 3871
rect 294 3871 297 3948
rect 326 3942 329 3988
rect 366 3972 369 3978
rect 358 3962 361 3968
rect 374 3962 377 3978
rect 406 3962 409 3988
rect 418 3968 422 3971
rect 438 3962 441 4008
rect 494 3982 497 4148
rect 518 4142 521 4148
rect 506 4138 510 4141
rect 526 4132 529 4168
rect 574 4162 577 4168
rect 538 4148 542 4151
rect 582 4142 585 4148
rect 554 4128 558 4131
rect 502 4092 505 4128
rect 518 4092 521 4108
rect 542 4092 545 4118
rect 590 4092 593 4158
rect 614 4152 617 4168
rect 626 4158 630 4161
rect 662 4161 665 4178
rect 678 4162 681 4168
rect 662 4158 673 4161
rect 670 4152 673 4158
rect 658 4148 662 4151
rect 546 4078 550 4081
rect 510 4022 513 4078
rect 534 4062 537 4068
rect 550 4062 553 4068
rect 558 4062 561 4078
rect 574 4072 577 4088
rect 522 4058 526 4061
rect 458 3968 462 3971
rect 502 3962 505 4008
rect 542 3992 545 4038
rect 574 3992 577 4058
rect 598 4051 601 4118
rect 622 4092 625 4138
rect 634 4128 638 4131
rect 606 4072 609 4088
rect 646 4071 649 4128
rect 678 4092 681 4118
rect 686 4092 689 4138
rect 694 4112 697 4148
rect 702 4092 705 4168
rect 710 4102 713 4138
rect 718 4092 721 4208
rect 750 4192 753 4258
rect 730 4158 734 4161
rect 758 4152 761 4158
rect 766 4152 769 4308
rect 774 4292 777 4338
rect 782 4292 785 4348
rect 790 4292 793 4358
rect 802 4348 806 4351
rect 822 4342 825 4408
rect 838 4392 841 4528
rect 848 4503 850 4507
rect 854 4503 857 4507
rect 861 4503 864 4507
rect 870 4492 873 4658
rect 894 4592 897 4668
rect 902 4592 905 4708
rect 902 4522 905 4548
rect 854 4441 857 4488
rect 890 4468 894 4471
rect 866 4458 870 4461
rect 874 4448 878 4451
rect 886 4442 889 4458
rect 894 4442 897 4448
rect 854 4438 862 4441
rect 862 4392 865 4418
rect 882 4348 886 4351
rect 834 4338 838 4341
rect 814 4332 817 4338
rect 798 4272 801 4328
rect 810 4258 814 4261
rect 774 4252 777 4258
rect 782 4252 785 4258
rect 814 4212 817 4228
rect 814 4192 817 4198
rect 754 4138 758 4141
rect 790 4122 793 4148
rect 822 4132 825 4338
rect 848 4303 850 4307
rect 854 4303 857 4307
rect 861 4303 864 4307
rect 874 4288 878 4291
rect 858 4268 862 4271
rect 838 4262 841 4268
rect 874 4258 878 4261
rect 870 4242 873 4248
rect 854 4192 857 4218
rect 878 4212 881 4238
rect 886 4162 889 4328
rect 894 4321 897 4338
rect 902 4332 905 4518
rect 910 4502 913 4728
rect 926 4702 929 4728
rect 942 4722 945 4738
rect 958 4732 961 4778
rect 966 4721 969 4958
rect 974 4952 977 4968
rect 982 4942 985 4958
rect 990 4942 993 4948
rect 1006 4942 1009 4968
rect 1046 4962 1049 5008
rect 1014 4942 1017 4958
rect 1062 4952 1065 4958
rect 982 4932 985 4938
rect 1014 4892 1017 4938
rect 1002 4888 1006 4891
rect 974 4842 977 4868
rect 982 4862 985 4878
rect 1006 4862 1009 4878
rect 1022 4862 1025 4868
rect 998 4858 1006 4861
rect 998 4852 1001 4858
rect 1030 4842 1033 4858
rect 1038 4841 1041 4938
rect 1046 4882 1049 4948
rect 1170 4948 1174 4951
rect 1134 4942 1137 4947
rect 1170 4938 1174 4941
rect 1054 4892 1057 4928
rect 1074 4918 1078 4921
rect 1150 4892 1153 4938
rect 1182 4892 1185 5058
rect 1198 5051 1201 5128
rect 1230 5082 1233 5088
rect 1234 5068 1238 5071
rect 1274 5068 1278 5071
rect 1246 5052 1249 5068
rect 1274 5058 1278 5061
rect 1190 5048 1201 5051
rect 1050 4878 1054 4881
rect 1082 4868 1086 4871
rect 1178 4868 1182 4871
rect 1082 4858 1086 4861
rect 1082 4848 1086 4851
rect 1034 4838 1041 4841
rect 974 4792 977 4838
rect 1094 4832 1097 4858
rect 1102 4842 1105 4848
rect 1034 4828 1038 4831
rect 982 4762 985 4778
rect 1018 4768 1022 4771
rect 1038 4762 1041 4768
rect 986 4748 990 4751
rect 1034 4748 1038 4751
rect 974 4732 977 4748
rect 958 4718 969 4721
rect 934 4702 937 4718
rect 958 4692 961 4718
rect 938 4688 942 4691
rect 966 4682 969 4688
rect 950 4672 953 4678
rect 918 4662 921 4668
rect 938 4658 942 4661
rect 934 4622 937 4648
rect 918 4532 921 4558
rect 926 4542 929 4558
rect 942 4542 945 4558
rect 950 4552 953 4558
rect 966 4541 969 4668
rect 990 4662 993 4698
rect 998 4682 1001 4748
rect 1006 4702 1009 4738
rect 1018 4718 1022 4721
rect 1046 4712 1049 4758
rect 1094 4752 1097 4818
rect 1118 4812 1121 4848
rect 1126 4832 1129 4858
rect 1154 4848 1158 4851
rect 1134 4842 1137 4848
rect 1166 4832 1169 4868
rect 1178 4858 1182 4861
rect 1190 4851 1193 5048
rect 1222 4962 1225 4968
rect 1230 4952 1233 5048
rect 1254 5002 1257 5058
rect 1262 4972 1265 5018
rect 1270 4962 1273 5048
rect 1278 4952 1281 4998
rect 1294 4962 1297 4968
rect 1334 4952 1337 5038
rect 1342 4992 1345 5068
rect 1406 5062 1409 5068
rect 1352 5003 1354 5007
rect 1358 5003 1361 5007
rect 1365 5003 1368 5007
rect 1350 4962 1353 4968
rect 1306 4948 1310 4951
rect 1198 4922 1201 4948
rect 1222 4942 1225 4948
rect 1270 4932 1273 4938
rect 1250 4928 1254 4931
rect 1202 4918 1209 4921
rect 1206 4852 1209 4918
rect 1214 4872 1217 4878
rect 1222 4862 1225 4928
rect 1270 4892 1273 4928
rect 1234 4878 1238 4881
rect 1234 4868 1238 4871
rect 1230 4862 1233 4868
rect 1190 4848 1198 4851
rect 1182 4842 1185 4848
rect 1126 4792 1129 4818
rect 1158 4782 1161 4818
rect 1158 4762 1161 4768
rect 1102 4752 1105 4758
rect 1146 4748 1153 4751
rect 1054 4732 1057 4738
rect 1070 4732 1073 4738
rect 998 4672 1001 4678
rect 1006 4652 1009 4668
rect 978 4648 982 4651
rect 1014 4622 1017 4628
rect 1022 4622 1025 4668
rect 1042 4658 1046 4661
rect 1034 4648 1038 4651
rect 1030 4612 1033 4648
rect 1054 4641 1057 4708
rect 1078 4692 1081 4748
rect 1110 4742 1113 4748
rect 1138 4738 1142 4741
rect 1098 4728 1102 4731
rect 1130 4728 1134 4731
rect 1150 4722 1153 4748
rect 1158 4732 1161 4738
rect 1086 4702 1089 4718
rect 1102 4682 1105 4698
rect 1074 4658 1078 4661
rect 1098 4658 1102 4661
rect 1050 4638 1057 4641
rect 1062 4642 1065 4648
rect 1102 4642 1105 4648
rect 1054 4632 1057 4638
rect 1078 4632 1081 4638
rect 962 4538 969 4541
rect 974 4532 977 4538
rect 934 4482 937 4498
rect 918 4402 921 4458
rect 934 4392 937 4458
rect 942 4452 945 4518
rect 966 4472 969 4518
rect 982 4492 985 4578
rect 1038 4562 1041 4618
rect 1046 4562 1049 4578
rect 1070 4561 1073 4618
rect 1110 4582 1113 4658
rect 1118 4592 1121 4718
rect 1126 4662 1129 4698
rect 1134 4682 1137 4698
rect 1134 4672 1137 4678
rect 1142 4672 1145 4678
rect 1158 4662 1161 4688
rect 1166 4671 1169 4758
rect 1182 4752 1185 4778
rect 1174 4742 1177 4748
rect 1190 4742 1193 4848
rect 1238 4772 1241 4818
rect 1246 4762 1249 4828
rect 1198 4752 1201 4758
rect 1246 4752 1249 4758
rect 1190 4732 1193 4738
rect 1182 4692 1185 4728
rect 1198 4682 1201 4748
rect 1206 4742 1209 4748
rect 1178 4678 1182 4681
rect 1166 4668 1177 4671
rect 1158 4652 1161 4658
rect 1118 4572 1121 4578
rect 1062 4558 1073 4561
rect 1106 4568 1110 4571
rect 1018 4538 1022 4541
rect 1030 4541 1033 4548
rect 1062 4542 1065 4558
rect 1078 4542 1081 4568
rect 1126 4562 1129 4648
rect 1118 4552 1121 4558
rect 1030 4538 1038 4541
rect 1070 4532 1073 4538
rect 990 4522 993 4528
rect 978 4478 982 4481
rect 986 4468 990 4471
rect 950 4462 953 4468
rect 998 4452 1001 4458
rect 958 4442 961 4448
rect 950 4422 953 4428
rect 922 4368 926 4371
rect 950 4362 953 4388
rect 970 4368 974 4371
rect 934 4342 937 4348
rect 942 4322 945 4358
rect 962 4348 966 4351
rect 958 4332 961 4338
rect 974 4332 977 4338
rect 982 4332 985 4388
rect 1006 4352 1009 4398
rect 1014 4372 1017 4508
rect 1070 4472 1073 4478
rect 1046 4462 1049 4468
rect 1034 4458 1038 4461
rect 1014 4342 1017 4368
rect 1030 4342 1033 4368
rect 1078 4362 1081 4528
rect 1094 4471 1097 4518
rect 1126 4492 1129 4558
rect 1134 4542 1137 4588
rect 1146 4558 1150 4561
rect 1162 4558 1166 4561
rect 1174 4552 1177 4668
rect 1182 4552 1185 4568
rect 1190 4562 1193 4678
rect 1206 4672 1209 4738
rect 1222 4672 1225 4718
rect 1174 4532 1177 4548
rect 1198 4541 1201 4658
rect 1206 4652 1209 4668
rect 1230 4662 1233 4728
rect 1238 4702 1241 4748
rect 1246 4712 1249 4718
rect 1238 4672 1241 4698
rect 1246 4672 1249 4678
rect 1206 4562 1209 4648
rect 1230 4642 1233 4658
rect 1246 4652 1249 4658
rect 1230 4592 1233 4618
rect 1254 4612 1257 4868
rect 1326 4862 1329 4918
rect 1278 4762 1281 4818
rect 1334 4772 1337 4948
rect 1342 4902 1345 4948
rect 1374 4932 1377 5059
rect 1382 4932 1385 5028
rect 1438 4992 1441 5128
rect 1462 5092 1465 5128
rect 1542 5128 1554 5131
rect 1662 5128 1666 5132
rect 1894 5128 1898 5132
rect 1542 5092 1545 5128
rect 1662 5102 1665 5128
rect 1872 5103 1874 5107
rect 1878 5103 1881 5107
rect 1885 5103 1888 5107
rect 1730 5078 1734 5081
rect 1822 5072 1825 5078
rect 1538 5068 1542 5071
rect 1586 5068 1590 5071
rect 1666 5068 1670 5071
rect 1738 5068 1742 5071
rect 1474 5058 1478 5061
rect 1482 5058 1489 5061
rect 1350 4882 1353 4888
rect 1382 4872 1385 4928
rect 1390 4872 1393 4958
rect 1454 4952 1457 4968
rect 1410 4948 1414 4951
rect 1434 4948 1438 4951
rect 1398 4932 1401 4938
rect 1406 4902 1409 4938
rect 1414 4882 1417 4948
rect 1422 4892 1425 4898
rect 1430 4892 1433 4928
rect 1470 4892 1473 4948
rect 1486 4942 1489 5058
rect 1570 5058 1574 5061
rect 1558 4992 1561 5058
rect 1654 5012 1657 5018
rect 1654 4992 1657 4998
rect 1546 4968 1550 4971
rect 1590 4952 1593 4958
rect 1710 4952 1713 4958
rect 1514 4948 1518 4951
rect 1730 4948 1734 4951
rect 1494 4942 1497 4948
rect 1486 4892 1489 4938
rect 1590 4882 1593 4948
rect 1614 4932 1617 4948
rect 1474 4878 1478 4881
rect 1654 4872 1657 4938
rect 1742 4892 1745 5068
rect 1802 5058 1806 5061
rect 1846 5002 1849 5058
rect 1806 4912 1809 4948
rect 1894 4942 1897 5128
rect 2888 5103 2890 5107
rect 2894 5103 2897 5107
rect 2901 5103 2904 5107
rect 3920 5103 3922 5107
rect 3926 5103 3929 5107
rect 3933 5103 3936 5107
rect 4936 5103 4938 5107
rect 4942 5103 4945 5107
rect 4949 5103 4952 5107
rect 2306 5088 2310 5091
rect 2618 5088 2622 5091
rect 4146 5088 4150 5091
rect 2454 5082 2457 5088
rect 2526 5082 2529 5088
rect 4238 5082 4241 5088
rect 4486 5082 4489 5088
rect 2426 5078 2430 5081
rect 2466 5078 2470 5081
rect 4498 5078 4502 5081
rect 1934 5072 1937 5078
rect 2126 5072 2129 5078
rect 2410 5068 2414 5071
rect 2442 5068 2446 5071
rect 1982 5062 1985 5068
rect 2058 5058 2062 5061
rect 2222 5062 2225 5068
rect 2246 5062 2249 5068
rect 2318 5062 2321 5068
rect 1906 5018 1910 5021
rect 1942 4992 1945 4998
rect 1922 4958 1926 4961
rect 1934 4951 1937 4958
rect 1934 4948 1942 4951
rect 1898 4938 1902 4941
rect 1898 4928 1902 4931
rect 1862 4922 1865 4928
rect 1874 4918 1878 4921
rect 1726 4872 1729 4888
rect 1442 4866 1446 4869
rect 1498 4868 1502 4871
rect 1454 4862 1457 4868
rect 1458 4858 1462 4861
rect 1578 4858 1582 4861
rect 1352 4803 1354 4807
rect 1358 4803 1361 4807
rect 1365 4803 1368 4807
rect 1406 4792 1409 4858
rect 1314 4758 1318 4761
rect 1278 4752 1281 4758
rect 1266 4748 1270 4751
rect 1298 4748 1302 4751
rect 1334 4751 1337 4758
rect 1326 4748 1337 4751
rect 1270 4732 1273 4738
rect 1266 4688 1270 4691
rect 1278 4671 1281 4748
rect 1286 4702 1289 4738
rect 1302 4732 1305 4738
rect 1310 4672 1313 4698
rect 1318 4672 1321 4678
rect 1278 4668 1289 4671
rect 1270 4632 1273 4668
rect 1278 4592 1281 4658
rect 1286 4652 1289 4668
rect 1314 4658 1318 4661
rect 1302 4642 1305 4658
rect 1326 4652 1329 4748
rect 1306 4618 1310 4621
rect 1238 4562 1241 4568
rect 1294 4562 1297 4608
rect 1302 4582 1305 4588
rect 1306 4568 1310 4571
rect 1218 4558 1222 4561
rect 1210 4548 1214 4551
rect 1266 4548 1270 4551
rect 1198 4538 1206 4541
rect 1242 4538 1246 4541
rect 1090 4468 1097 4471
rect 1086 4442 1089 4468
rect 1098 4458 1102 4461
rect 1114 4458 1118 4461
rect 1098 4448 1102 4451
rect 1106 4438 1110 4441
rect 1102 4392 1105 4428
rect 1042 4348 1046 4351
rect 1094 4342 1097 4388
rect 1110 4381 1113 4418
rect 1134 4382 1137 4478
rect 1142 4472 1145 4478
rect 1150 4472 1153 4518
rect 1158 4512 1161 4518
rect 1166 4492 1169 4518
rect 1174 4512 1177 4528
rect 1182 4522 1185 4538
rect 1178 4468 1182 4471
rect 1110 4378 1121 4381
rect 1110 4332 1113 4368
rect 1118 4352 1121 4378
rect 1134 4362 1137 4378
rect 1150 4372 1153 4468
rect 1158 4462 1161 4468
rect 1158 4352 1161 4458
rect 1166 4452 1169 4468
rect 1182 4452 1185 4458
rect 1190 4452 1193 4538
rect 1206 4462 1209 4538
rect 1214 4522 1217 4538
rect 1242 4528 1246 4531
rect 1254 4522 1257 4548
rect 1222 4482 1225 4488
rect 1214 4452 1217 4468
rect 1222 4452 1225 4458
rect 1230 4402 1233 4518
rect 1254 4481 1257 4518
rect 1250 4478 1257 4481
rect 1262 4492 1265 4538
rect 1278 4522 1281 4548
rect 1262 4482 1265 4488
rect 1242 4468 1246 4471
rect 1254 4462 1257 4478
rect 1270 4461 1273 4518
rect 1294 4482 1297 4558
rect 1310 4492 1313 4558
rect 1318 4552 1321 4618
rect 1326 4562 1329 4648
rect 1334 4642 1337 4738
rect 1342 4732 1345 4738
rect 1358 4692 1361 4788
rect 1366 4742 1369 4778
rect 1386 4768 1390 4771
rect 1366 4692 1369 4738
rect 1382 4692 1385 4738
rect 1342 4682 1345 4688
rect 1366 4642 1369 4678
rect 1402 4668 1406 4671
rect 1410 4658 1414 4661
rect 1326 4502 1329 4558
rect 1334 4532 1337 4638
rect 1366 4622 1369 4638
rect 1352 4603 1354 4607
rect 1358 4603 1361 4607
rect 1365 4603 1368 4607
rect 1370 4548 1374 4551
rect 1338 4518 1342 4521
rect 1326 4482 1329 4488
rect 1350 4482 1353 4548
rect 1382 4542 1385 4588
rect 1358 4532 1361 4538
rect 1382 4532 1385 4538
rect 1358 4492 1361 4528
rect 1398 4522 1401 4658
rect 1406 4642 1409 4648
rect 1422 4642 1425 4668
rect 1414 4632 1417 4638
rect 1422 4592 1425 4638
rect 1430 4562 1433 4818
rect 1502 4792 1505 4858
rect 1654 4822 1657 4868
rect 1662 4862 1665 4868
rect 1742 4862 1745 4868
rect 1854 4862 1857 4918
rect 1862 4892 1865 4908
rect 1872 4903 1874 4907
rect 1878 4903 1881 4907
rect 1885 4903 1888 4907
rect 1914 4888 1921 4891
rect 1910 4872 1913 4888
rect 1770 4858 1774 4861
rect 1882 4858 1886 4861
rect 1510 4752 1513 4818
rect 1518 4752 1521 4778
rect 1574 4752 1577 4758
rect 1530 4748 1534 4751
rect 1618 4748 1622 4751
rect 1446 4742 1449 4747
rect 1462 4732 1465 4738
rect 1438 4692 1441 4698
rect 1462 4682 1465 4688
rect 1406 4522 1409 4548
rect 1382 4492 1385 4518
rect 1282 4478 1286 4481
rect 1314 4478 1318 4481
rect 1266 4458 1273 4461
rect 1286 4452 1289 4468
rect 1294 4462 1297 4468
rect 1254 4442 1257 4448
rect 1302 4412 1305 4458
rect 1146 4348 1150 4351
rect 894 4318 905 4321
rect 902 4292 905 4318
rect 958 4292 961 4318
rect 918 4192 921 4268
rect 926 4262 929 4278
rect 974 4262 977 4328
rect 982 4272 985 4278
rect 990 4272 993 4318
rect 954 4258 958 4261
rect 1014 4252 1017 4328
rect 1030 4292 1033 4328
rect 1038 4282 1041 4328
rect 1026 4268 1030 4271
rect 1022 4252 1025 4258
rect 954 4248 958 4251
rect 946 4238 950 4241
rect 842 4148 846 4151
rect 638 4068 649 4071
rect 706 4068 710 4071
rect 614 4062 617 4068
rect 638 4052 641 4068
rect 670 4062 673 4068
rect 594 4048 601 4051
rect 514 3988 518 3991
rect 610 3988 614 3991
rect 466 3958 470 3961
rect 374 3952 377 3958
rect 526 3952 529 3978
rect 598 3972 601 3978
rect 562 3968 566 3971
rect 582 3962 585 3968
rect 622 3962 625 3978
rect 630 3952 633 4048
rect 638 4002 641 4048
rect 646 3992 649 4058
rect 658 4038 662 4041
rect 662 4022 665 4028
rect 678 3972 681 4068
rect 686 4042 689 4048
rect 678 3962 681 3968
rect 686 3952 689 4038
rect 694 4012 697 4058
rect 718 4052 721 4088
rect 766 4082 769 4088
rect 726 4072 729 4078
rect 694 3992 697 4008
rect 702 3982 705 4018
rect 702 3952 705 3968
rect 694 3948 702 3951
rect 326 3912 329 3938
rect 290 3868 297 3871
rect 170 3858 201 3861
rect 158 3782 161 3858
rect 198 3841 201 3858
rect 206 3852 209 3858
rect 214 3841 217 3848
rect 198 3838 217 3841
rect 126 3672 129 3678
rect 134 3652 137 3758
rect 206 3742 209 3798
rect 142 3682 145 3698
rect 106 3558 110 3561
rect 130 3548 134 3551
rect 70 3542 73 3547
rect 118 3542 121 3548
rect 86 3532 89 3538
rect 6 3462 9 3468
rect 22 3342 25 3418
rect 10 3338 14 3341
rect 10 3288 14 3291
rect 22 3142 25 3338
rect 62 3302 65 3318
rect 70 3282 73 3528
rect 86 3521 89 3528
rect 102 3522 105 3528
rect 86 3518 97 3521
rect 94 3492 97 3518
rect 130 3468 134 3471
rect 78 3362 81 3368
rect 110 3352 113 3448
rect 118 3372 121 3418
rect 98 3348 102 3351
rect 142 3342 145 3678
rect 150 3672 153 3738
rect 198 3732 201 3738
rect 190 3692 193 3718
rect 198 3712 201 3728
rect 206 3702 209 3738
rect 214 3732 217 3740
rect 222 3692 225 3818
rect 230 3792 233 3868
rect 262 3862 265 3868
rect 238 3832 241 3858
rect 286 3852 289 3868
rect 302 3852 305 3908
rect 354 3878 358 3881
rect 366 3872 369 3948
rect 390 3942 393 3948
rect 406 3942 409 3948
rect 430 3942 433 3948
rect 378 3938 382 3941
rect 318 3862 321 3868
rect 366 3862 369 3868
rect 374 3862 377 3888
rect 262 3842 265 3848
rect 250 3788 254 3791
rect 230 3752 233 3788
rect 194 3678 198 3681
rect 246 3672 249 3768
rect 254 3762 257 3768
rect 178 3668 182 3671
rect 210 3668 214 3671
rect 150 3652 153 3668
rect 254 3662 257 3748
rect 262 3742 265 3838
rect 278 3832 281 3848
rect 310 3842 313 3858
rect 278 3792 281 3808
rect 310 3802 313 3838
rect 318 3791 321 3858
rect 328 3803 330 3807
rect 334 3803 337 3807
rect 341 3803 344 3807
rect 318 3788 326 3791
rect 278 3762 281 3778
rect 278 3752 281 3758
rect 294 3742 297 3758
rect 310 3742 313 3758
rect 270 3672 273 3738
rect 298 3728 302 3731
rect 318 3672 321 3738
rect 350 3732 353 3828
rect 358 3792 361 3858
rect 374 3852 377 3858
rect 366 3752 369 3818
rect 362 3748 366 3751
rect 374 3742 377 3838
rect 382 3832 385 3868
rect 390 3822 393 3858
rect 406 3852 409 3928
rect 446 3922 449 3938
rect 454 3932 457 3948
rect 430 3892 433 3908
rect 470 3892 473 3938
rect 478 3922 481 3938
rect 486 3932 489 3948
rect 510 3932 513 3948
rect 550 3932 553 3948
rect 574 3942 577 3948
rect 438 3872 441 3878
rect 486 3872 489 3878
rect 502 3872 505 3918
rect 510 3892 513 3928
rect 526 3922 529 3928
rect 526 3892 529 3918
rect 406 3772 409 3848
rect 414 3762 417 3848
rect 422 3792 425 3868
rect 450 3848 454 3851
rect 462 3841 465 3858
rect 494 3852 497 3858
rect 518 3852 521 3878
rect 534 3862 537 3878
rect 566 3872 569 3908
rect 582 3892 585 3948
rect 606 3942 609 3948
rect 638 3922 641 3948
rect 646 3932 649 3938
rect 630 3882 633 3888
rect 594 3878 598 3881
rect 574 3872 577 3878
rect 654 3862 657 3918
rect 686 3912 689 3928
rect 694 3872 697 3948
rect 702 3862 705 3938
rect 726 3932 729 3978
rect 734 3972 737 4018
rect 734 3942 737 3948
rect 746 3938 750 3941
rect 710 3872 713 3878
rect 454 3838 465 3841
rect 474 3838 478 3841
rect 390 3742 393 3758
rect 398 3752 401 3758
rect 418 3748 422 3751
rect 326 3672 329 3708
rect 170 3658 174 3661
rect 202 3658 206 3661
rect 262 3622 265 3658
rect 150 3552 153 3558
rect 158 3552 161 3558
rect 158 3492 161 3538
rect 174 3532 177 3538
rect 198 3482 201 3538
rect 206 3532 209 3548
rect 166 3462 169 3468
rect 206 3462 209 3468
rect 114 3338 118 3341
rect 70 3263 73 3268
rect 86 3262 89 3338
rect 102 3331 105 3338
rect 102 3328 113 3331
rect 110 3292 113 3328
rect 102 3282 105 3288
rect 118 3272 121 3338
rect 110 3192 113 3218
rect 70 3142 73 3148
rect 86 3142 89 3148
rect 10 3138 14 3141
rect 6 3072 9 3138
rect 102 3111 105 3147
rect 94 3108 105 3111
rect 94 3092 97 3108
rect 126 3082 129 3118
rect 78 3062 81 3078
rect 86 3062 89 3068
rect 158 3062 161 3418
rect 166 3382 169 3388
rect 222 3362 225 3508
rect 246 3502 249 3618
rect 294 3612 297 3618
rect 328 3603 330 3607
rect 334 3603 337 3607
rect 341 3603 344 3607
rect 374 3602 377 3738
rect 398 3732 401 3738
rect 446 3732 449 3768
rect 406 3692 409 3698
rect 430 3692 433 3728
rect 446 3702 449 3728
rect 454 3682 457 3838
rect 462 3832 465 3838
rect 470 3752 473 3818
rect 478 3762 481 3818
rect 462 3722 465 3748
rect 550 3742 553 3748
rect 566 3742 569 3748
rect 486 3712 489 3738
rect 590 3732 593 3748
rect 598 3712 601 3818
rect 630 3772 633 3858
rect 702 3832 705 3858
rect 718 3852 721 3918
rect 750 3863 753 3928
rect 758 3922 761 3948
rect 766 3892 769 3928
rect 642 3768 646 3771
rect 758 3752 761 3868
rect 662 3742 665 3748
rect 678 3732 681 3747
rect 758 3742 761 3748
rect 646 3692 649 3728
rect 474 3688 478 3691
rect 566 3682 569 3688
rect 674 3678 678 3681
rect 398 3672 401 3678
rect 426 3668 430 3671
rect 446 3662 449 3668
rect 394 3658 398 3661
rect 418 3658 425 3661
rect 262 3542 265 3548
rect 302 3542 305 3558
rect 326 3542 329 3548
rect 306 3538 310 3541
rect 258 3518 262 3521
rect 286 3482 289 3538
rect 314 3528 318 3531
rect 326 3492 329 3538
rect 342 3532 345 3548
rect 366 3542 369 3568
rect 422 3562 425 3658
rect 462 3612 465 3678
rect 526 3662 529 3678
rect 590 3672 593 3678
rect 582 3662 585 3668
rect 638 3662 641 3668
rect 686 3662 689 3708
rect 742 3682 745 3718
rect 754 3678 758 3681
rect 718 3662 721 3678
rect 774 3672 777 3938
rect 782 3872 785 4068
rect 798 4063 801 4118
rect 814 4062 817 4128
rect 830 4062 833 4148
rect 848 4103 850 4107
rect 854 4103 857 4107
rect 861 4103 864 4107
rect 870 4092 873 4138
rect 894 4132 897 4168
rect 878 4062 881 4078
rect 902 4062 905 4138
rect 910 4072 913 4168
rect 974 4142 977 4168
rect 1046 4151 1049 4288
rect 1054 4282 1057 4308
rect 1086 4282 1089 4318
rect 1134 4292 1137 4328
rect 1174 4292 1177 4368
rect 1186 4358 1190 4361
rect 1186 4348 1190 4351
rect 1222 4342 1225 4358
rect 1246 4342 1249 4408
rect 1310 4392 1313 4478
rect 1350 4452 1353 4458
rect 1374 4452 1377 4478
rect 1390 4472 1393 4488
rect 1414 4462 1417 4558
rect 1438 4552 1441 4638
rect 1454 4552 1457 4668
rect 1430 4501 1433 4538
rect 1454 4512 1457 4548
rect 1462 4542 1465 4678
rect 1470 4562 1473 4688
rect 1478 4572 1481 4618
rect 1486 4561 1489 4748
rect 1478 4558 1489 4561
rect 1470 4552 1473 4558
rect 1478 4552 1481 4558
rect 1502 4552 1505 4558
rect 1466 4538 1470 4541
rect 1430 4498 1438 4501
rect 1438 4462 1441 4498
rect 1446 4462 1449 4468
rect 1470 4462 1473 4468
rect 1466 4458 1470 4461
rect 1378 4448 1382 4451
rect 1426 4438 1430 4441
rect 1326 4372 1329 4418
rect 1352 4403 1354 4407
rect 1358 4403 1361 4407
rect 1365 4403 1368 4407
rect 1182 4282 1185 4338
rect 1246 4332 1249 4338
rect 1198 4292 1201 4318
rect 1098 4278 1102 4281
rect 1078 4262 1081 4268
rect 1102 4262 1105 4268
rect 1118 4262 1121 4268
rect 1142 4262 1145 4268
rect 1066 4258 1070 4261
rect 1086 4232 1089 4238
rect 1126 4232 1129 4248
rect 1150 4232 1153 4268
rect 1162 4258 1166 4261
rect 1182 4222 1185 4278
rect 1190 4272 1193 4278
rect 1254 4262 1257 4358
rect 1326 4352 1329 4358
rect 1262 4332 1265 4338
rect 1310 4292 1313 4348
rect 1382 4342 1385 4348
rect 1390 4342 1393 4398
rect 1414 4352 1417 4398
rect 1406 4342 1409 4348
rect 1326 4272 1329 4328
rect 1358 4282 1361 4318
rect 1346 4278 1350 4281
rect 1298 4268 1302 4271
rect 1326 4262 1329 4268
rect 1382 4262 1385 4338
rect 1078 4172 1081 4218
rect 1246 4192 1249 4258
rect 1170 4168 1174 4171
rect 1206 4162 1209 4168
rect 1166 4158 1182 4161
rect 1166 4152 1169 4158
rect 1222 4152 1225 4158
rect 1246 4152 1249 4178
rect 1114 4148 1118 4151
rect 1178 4148 1182 4151
rect 922 4138 926 4141
rect 946 4118 950 4121
rect 918 4072 921 4118
rect 982 4082 985 4118
rect 942 4062 945 4068
rect 998 4062 1001 4068
rect 914 4058 918 4061
rect 838 4052 841 4058
rect 882 4048 886 4051
rect 938 4048 942 4051
rect 902 4042 905 4048
rect 950 4042 953 4058
rect 990 4042 993 4058
rect 838 3952 841 4008
rect 854 3982 857 4018
rect 934 3972 937 4038
rect 898 3948 902 3951
rect 790 3902 793 3948
rect 798 3942 801 3948
rect 838 3942 841 3948
rect 958 3942 961 3958
rect 978 3948 982 3951
rect 966 3942 969 3948
rect 806 3922 809 3928
rect 822 3922 825 3928
rect 822 3892 825 3918
rect 848 3903 850 3907
rect 854 3903 857 3907
rect 861 3903 864 3907
rect 846 3862 849 3868
rect 870 3862 873 3878
rect 886 3872 889 3928
rect 990 3922 993 3958
rect 954 3918 958 3921
rect 918 3892 921 3908
rect 930 3888 934 3891
rect 910 3752 913 3868
rect 918 3752 921 3888
rect 954 3878 958 3881
rect 970 3878 974 3881
rect 938 3868 942 3871
rect 982 3862 985 3868
rect 938 3858 942 3861
rect 990 3852 993 3898
rect 850 3748 854 3751
rect 882 3748 886 3751
rect 734 3662 737 3668
rect 782 3662 785 3748
rect 790 3742 793 3748
rect 910 3742 913 3748
rect 934 3742 937 3748
rect 874 3738 878 3741
rect 918 3732 921 3738
rect 894 3722 897 3728
rect 842 3718 846 3721
rect 506 3658 510 3661
rect 610 3658 614 3661
rect 658 3658 662 3661
rect 762 3658 766 3661
rect 510 3592 513 3658
rect 590 3652 593 3658
rect 622 3652 625 3658
rect 490 3568 494 3571
rect 386 3558 390 3561
rect 434 3548 438 3551
rect 486 3541 489 3558
rect 542 3552 545 3568
rect 566 3562 569 3568
rect 514 3548 518 3551
rect 494 3541 497 3548
rect 526 3542 529 3548
rect 486 3538 497 3541
rect 506 3538 510 3541
rect 390 3532 393 3538
rect 342 3522 345 3528
rect 274 3468 278 3471
rect 286 3462 289 3478
rect 298 3468 302 3471
rect 298 3458 302 3461
rect 270 3452 273 3458
rect 306 3448 310 3451
rect 262 3442 265 3448
rect 246 3391 249 3438
rect 318 3432 321 3458
rect 342 3422 345 3468
rect 406 3462 409 3538
rect 442 3488 446 3491
rect 386 3458 390 3461
rect 328 3403 330 3407
rect 334 3403 337 3407
rect 341 3403 344 3407
rect 246 3388 257 3391
rect 178 3338 182 3341
rect 194 3318 198 3321
rect 190 3252 193 3268
rect 206 3262 209 3358
rect 222 3342 225 3358
rect 254 3342 257 3388
rect 350 3372 353 3378
rect 262 3352 265 3368
rect 318 3362 321 3368
rect 374 3362 377 3368
rect 390 3352 393 3428
rect 406 3421 409 3458
rect 406 3418 417 3421
rect 214 3272 217 3318
rect 210 3258 217 3261
rect 198 3252 201 3258
rect 174 3172 177 3218
rect 214 3162 217 3258
rect 182 3142 185 3148
rect 198 3132 201 3147
rect 166 3112 169 3118
rect 166 3092 169 3108
rect 182 3092 185 3128
rect 214 3082 217 3118
rect 222 3102 225 3218
rect 278 3192 281 3278
rect 286 3272 289 3338
rect 290 3258 294 3261
rect 334 3222 337 3348
rect 398 3342 401 3418
rect 414 3342 417 3418
rect 438 3352 441 3418
rect 342 3302 345 3338
rect 398 3322 401 3338
rect 414 3321 417 3338
rect 406 3318 417 3321
rect 382 3262 385 3308
rect 406 3272 409 3318
rect 446 3302 449 3468
rect 454 3462 457 3498
rect 478 3492 481 3528
rect 458 3418 462 3421
rect 454 3292 457 3408
rect 470 3401 473 3448
rect 478 3412 481 3448
rect 470 3398 481 3401
rect 478 3332 481 3398
rect 438 3272 441 3288
rect 450 3278 454 3281
rect 474 3258 478 3261
rect 486 3222 489 3538
rect 542 3532 545 3548
rect 550 3532 553 3558
rect 590 3552 593 3608
rect 630 3582 633 3658
rect 610 3548 614 3551
rect 626 3548 630 3551
rect 566 3532 569 3548
rect 638 3542 641 3658
rect 702 3652 705 3658
rect 726 3652 729 3658
rect 662 3552 665 3628
rect 662 3542 665 3548
rect 678 3542 681 3588
rect 762 3568 766 3571
rect 774 3552 777 3638
rect 782 3622 785 3658
rect 798 3592 801 3668
rect 818 3659 822 3662
rect 790 3562 793 3568
rect 706 3548 710 3551
rect 806 3551 809 3618
rect 806 3548 814 3551
rect 582 3492 585 3538
rect 766 3532 769 3538
rect 658 3518 662 3521
rect 510 3472 513 3478
rect 502 3462 505 3468
rect 526 3462 529 3468
rect 494 3452 497 3458
rect 518 3442 521 3458
rect 542 3452 545 3488
rect 546 3448 550 3451
rect 558 3432 561 3458
rect 498 3378 502 3381
rect 558 3362 561 3368
rect 566 3362 569 3468
rect 574 3452 577 3478
rect 594 3458 598 3461
rect 502 3352 505 3358
rect 574 3352 577 3428
rect 606 3422 609 3518
rect 662 3463 665 3468
rect 598 3402 601 3418
rect 614 3362 617 3398
rect 550 3342 553 3348
rect 590 3342 593 3358
rect 602 3348 609 3351
rect 514 3338 518 3341
rect 582 3332 585 3338
rect 554 3328 558 3331
rect 518 3312 521 3318
rect 534 3312 537 3328
rect 534 3272 537 3308
rect 558 3282 561 3288
rect 558 3232 561 3259
rect 494 3222 497 3228
rect 328 3203 330 3207
rect 334 3203 337 3207
rect 341 3203 344 3207
rect 298 3148 302 3151
rect 230 3112 233 3138
rect 258 3118 262 3121
rect 218 3068 222 3071
rect 174 3062 177 3068
rect 106 3058 110 3061
rect 62 2942 65 3018
rect 70 2932 73 2947
rect 10 2918 14 2921
rect 42 2858 46 2861
rect 62 2752 65 2858
rect 86 2852 89 3058
rect 158 3052 161 3058
rect 142 2962 145 3018
rect 166 2972 169 3058
rect 198 3052 201 3058
rect 126 2942 129 2948
rect 102 2922 105 2928
rect 98 2888 102 2891
rect 110 2882 113 2918
rect 142 2872 145 2958
rect 150 2922 153 2948
rect 222 2942 225 2948
rect 166 2892 169 2928
rect 206 2902 209 2918
rect 110 2862 113 2868
rect 158 2862 161 2868
rect 182 2862 185 2878
rect 214 2872 217 2918
rect 146 2858 150 2861
rect 42 2748 46 2751
rect 62 2742 65 2748
rect 62 2662 65 2738
rect 94 2682 97 2688
rect 102 2672 105 2838
rect 134 2832 137 2858
rect 110 2792 113 2828
rect 182 2822 185 2858
rect 190 2852 193 2858
rect 198 2842 201 2868
rect 206 2862 209 2868
rect 118 2752 121 2818
rect 130 2748 134 2751
rect 42 2658 46 2661
rect 38 2552 41 2558
rect 62 2552 65 2658
rect 90 2578 94 2581
rect 62 2462 65 2548
rect 102 2542 105 2668
rect 110 2662 113 2668
rect 118 2622 121 2738
rect 142 2692 145 2758
rect 158 2732 161 2738
rect 150 2672 153 2688
rect 130 2668 134 2671
rect 126 2652 129 2658
rect 150 2652 153 2668
rect 162 2658 166 2661
rect 134 2622 137 2648
rect 134 2572 137 2578
rect 110 2562 113 2568
rect 126 2562 129 2568
rect 114 2548 118 2551
rect 102 2532 105 2538
rect 94 2472 97 2488
rect 102 2472 105 2528
rect 134 2512 137 2568
rect 114 2458 118 2461
rect 38 2452 41 2458
rect 62 2352 65 2458
rect 122 2448 126 2451
rect 142 2451 145 2618
rect 150 2562 153 2568
rect 158 2551 161 2588
rect 154 2548 161 2551
rect 150 2502 153 2548
rect 174 2542 177 2728
rect 182 2662 185 2708
rect 198 2692 201 2748
rect 194 2678 198 2681
rect 206 2672 209 2848
rect 222 2742 225 2938
rect 246 2932 249 2948
rect 230 2852 233 2898
rect 270 2871 273 3078
rect 278 2992 281 3118
rect 310 3092 313 3148
rect 326 3142 329 3168
rect 414 3152 417 3218
rect 562 3168 566 3171
rect 342 3142 345 3147
rect 374 3102 377 3138
rect 358 3072 361 3078
rect 270 2868 278 2871
rect 246 2852 249 2858
rect 254 2842 257 2868
rect 262 2801 265 2868
rect 270 2862 273 2868
rect 274 2848 278 2851
rect 254 2798 265 2801
rect 238 2682 241 2718
rect 226 2678 230 2681
rect 182 2592 185 2658
rect 190 2542 193 2668
rect 246 2662 249 2668
rect 254 2662 257 2798
rect 286 2772 289 3058
rect 294 2982 297 3058
rect 302 3022 305 3068
rect 326 3022 329 3058
rect 328 3003 330 3007
rect 334 3003 337 3007
rect 341 3003 344 3007
rect 310 2952 313 2958
rect 374 2952 377 3088
rect 390 3082 393 3108
rect 398 3062 401 3128
rect 406 3072 409 3118
rect 414 3082 417 3148
rect 422 3142 425 3148
rect 446 3142 449 3148
rect 502 3142 505 3148
rect 434 3128 438 3131
rect 406 2992 409 3068
rect 446 3062 449 3138
rect 462 3091 465 3128
rect 478 3112 481 3138
rect 482 3108 489 3111
rect 458 3088 465 3091
rect 486 3082 489 3108
rect 494 3062 497 3088
rect 510 3072 513 3158
rect 582 3152 585 3158
rect 566 3122 569 3128
rect 574 3112 577 3118
rect 558 3052 561 3058
rect 454 2982 457 3018
rect 318 2942 321 2948
rect 350 2942 353 2948
rect 326 2922 329 2928
rect 302 2912 305 2918
rect 342 2882 345 2898
rect 322 2878 326 2881
rect 294 2852 297 2878
rect 310 2842 313 2858
rect 282 2748 286 2751
rect 270 2742 273 2748
rect 270 2702 273 2738
rect 318 2722 321 2868
rect 350 2862 353 2938
rect 374 2912 377 2928
rect 370 2868 374 2871
rect 358 2862 361 2868
rect 362 2848 366 2851
rect 328 2803 330 2807
rect 334 2803 337 2807
rect 341 2803 344 2807
rect 338 2778 342 2781
rect 358 2742 361 2838
rect 382 2832 385 2858
rect 390 2812 393 2938
rect 398 2922 401 2928
rect 406 2911 409 2928
rect 398 2908 409 2911
rect 398 2892 401 2908
rect 438 2872 441 2928
rect 446 2902 449 2948
rect 534 2942 537 3038
rect 574 3032 577 3078
rect 554 3028 558 3031
rect 494 2882 497 2888
rect 502 2882 505 2918
rect 534 2912 537 2938
rect 542 2932 545 2948
rect 562 2888 566 2891
rect 534 2882 537 2888
rect 530 2868 534 2871
rect 398 2842 401 2848
rect 382 2772 385 2778
rect 270 2672 273 2678
rect 302 2672 305 2718
rect 306 2668 313 2671
rect 234 2658 238 2661
rect 198 2552 201 2558
rect 214 2552 217 2658
rect 158 2482 161 2538
rect 138 2448 145 2451
rect 150 2452 153 2468
rect 158 2452 161 2458
rect 110 2442 113 2448
rect 122 2348 126 2351
rect 38 2332 41 2348
rect 38 2262 41 2278
rect 62 2262 65 2348
rect 134 2342 137 2448
rect 142 2362 145 2418
rect 150 2352 153 2438
rect 158 2352 161 2358
rect 142 2342 145 2348
rect 122 2338 126 2341
rect 150 2292 153 2348
rect 166 2341 169 2518
rect 174 2462 177 2498
rect 214 2482 217 2538
rect 222 2522 225 2658
rect 274 2638 278 2641
rect 258 2568 262 2571
rect 274 2558 278 2561
rect 274 2548 278 2551
rect 262 2532 265 2538
rect 262 2502 265 2528
rect 182 2472 185 2478
rect 286 2472 289 2658
rect 302 2572 305 2658
rect 294 2562 297 2568
rect 294 2532 297 2558
rect 310 2492 313 2668
rect 318 2552 321 2708
rect 350 2682 353 2698
rect 350 2663 353 2668
rect 328 2603 330 2607
rect 334 2603 337 2607
rect 341 2603 344 2607
rect 358 2582 361 2738
rect 366 2712 369 2748
rect 382 2722 385 2768
rect 390 2742 393 2748
rect 406 2742 409 2748
rect 430 2742 433 2868
rect 446 2862 449 2868
rect 502 2862 505 2868
rect 574 2862 577 2878
rect 582 2872 585 3148
rect 590 3142 593 3298
rect 598 3292 601 3318
rect 606 3182 609 3348
rect 614 3331 617 3358
rect 622 3352 625 3408
rect 638 3352 641 3458
rect 638 3332 641 3348
rect 670 3332 673 3347
rect 678 3342 681 3468
rect 694 3462 697 3468
rect 694 3412 697 3448
rect 710 3442 713 3458
rect 718 3402 721 3468
rect 738 3378 742 3381
rect 750 3362 753 3368
rect 742 3352 745 3358
rect 614 3328 622 3331
rect 630 3312 633 3318
rect 614 3212 617 3258
rect 622 3252 625 3298
rect 654 3292 657 3328
rect 678 3292 681 3338
rect 742 3332 745 3348
rect 750 3342 753 3358
rect 758 3332 761 3478
rect 766 3462 769 3518
rect 774 3482 777 3548
rect 798 3542 801 3548
rect 774 3372 777 3458
rect 806 3402 809 3548
rect 822 3542 825 3588
rect 830 3552 833 3558
rect 830 3492 833 3538
rect 838 3531 841 3718
rect 848 3703 850 3707
rect 854 3703 857 3707
rect 861 3703 864 3707
rect 846 3672 849 3688
rect 878 3682 881 3688
rect 886 3552 889 3708
rect 926 3662 929 3698
rect 942 3672 945 3758
rect 974 3742 977 3747
rect 958 3692 961 3738
rect 958 3672 961 3678
rect 998 3672 1001 3988
rect 1006 3952 1009 4108
rect 1030 4072 1033 4138
rect 1046 4082 1049 4088
rect 1030 3992 1033 4038
rect 1062 3972 1065 3978
rect 1046 3962 1049 3968
rect 1078 3962 1081 3998
rect 1094 3962 1097 4088
rect 1126 4072 1129 4148
rect 1226 4138 1230 4141
rect 1174 4122 1177 4138
rect 1230 4132 1233 4138
rect 1238 4122 1241 4138
rect 1110 4052 1113 4059
rect 1058 3948 1062 3951
rect 1030 3942 1033 3948
rect 1014 3932 1017 3938
rect 1006 3862 1009 3868
rect 1006 3842 1009 3848
rect 1014 3832 1017 3928
rect 1022 3912 1025 3938
rect 1054 3932 1057 3938
rect 1078 3882 1081 3918
rect 1054 3872 1057 3878
rect 1094 3872 1097 3958
rect 1126 3952 1129 4068
rect 1150 4062 1153 4068
rect 1174 4062 1177 4098
rect 1190 4072 1193 4078
rect 1170 4058 1174 4061
rect 1130 3948 1134 3951
rect 1110 3872 1113 3918
rect 1118 3892 1121 3948
rect 1066 3858 1070 3861
rect 1038 3842 1041 3858
rect 1046 3852 1049 3858
rect 1078 3852 1081 3868
rect 1086 3852 1089 3858
rect 1094 3852 1097 3858
rect 1022 3802 1025 3818
rect 1054 3792 1057 3848
rect 1102 3802 1105 3858
rect 1094 3742 1097 3748
rect 970 3668 974 3671
rect 998 3662 1001 3668
rect 970 3658 974 3661
rect 910 3642 913 3648
rect 894 3552 897 3618
rect 918 3552 921 3658
rect 938 3648 942 3651
rect 950 3642 953 3658
rect 1006 3652 1009 3728
rect 1014 3672 1017 3678
rect 1030 3672 1033 3688
rect 1070 3672 1073 3738
rect 1110 3712 1113 3868
rect 1134 3862 1137 3918
rect 1142 3912 1145 4058
rect 1150 3992 1153 4058
rect 1158 4052 1161 4058
rect 1222 4042 1225 4059
rect 1222 3952 1225 3968
rect 1230 3952 1233 4068
rect 1238 3932 1241 4118
rect 1246 4092 1249 4148
rect 1254 4142 1257 4258
rect 1270 4238 1278 4241
rect 1282 4238 1286 4241
rect 1270 4162 1273 4238
rect 1294 4182 1297 4258
rect 1366 4252 1369 4258
rect 1352 4203 1354 4207
rect 1358 4203 1361 4207
rect 1365 4203 1368 4207
rect 1286 4152 1289 4158
rect 1382 4152 1385 4218
rect 1254 4062 1257 4138
rect 1286 4112 1289 4148
rect 1294 4132 1297 4138
rect 1310 4132 1313 4138
rect 1326 4122 1329 4147
rect 1390 4132 1393 4338
rect 1446 4332 1449 4458
rect 1466 4448 1470 4451
rect 1470 4352 1473 4358
rect 1442 4318 1446 4321
rect 1438 4282 1441 4288
rect 1418 4278 1422 4281
rect 1398 4272 1401 4278
rect 1426 4268 1430 4271
rect 1410 4258 1414 4261
rect 1422 4242 1425 4258
rect 1310 4092 1313 4118
rect 1290 4088 1294 4091
rect 1302 4062 1305 4068
rect 1334 4061 1337 4128
rect 1386 4118 1390 4121
rect 1358 4082 1361 4118
rect 1330 4058 1337 4061
rect 1342 4062 1345 4078
rect 1370 4068 1374 4071
rect 1390 4062 1393 4088
rect 1398 4072 1401 4178
rect 1414 4132 1417 4168
rect 1438 4152 1441 4278
rect 1446 4262 1449 4268
rect 1454 4262 1457 4318
rect 1446 4182 1449 4258
rect 1470 4192 1473 4248
rect 1478 4212 1481 4548
rect 1498 4538 1502 4541
rect 1510 4512 1513 4748
rect 1534 4672 1537 4678
rect 1550 4662 1553 4718
rect 1558 4702 1561 4748
rect 1566 4742 1569 4748
rect 1582 4742 1585 4748
rect 1598 4732 1601 4738
rect 1566 4682 1569 4728
rect 1606 4722 1609 4728
rect 1570 4659 1574 4662
rect 1590 4662 1593 4718
rect 1630 4712 1633 4818
rect 1654 4752 1657 4798
rect 1646 4742 1649 4748
rect 1638 4722 1641 4728
rect 1646 4722 1649 4738
rect 1646 4692 1649 4698
rect 1662 4672 1665 4858
rect 1838 4792 1841 4818
rect 1846 4782 1849 4858
rect 1854 4782 1857 4858
rect 1862 4792 1865 4858
rect 1802 4748 1806 4751
rect 1674 4738 1678 4741
rect 1678 4702 1681 4728
rect 1686 4692 1689 4748
rect 1598 4662 1601 4668
rect 1574 4552 1577 4558
rect 1542 4542 1545 4547
rect 1486 4482 1489 4488
rect 1526 4472 1529 4538
rect 1578 4488 1582 4491
rect 1518 4452 1521 4459
rect 1590 4452 1593 4518
rect 1606 4462 1609 4608
rect 1662 4562 1665 4668
rect 1682 4659 1686 4662
rect 1694 4592 1697 4748
rect 1726 4742 1729 4748
rect 1830 4742 1833 4748
rect 1710 4652 1713 4658
rect 1614 4552 1617 4558
rect 1654 4542 1657 4547
rect 1662 4542 1665 4558
rect 1726 4552 1729 4708
rect 1742 4692 1745 4698
rect 1758 4672 1761 4718
rect 1782 4682 1785 4728
rect 1798 4682 1801 4688
rect 1774 4662 1777 4668
rect 1782 4662 1785 4668
rect 1750 4632 1753 4658
rect 1814 4652 1817 4668
rect 1846 4662 1849 4778
rect 1854 4752 1857 4758
rect 1870 4751 1873 4788
rect 1878 4762 1881 4858
rect 1870 4748 1878 4751
rect 1886 4732 1889 4748
rect 1898 4738 1902 4741
rect 1872 4703 1874 4707
rect 1878 4703 1881 4707
rect 1885 4703 1888 4707
rect 1890 4688 1894 4691
rect 1918 4672 1921 4888
rect 1830 4652 1833 4659
rect 1742 4602 1745 4618
rect 1742 4582 1745 4588
rect 1638 4492 1641 4538
rect 1686 4502 1689 4508
rect 1686 4492 1689 4498
rect 1718 4482 1721 4518
rect 1614 4472 1617 4478
rect 1670 4472 1673 4478
rect 1626 4468 1630 4471
rect 1586 4448 1590 4451
rect 1566 4352 1569 4448
rect 1598 4382 1601 4458
rect 1614 4362 1617 4468
rect 1654 4462 1657 4468
rect 1626 4458 1630 4461
rect 1702 4442 1705 4458
rect 1622 4362 1625 4368
rect 1594 4358 1598 4361
rect 1490 4348 1494 4351
rect 1538 4348 1542 4351
rect 1566 4342 1569 4348
rect 1518 4291 1521 4338
rect 1542 4332 1545 4338
rect 1558 4322 1561 4328
rect 1518 4288 1529 4291
rect 1510 4272 1513 4278
rect 1526 4272 1529 4288
rect 1550 4272 1553 4318
rect 1486 4262 1489 4268
rect 1542 4263 1545 4268
rect 1502 4242 1505 4258
rect 1498 4218 1502 4221
rect 1486 4162 1489 4168
rect 1446 4158 1454 4161
rect 1438 4142 1441 4148
rect 1294 4042 1297 4058
rect 1286 4002 1289 4018
rect 1302 4012 1305 4058
rect 1352 4003 1354 4007
rect 1358 4003 1361 4007
rect 1365 4003 1368 4007
rect 1274 3988 1278 3991
rect 1286 3972 1289 3978
rect 1310 3962 1313 3988
rect 1350 3972 1353 3978
rect 1374 3952 1377 3958
rect 1382 3952 1385 4058
rect 1422 4052 1425 4118
rect 1446 4092 1449 4158
rect 1462 4152 1465 4158
rect 1502 4152 1505 4208
rect 1510 4192 1513 4258
rect 1566 4192 1569 4338
rect 1574 4302 1577 4348
rect 1582 4332 1585 4338
rect 1590 4312 1593 4358
rect 1618 4348 1622 4351
rect 1606 4342 1609 4348
rect 1682 4348 1686 4351
rect 1654 4342 1657 4347
rect 1598 4332 1601 4338
rect 1506 4148 1510 4151
rect 1454 4138 1462 4141
rect 1430 4072 1433 4078
rect 1454 4072 1457 4138
rect 1470 4131 1473 4148
rect 1462 4128 1473 4131
rect 1462 4112 1465 4128
rect 1394 4048 1398 4051
rect 1446 4042 1449 4048
rect 1406 3961 1409 4018
rect 1454 3992 1457 4068
rect 1462 4062 1465 4108
rect 1462 3982 1465 4058
rect 1478 4052 1481 4078
rect 1518 4071 1521 4138
rect 1526 4132 1529 4188
rect 1550 4152 1553 4178
rect 1574 4162 1577 4298
rect 1606 4292 1609 4298
rect 1610 4268 1614 4271
rect 1622 4262 1625 4298
rect 1662 4292 1665 4298
rect 1674 4278 1678 4281
rect 1654 4272 1657 4278
rect 1566 4132 1569 4138
rect 1534 4122 1537 4128
rect 1566 4118 1574 4121
rect 1534 4092 1537 4108
rect 1566 4082 1569 4118
rect 1558 4078 1566 4081
rect 1514 4068 1521 4071
rect 1530 4068 1534 4071
rect 1502 4062 1505 4068
rect 1502 4042 1505 4048
rect 1510 4022 1513 4068
rect 1518 3992 1521 4038
rect 1502 3962 1505 3978
rect 1406 3958 1414 3961
rect 1502 3952 1505 3958
rect 1290 3948 1294 3951
rect 1330 3948 1334 3951
rect 1514 3948 1518 3951
rect 1394 3938 1398 3941
rect 1278 3932 1281 3938
rect 1174 3912 1177 3918
rect 1142 3782 1145 3908
rect 1150 3882 1153 3908
rect 1174 3882 1177 3888
rect 1202 3878 1206 3881
rect 1150 3862 1153 3878
rect 1182 3872 1185 3878
rect 1214 3872 1217 3908
rect 1222 3862 1225 3878
rect 1238 3872 1241 3878
rect 1246 3862 1249 3908
rect 1334 3902 1337 3938
rect 1334 3872 1337 3878
rect 1382 3872 1385 3878
rect 1318 3863 1321 3868
rect 1178 3858 1182 3861
rect 1194 3858 1201 3861
rect 1154 3768 1158 3771
rect 1158 3752 1161 3758
rect 1174 3752 1177 3798
rect 1190 3742 1193 3758
rect 1198 3752 1201 3858
rect 1366 3862 1369 3868
rect 1414 3862 1417 3948
rect 1422 3872 1425 3878
rect 1378 3858 1382 3861
rect 1206 3852 1209 3858
rect 1254 3842 1257 3848
rect 1226 3818 1230 3821
rect 1206 3752 1209 3768
rect 1214 3742 1217 3788
rect 1238 3752 1241 3768
rect 1222 3742 1225 3748
rect 1162 3738 1166 3741
rect 1250 3738 1254 3741
rect 1118 3732 1121 3738
rect 1182 3722 1185 3738
rect 1190 3692 1193 3708
rect 1254 3702 1257 3718
rect 1262 3692 1265 3858
rect 1398 3852 1401 3858
rect 1352 3803 1354 3807
rect 1358 3803 1361 3807
rect 1365 3803 1368 3807
rect 1374 3752 1377 3778
rect 1414 3772 1417 3858
rect 1422 3832 1425 3868
rect 1430 3852 1433 3918
rect 1438 3772 1441 3898
rect 1446 3891 1449 3938
rect 1470 3932 1473 3948
rect 1486 3942 1489 3948
rect 1510 3932 1513 3938
rect 1454 3902 1457 3918
rect 1486 3892 1489 3928
rect 1526 3922 1529 4068
rect 1550 4062 1553 4068
rect 1534 3962 1537 4028
rect 1558 3952 1561 4078
rect 1582 4072 1585 4138
rect 1606 4092 1609 4128
rect 1622 4122 1625 4218
rect 1630 4112 1633 4148
rect 1606 4082 1609 4088
rect 1598 4062 1601 4068
rect 1574 4042 1577 4048
rect 1590 4012 1593 4058
rect 1622 3952 1625 4038
rect 1542 3942 1545 3948
rect 1598 3942 1601 3948
rect 1546 3928 1550 3931
rect 1446 3888 1457 3891
rect 1454 3872 1457 3888
rect 1486 3882 1489 3888
rect 1446 3832 1449 3858
rect 1454 3822 1457 3868
rect 1462 3862 1465 3878
rect 1558 3871 1561 3938
rect 1598 3882 1601 3888
rect 1626 3878 1630 3881
rect 1554 3868 1561 3871
rect 1546 3858 1550 3861
rect 1626 3858 1630 3861
rect 1446 3802 1449 3818
rect 1470 3812 1473 3818
rect 1454 3772 1457 3788
rect 1482 3768 1486 3771
rect 1310 3742 1313 3748
rect 1386 3738 1390 3741
rect 1302 3732 1305 3738
rect 1146 3688 1150 3691
rect 1110 3682 1113 3688
rect 1242 3678 1246 3681
rect 1114 3668 1118 3671
rect 886 3542 889 3548
rect 858 3538 862 3541
rect 906 3538 910 3541
rect 838 3528 846 3531
rect 906 3528 910 3531
rect 870 3522 873 3528
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 861 3503 864 3507
rect 870 3492 873 3518
rect 878 3492 881 3498
rect 902 3492 905 3508
rect 818 3488 822 3491
rect 918 3482 921 3548
rect 926 3542 929 3598
rect 954 3588 958 3591
rect 966 3542 969 3638
rect 1046 3622 1049 3659
rect 994 3618 998 3621
rect 1054 3592 1057 3598
rect 1018 3568 1022 3571
rect 994 3558 998 3561
rect 974 3552 977 3558
rect 1050 3548 1054 3551
rect 818 3478 822 3481
rect 890 3478 894 3481
rect 914 3468 918 3471
rect 914 3458 918 3461
rect 774 3342 777 3368
rect 798 3342 801 3348
rect 838 3342 841 3458
rect 862 3452 865 3458
rect 926 3442 929 3458
rect 862 3352 865 3418
rect 702 3302 705 3328
rect 638 3262 641 3278
rect 638 3242 641 3248
rect 646 3202 649 3268
rect 670 3262 673 3268
rect 654 3242 657 3248
rect 678 3242 681 3268
rect 686 3202 689 3268
rect 694 3262 697 3278
rect 742 3272 745 3308
rect 758 3282 761 3328
rect 774 3292 777 3338
rect 854 3322 857 3338
rect 862 3332 865 3348
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 861 3303 864 3307
rect 774 3282 777 3288
rect 850 3278 854 3281
rect 734 3262 737 3268
rect 710 3242 713 3248
rect 734 3232 737 3238
rect 626 3168 630 3171
rect 638 3152 641 3178
rect 706 3158 710 3161
rect 602 3148 606 3151
rect 674 3148 678 3151
rect 690 3148 694 3151
rect 610 3138 614 3141
rect 590 3132 593 3138
rect 594 3088 598 3091
rect 598 3062 601 3068
rect 606 3062 609 3128
rect 614 3062 617 3068
rect 622 3062 625 3148
rect 678 3142 681 3148
rect 718 3142 721 3148
rect 742 3142 745 3268
rect 774 3242 777 3259
rect 838 3242 841 3248
rect 870 3242 873 3438
rect 886 3342 889 3358
rect 926 3342 929 3348
rect 898 3328 902 3331
rect 910 3282 913 3328
rect 886 3262 889 3278
rect 910 3252 913 3258
rect 918 3252 921 3258
rect 934 3232 937 3518
rect 966 3502 969 3538
rect 1006 3512 1009 3548
rect 1038 3542 1041 3548
rect 1070 3542 1073 3668
rect 1126 3642 1129 3658
rect 1142 3632 1145 3648
rect 1150 3642 1153 3668
rect 1158 3662 1161 3678
rect 1270 3672 1273 3678
rect 1250 3668 1254 3671
rect 1206 3662 1209 3668
rect 1178 3648 1182 3651
rect 1166 3592 1169 3608
rect 1154 3588 1158 3591
rect 1094 3552 1097 3568
rect 1102 3552 1105 3568
rect 1158 3552 1161 3558
rect 1182 3542 1185 3628
rect 1190 3602 1193 3658
rect 1222 3642 1225 3658
rect 1246 3652 1249 3658
rect 1278 3622 1281 3668
rect 1286 3662 1289 3698
rect 1358 3692 1361 3738
rect 1310 3682 1313 3688
rect 1310 3672 1313 3678
rect 1358 3672 1361 3688
rect 1298 3668 1302 3671
rect 1306 3648 1310 3651
rect 1366 3632 1369 3738
rect 1398 3702 1401 3758
rect 1414 3752 1417 3768
rect 1418 3738 1422 3741
rect 1438 3741 1441 3768
rect 1502 3752 1505 3858
rect 1606 3852 1609 3858
rect 1638 3822 1641 4248
rect 1646 4192 1649 4258
rect 1678 4172 1681 4248
rect 1686 4192 1689 4278
rect 1702 4272 1705 4428
rect 1710 4282 1713 4478
rect 1718 4352 1721 4418
rect 1726 4412 1729 4548
rect 1742 4482 1745 4518
rect 1750 4512 1753 4628
rect 1758 4542 1761 4598
rect 1774 4562 1777 4638
rect 1770 4558 1774 4561
rect 1742 4462 1745 4478
rect 1750 4372 1753 4508
rect 1766 4362 1769 4518
rect 1774 4472 1777 4538
rect 1782 4522 1785 4558
rect 1782 4472 1785 4488
rect 1790 4462 1793 4538
rect 1806 4532 1809 4538
rect 1806 4518 1814 4521
rect 1806 4482 1809 4518
rect 1862 4512 1865 4548
rect 1878 4542 1881 4638
rect 1838 4492 1841 4508
rect 1872 4503 1874 4507
rect 1878 4503 1881 4507
rect 1885 4503 1888 4507
rect 1894 4502 1897 4618
rect 1918 4542 1921 4668
rect 1846 4462 1849 4468
rect 1854 4462 1857 4478
rect 1910 4472 1913 4538
rect 1918 4482 1921 4538
rect 1826 4458 1830 4461
rect 1786 4448 1790 4451
rect 1798 4432 1801 4448
rect 1726 4352 1729 4358
rect 1698 4268 1702 4271
rect 1718 4271 1721 4318
rect 1710 4268 1721 4271
rect 1710 4262 1713 4268
rect 1726 4262 1729 4308
rect 1734 4272 1737 4328
rect 1742 4302 1745 4348
rect 1766 4342 1769 4348
rect 1750 4282 1753 4338
rect 1782 4322 1785 4347
rect 1758 4292 1761 4318
rect 1734 4252 1737 4268
rect 1742 4262 1745 4268
rect 1750 4262 1753 4278
rect 1766 4272 1769 4278
rect 1774 4262 1777 4298
rect 1766 4258 1774 4261
rect 1694 4242 1697 4248
rect 1758 4242 1761 4248
rect 1726 4192 1729 4218
rect 1654 4142 1657 4158
rect 1654 4072 1657 4138
rect 1662 4052 1665 4058
rect 1670 4042 1673 4158
rect 1686 4032 1689 4148
rect 1694 4142 1697 4188
rect 1734 4152 1737 4158
rect 1694 4132 1697 4138
rect 1710 4082 1713 4088
rect 1722 4078 1726 4081
rect 1734 4072 1737 4098
rect 1742 4092 1745 4208
rect 1766 4202 1769 4258
rect 1786 4248 1790 4251
rect 1774 4242 1777 4248
rect 1758 4142 1761 4148
rect 1758 4082 1761 4088
rect 1746 4078 1750 4081
rect 1774 4062 1777 4078
rect 1782 4072 1785 4188
rect 1798 4182 1801 4248
rect 1798 4062 1801 4148
rect 1806 4071 1809 4458
rect 1814 4322 1817 4338
rect 1846 4312 1849 4318
rect 1814 4262 1817 4308
rect 1854 4292 1857 4358
rect 1870 4352 1873 4458
rect 1910 4392 1913 4458
rect 1926 4382 1929 4548
rect 1934 4542 1937 4948
rect 1942 4742 1945 4748
rect 1950 4702 1953 4938
rect 1958 4932 1961 5018
rect 1966 5002 1969 5058
rect 1982 4942 1985 5058
rect 2086 5032 2089 5059
rect 2150 5052 2153 5058
rect 2342 5042 2345 5058
rect 2026 5018 2030 5021
rect 2014 4952 2017 5018
rect 2134 4992 2137 4998
rect 1998 4892 2001 4947
rect 2030 4882 2033 4918
rect 1982 4862 1985 4878
rect 2046 4872 2049 4968
rect 2074 4958 2078 4961
rect 2150 4952 2153 4958
rect 2190 4952 2193 5038
rect 2206 4992 2209 5018
rect 2218 4958 2222 4961
rect 2198 4952 2201 4958
rect 2130 4948 2134 4951
rect 2070 4932 2073 4948
rect 2086 4922 2089 4948
rect 2094 4922 2097 4938
rect 2158 4932 2161 4948
rect 2058 4918 2062 4921
rect 2102 4912 2105 4918
rect 1990 4862 1993 4868
rect 2018 4858 2022 4861
rect 1966 4772 1969 4818
rect 2046 4762 2049 4868
rect 2070 4862 2073 4868
rect 2102 4762 2105 4768
rect 2110 4762 2113 4928
rect 2166 4872 2169 4878
rect 2146 4858 2150 4861
rect 2158 4852 2161 4858
rect 2142 4822 2145 4848
rect 1966 4752 1969 4758
rect 2046 4752 2049 4758
rect 2118 4752 2121 4778
rect 2070 4742 2073 4747
rect 2126 4742 2129 4788
rect 2134 4742 2137 4758
rect 2142 4752 2145 4818
rect 2174 4802 2177 4948
rect 2182 4862 2185 4948
rect 2190 4932 2193 4938
rect 2206 4932 2209 4948
rect 2238 4942 2241 4948
rect 2222 4932 2225 4938
rect 2182 4802 2185 4858
rect 2158 4762 2161 4778
rect 2162 4748 2166 4751
rect 1990 4718 1998 4721
rect 1990 4682 1993 4718
rect 2006 4712 2009 4718
rect 2022 4692 2025 4738
rect 2078 4672 2081 4698
rect 1994 4668 1998 4671
rect 2058 4668 2062 4671
rect 2014 4662 2017 4668
rect 2086 4662 2089 4678
rect 2006 4652 2009 4658
rect 1974 4612 1977 4618
rect 1950 4552 1953 4558
rect 1958 4542 1961 4548
rect 1938 4538 1942 4541
rect 1958 4418 1966 4421
rect 1958 4372 1961 4418
rect 1894 4352 1897 4368
rect 1942 4362 1945 4368
rect 1930 4358 1934 4361
rect 1862 4342 1865 4348
rect 1878 4332 1881 4338
rect 1872 4303 1874 4307
rect 1878 4303 1881 4307
rect 1885 4303 1888 4307
rect 1902 4282 1905 4318
rect 1822 4272 1825 4278
rect 1814 4252 1817 4258
rect 1814 4222 1817 4228
rect 1814 4192 1817 4198
rect 1822 4132 1825 4268
rect 1830 4262 1833 4268
rect 1918 4262 1921 4298
rect 1838 4252 1841 4258
rect 1926 4252 1929 4348
rect 1934 4262 1937 4338
rect 1838 4192 1841 4248
rect 1830 4162 1833 4168
rect 1822 4122 1825 4128
rect 1830 4112 1833 4118
rect 1846 4092 1849 4148
rect 1854 4142 1857 4148
rect 1806 4068 1814 4071
rect 1722 4058 1726 4061
rect 1826 4058 1830 4061
rect 1702 3992 1705 4058
rect 1750 3982 1753 4058
rect 1790 4052 1793 4058
rect 1806 4042 1809 4058
rect 1826 4048 1830 4051
rect 1658 3968 1662 3971
rect 1694 3962 1697 3968
rect 1646 3852 1649 3868
rect 1654 3862 1657 3958
rect 1666 3948 1670 3951
rect 1682 3938 1686 3941
rect 1662 3932 1665 3938
rect 1670 3892 1673 3928
rect 1662 3872 1665 3878
rect 1678 3832 1681 3858
rect 1474 3748 1478 3751
rect 1518 3751 1521 3768
rect 1434 3738 1441 3741
rect 1486 3732 1489 3738
rect 1406 3662 1409 3668
rect 1430 3662 1433 3678
rect 1478 3672 1481 3678
rect 1374 3652 1377 3659
rect 1352 3603 1354 3607
rect 1358 3603 1361 3607
rect 1365 3603 1368 3607
rect 1338 3588 1342 3591
rect 1214 3572 1217 3588
rect 1190 3562 1193 3568
rect 1026 3538 1030 3541
rect 1174 3532 1177 3538
rect 1038 3522 1041 3528
rect 1070 3492 1073 3498
rect 1190 3492 1193 3548
rect 1066 3488 1070 3491
rect 942 3452 945 3488
rect 1094 3482 1097 3488
rect 966 3462 969 3478
rect 1202 3468 1206 3471
rect 954 3458 958 3461
rect 974 3451 977 3468
rect 966 3448 977 3451
rect 942 3392 945 3438
rect 950 3348 958 3351
rect 950 3262 953 3348
rect 966 3342 969 3448
rect 974 3352 977 3398
rect 990 3371 993 3468
rect 1006 3452 1009 3459
rect 1038 3372 1041 3458
rect 1078 3442 1081 3458
rect 1094 3402 1097 3418
rect 1118 3392 1121 3468
rect 1214 3462 1217 3558
rect 1230 3552 1233 3558
rect 1342 3552 1345 3578
rect 1238 3542 1241 3548
rect 1270 3481 1273 3538
rect 1278 3512 1281 3538
rect 1286 3522 1289 3548
rect 1346 3538 1350 3541
rect 1390 3532 1393 3558
rect 1294 3492 1297 3528
rect 1366 3512 1369 3518
rect 1262 3478 1273 3481
rect 1238 3462 1241 3468
rect 1254 3462 1257 3478
rect 1262 3472 1265 3478
rect 1310 3472 1313 3508
rect 1274 3468 1278 3471
rect 1146 3458 1150 3461
rect 1282 3458 1286 3461
rect 1234 3448 1238 3451
rect 1198 3442 1201 3448
rect 1254 3422 1257 3458
rect 1290 3448 1294 3451
rect 1310 3392 1313 3468
rect 1334 3462 1337 3508
rect 1390 3492 1393 3528
rect 1406 3472 1409 3658
rect 1414 3542 1417 3618
rect 1422 3562 1425 3658
rect 1422 3552 1425 3558
rect 1430 3552 1433 3658
rect 1438 3652 1441 3658
rect 1454 3652 1457 3668
rect 1474 3658 1478 3661
rect 1486 3642 1489 3698
rect 1502 3692 1505 3738
rect 1506 3668 1510 3671
rect 1542 3662 1545 3798
rect 1578 3788 1582 3791
rect 1614 3752 1617 3758
rect 1646 3752 1649 3808
rect 1602 3748 1606 3751
rect 1670 3742 1673 3748
rect 1642 3738 1646 3741
rect 1634 3728 1638 3731
rect 1650 3728 1654 3731
rect 1550 3722 1553 3728
rect 1550 3692 1553 3718
rect 1662 3701 1665 3718
rect 1654 3698 1665 3701
rect 1566 3672 1569 3678
rect 1578 3668 1582 3671
rect 1506 3658 1510 3661
rect 1578 3658 1582 3661
rect 1598 3652 1601 3688
rect 1618 3658 1622 3661
rect 1550 3642 1553 3648
rect 1582 3642 1585 3648
rect 1606 3642 1609 3648
rect 1622 3642 1625 3648
rect 1462 3592 1465 3608
rect 1486 3602 1489 3638
rect 1446 3562 1449 3568
rect 1414 3492 1417 3538
rect 1352 3403 1354 3407
rect 1358 3403 1361 3407
rect 1365 3403 1368 3407
rect 1422 3402 1425 3538
rect 1430 3512 1433 3548
rect 1454 3532 1457 3558
rect 1470 3542 1473 3588
rect 1478 3552 1481 3558
rect 1494 3542 1497 3638
rect 1630 3632 1633 3668
rect 1654 3662 1657 3698
rect 1666 3688 1670 3691
rect 1638 3642 1641 3648
rect 1654 3632 1657 3638
rect 1662 3632 1665 3668
rect 1678 3661 1681 3748
rect 1686 3702 1689 3868
rect 1694 3862 1697 3958
rect 1702 3892 1705 3968
rect 1750 3952 1753 3978
rect 1774 3972 1777 4018
rect 1806 4002 1809 4018
rect 1790 3952 1793 3958
rect 1762 3948 1766 3951
rect 1754 3938 1758 3941
rect 1798 3941 1801 3948
rect 1786 3938 1801 3941
rect 1806 3942 1809 3948
rect 1718 3922 1721 3938
rect 1718 3902 1721 3918
rect 1734 3912 1737 3918
rect 1710 3862 1713 3878
rect 1750 3862 1753 3898
rect 1790 3892 1793 3928
rect 1806 3912 1809 3938
rect 1814 3932 1817 3938
rect 1822 3902 1825 3918
rect 1830 3892 1833 4008
rect 1838 3892 1841 4078
rect 1862 4071 1865 4238
rect 1926 4222 1929 4248
rect 1958 4242 1961 4328
rect 1974 4312 1977 4528
rect 2014 4492 2017 4658
rect 2038 4632 2041 4658
rect 2050 4648 2054 4651
rect 2070 4632 2073 4658
rect 2094 4642 2097 4668
rect 2094 4592 2097 4638
rect 2038 4552 2041 4558
rect 2102 4502 2105 4718
rect 2118 4682 2121 4708
rect 2150 4692 2153 4738
rect 2110 4672 2113 4678
rect 2110 4562 2113 4618
rect 2134 4552 2137 4558
rect 2110 4532 2113 4548
rect 2022 4472 2025 4498
rect 2070 4472 2073 4488
rect 2106 4468 2110 4471
rect 1998 4452 2001 4458
rect 2018 4448 2022 4451
rect 2034 4448 2038 4451
rect 1990 4351 1993 4358
rect 1990 4322 1993 4328
rect 1998 4312 2001 4418
rect 2046 4322 2049 4468
rect 2078 4462 2081 4468
rect 2118 4462 2121 4548
rect 2158 4492 2161 4718
rect 2174 4711 2177 4798
rect 2190 4792 2193 4858
rect 2206 4812 2209 4928
rect 2238 4872 2241 4938
rect 2254 4932 2257 4947
rect 2262 4932 2265 5018
rect 2302 4872 2305 5008
rect 2350 4992 2353 5048
rect 2446 5022 2449 5058
rect 2454 5052 2457 5078
rect 3566 5072 3569 5078
rect 5014 5072 5017 5078
rect 5022 5072 5025 5078
rect 2506 5068 2510 5071
rect 2746 5068 2750 5071
rect 3074 5068 3078 5071
rect 3114 5068 3118 5071
rect 3186 5068 3190 5071
rect 3922 5068 3926 5071
rect 3962 5068 3966 5071
rect 4034 5068 4038 5071
rect 4858 5068 4862 5071
rect 5050 5068 5054 5071
rect 5234 5068 5238 5071
rect 2402 5018 2406 5021
rect 2384 5003 2386 5007
rect 2390 5003 2393 5007
rect 2397 5003 2400 5007
rect 2318 4952 2321 4968
rect 2390 4952 2393 4988
rect 2354 4948 2358 4951
rect 2326 4942 2329 4948
rect 2334 4942 2337 4948
rect 2326 4882 2329 4938
rect 2222 4852 2225 4859
rect 2326 4852 2329 4858
rect 2182 4732 2185 4738
rect 2166 4708 2177 4711
rect 2166 4662 2169 4708
rect 2190 4672 2193 4768
rect 2214 4752 2217 4778
rect 2222 4752 2225 4798
rect 2254 4762 2257 4768
rect 2274 4748 2278 4751
rect 2206 4742 2209 4748
rect 2286 4741 2289 4818
rect 2334 4812 2337 4938
rect 2390 4932 2393 4948
rect 2406 4942 2409 4978
rect 2418 4958 2422 4961
rect 2406 4922 2409 4938
rect 2430 4932 2433 5018
rect 2454 4992 2457 5038
rect 2478 5002 2481 5058
rect 2486 5042 2489 5068
rect 2542 5062 2545 5068
rect 2558 5063 2561 5068
rect 2638 5062 2641 5068
rect 2662 5062 2665 5068
rect 2478 4952 2481 4998
rect 2442 4948 2446 4951
rect 2490 4948 2494 4951
rect 2470 4942 2473 4948
rect 2422 4922 2425 4928
rect 2414 4882 2417 4888
rect 2294 4752 2297 4758
rect 2350 4752 2353 4858
rect 2384 4803 2386 4807
rect 2390 4803 2393 4807
rect 2397 4803 2400 4807
rect 2414 4752 2417 4808
rect 2422 4762 2425 4918
rect 2430 4872 2433 4928
rect 2454 4862 2457 4878
rect 2478 4862 2481 4948
rect 2486 4932 2489 4938
rect 2502 4901 2505 5058
rect 2510 5042 2513 5058
rect 2518 4992 2521 5028
rect 2558 4952 2561 4978
rect 2570 4958 2574 4961
rect 2582 4952 2585 4968
rect 2614 4952 2617 5048
rect 2742 5042 2745 5058
rect 2766 5042 2769 5068
rect 2790 5062 2793 5068
rect 2894 5062 2897 5068
rect 3022 5063 3025 5068
rect 2818 5058 2822 5061
rect 2774 5052 2777 5058
rect 2722 5018 2726 5021
rect 2626 4958 2630 4961
rect 2638 4952 2641 5018
rect 2790 4982 2793 5058
rect 2662 4962 2665 4968
rect 2494 4898 2505 4901
rect 2530 4948 2534 4951
rect 2562 4948 2566 4951
rect 2642 4948 2646 4951
rect 2694 4951 2697 4958
rect 2510 4942 2513 4948
rect 2542 4942 2545 4948
rect 2550 4942 2553 4948
rect 2790 4942 2793 4978
rect 2858 4968 2862 4971
rect 2866 4948 2870 4951
rect 2642 4938 2646 4941
rect 2494 4882 2497 4898
rect 2502 4862 2505 4868
rect 2434 4858 2438 4861
rect 2430 4782 2433 4858
rect 2438 4842 2441 4848
rect 2462 4792 2465 4858
rect 2510 4812 2513 4938
rect 2542 4852 2545 4938
rect 2598 4922 2601 4928
rect 2574 4892 2577 4918
rect 2558 4882 2561 4888
rect 2570 4878 2574 4881
rect 2590 4872 2593 4918
rect 2630 4902 2633 4918
rect 2582 4862 2585 4868
rect 2610 4858 2614 4861
rect 2638 4861 2641 4938
rect 2662 4892 2665 4928
rect 2670 4882 2673 4918
rect 2650 4878 2654 4881
rect 2638 4858 2646 4861
rect 2282 4738 2289 4741
rect 2166 4642 2169 4658
rect 2174 4622 2177 4658
rect 2190 4562 2193 4668
rect 2206 4662 2209 4738
rect 2278 4732 2281 4738
rect 2334 4722 2337 4748
rect 2214 4662 2217 4668
rect 2230 4582 2233 4718
rect 2286 4702 2289 4718
rect 2270 4682 2273 4688
rect 2310 4682 2313 4688
rect 2358 4682 2361 4738
rect 2390 4712 2393 4718
rect 2294 4672 2297 4678
rect 2278 4642 2281 4658
rect 2286 4652 2289 4668
rect 2326 4652 2329 4658
rect 2194 4558 2201 4561
rect 2190 4542 2193 4548
rect 2066 4458 2070 4461
rect 2090 4458 2094 4461
rect 2130 4458 2134 4461
rect 2054 4322 2057 4328
rect 1990 4262 1993 4308
rect 2022 4292 2025 4298
rect 1970 4248 1974 4251
rect 1998 4242 2001 4268
rect 2014 4262 2017 4268
rect 2038 4262 2041 4298
rect 2062 4292 2065 4298
rect 1878 4152 1881 4188
rect 1886 4162 1889 4168
rect 1934 4162 1937 4168
rect 1894 4158 1902 4161
rect 1874 4138 1878 4141
rect 1872 4103 1874 4107
rect 1878 4103 1881 4107
rect 1885 4103 1888 4107
rect 1894 4081 1897 4158
rect 1902 4152 1905 4158
rect 1930 4148 1934 4151
rect 1906 4138 1910 4141
rect 1902 4092 1905 4118
rect 1918 4112 1921 4148
rect 1950 4142 1953 4238
rect 1970 4228 1974 4231
rect 1990 4212 1993 4218
rect 1998 4202 2001 4238
rect 2046 4202 2049 4258
rect 2054 4232 2057 4278
rect 2070 4262 2073 4368
rect 2086 4292 2089 4358
rect 2110 4352 2113 4398
rect 2098 4348 2102 4351
rect 2118 4292 2121 4458
rect 2158 4402 2161 4438
rect 2154 4358 2158 4361
rect 2174 4352 2177 4528
rect 2198 4472 2201 4558
rect 2218 4548 2222 4551
rect 2206 4522 2209 4528
rect 2190 4462 2193 4468
rect 2222 4462 2225 4538
rect 2262 4532 2265 4548
rect 2238 4472 2241 4478
rect 2182 4342 2185 4368
rect 2198 4352 2201 4418
rect 2270 4411 2273 4618
rect 2278 4422 2281 4638
rect 2326 4572 2329 4648
rect 2366 4642 2369 4658
rect 2384 4603 2386 4607
rect 2390 4603 2393 4607
rect 2397 4603 2400 4607
rect 2394 4558 2398 4561
rect 2358 4552 2361 4558
rect 2286 4542 2289 4548
rect 2310 4518 2318 4521
rect 2310 4482 2313 4518
rect 2302 4452 2305 4458
rect 2270 4408 2281 4411
rect 2222 4352 2225 4358
rect 2238 4352 2241 4358
rect 2190 4342 2193 4348
rect 2150 4322 2153 4328
rect 2090 4278 2094 4281
rect 2030 4162 2033 4168
rect 2054 4152 2057 4218
rect 2094 4192 2097 4278
rect 2142 4272 2145 4278
rect 2142 4262 2145 4268
rect 2130 4258 2134 4261
rect 2102 4252 2105 4258
rect 2078 4162 2081 4168
rect 2070 4152 2073 4158
rect 1966 4142 1969 4147
rect 2046 4132 2049 4138
rect 1890 4078 1897 4081
rect 1858 4068 1865 4071
rect 1934 4072 1937 4078
rect 1950 4072 1953 4078
rect 1962 4058 1966 4061
rect 1846 4002 1849 4058
rect 1854 4012 1857 4058
rect 1918 4052 1921 4058
rect 1862 4042 1865 4048
rect 1874 3948 1878 3951
rect 1902 3942 1905 3948
rect 1778 3878 1782 3881
rect 1814 3872 1817 3878
rect 1822 3868 1830 3871
rect 1758 3862 1761 3868
rect 1822 3862 1825 3868
rect 1722 3858 1726 3861
rect 1810 3858 1814 3861
rect 1834 3848 1838 3851
rect 1694 3792 1697 3798
rect 1702 3782 1705 3848
rect 1710 3748 1718 3751
rect 1726 3751 1729 3818
rect 1766 3812 1769 3818
rect 1790 3792 1793 3818
rect 1750 3752 1753 3768
rect 1726 3748 1734 3751
rect 1710 3712 1713 3748
rect 1670 3658 1681 3661
rect 1718 3682 1721 3738
rect 1742 3732 1745 3738
rect 1730 3728 1734 3731
rect 1766 3682 1769 3728
rect 1502 3572 1505 3618
rect 1630 3602 1633 3628
rect 1662 3592 1665 3628
rect 1526 3552 1529 3558
rect 1506 3548 1510 3551
rect 1582 3551 1585 3558
rect 1622 3552 1625 3568
rect 1670 3562 1673 3658
rect 1654 3552 1657 3558
rect 1582 3548 1590 3551
rect 1610 3548 1614 3551
rect 1642 3548 1649 3551
rect 1534 3542 1537 3548
rect 1482 3538 1486 3541
rect 1450 3518 1454 3521
rect 1470 3492 1473 3538
rect 990 3368 1001 3371
rect 966 3312 969 3338
rect 750 3162 753 3218
rect 762 3158 766 3161
rect 774 3152 777 3178
rect 786 3158 790 3161
rect 838 3152 841 3228
rect 870 3212 873 3218
rect 870 3162 873 3178
rect 870 3152 873 3158
rect 878 3152 881 3218
rect 902 3202 905 3218
rect 886 3162 889 3178
rect 918 3162 921 3218
rect 934 3212 937 3218
rect 934 3162 937 3208
rect 950 3202 953 3258
rect 786 3148 790 3151
rect 898 3148 902 3151
rect 914 3148 918 3151
rect 646 3122 649 3138
rect 630 3082 633 3088
rect 662 3082 665 3118
rect 678 3082 681 3098
rect 678 3072 681 3078
rect 658 3068 662 3071
rect 646 3052 649 3058
rect 602 2968 606 2971
rect 606 2952 609 2958
rect 614 2942 617 3018
rect 662 3002 665 3058
rect 694 3052 697 3059
rect 726 3021 729 3118
rect 754 3088 758 3091
rect 766 3062 769 3108
rect 774 3092 777 3138
rect 798 3122 801 3148
rect 822 3142 825 3148
rect 814 3132 817 3138
rect 774 3062 777 3068
rect 726 3018 737 3021
rect 754 3018 758 3021
rect 734 2992 737 3018
rect 766 3012 769 3058
rect 774 2992 777 3058
rect 782 2992 785 3118
rect 802 3068 809 3071
rect 806 3062 809 3068
rect 794 3058 798 3061
rect 814 3042 817 3078
rect 734 2982 737 2988
rect 638 2942 641 2948
rect 618 2938 622 2941
rect 626 2928 630 2931
rect 590 2872 593 2888
rect 638 2882 641 2938
rect 654 2932 657 2968
rect 678 2942 681 2948
rect 686 2932 689 2948
rect 694 2922 697 2938
rect 710 2932 713 2958
rect 718 2942 721 2948
rect 670 2902 673 2918
rect 646 2892 649 2898
rect 662 2882 665 2888
rect 686 2882 689 2918
rect 622 2872 625 2878
rect 638 2872 641 2878
rect 562 2858 569 2861
rect 494 2792 497 2818
rect 502 2782 505 2848
rect 510 2762 513 2768
rect 526 2752 529 2858
rect 534 2852 537 2858
rect 546 2838 550 2841
rect 558 2802 561 2848
rect 566 2832 569 2858
rect 598 2842 601 2858
rect 614 2842 617 2858
rect 630 2852 633 2858
rect 574 2772 577 2788
rect 614 2782 617 2818
rect 414 2651 417 2738
rect 430 2702 433 2738
rect 454 2732 457 2748
rect 518 2742 521 2748
rect 526 2742 529 2748
rect 478 2692 481 2738
rect 550 2732 553 2758
rect 566 2752 569 2758
rect 582 2752 585 2778
rect 630 2752 633 2798
rect 638 2752 641 2808
rect 650 2758 654 2761
rect 662 2752 665 2868
rect 678 2862 681 2878
rect 686 2752 689 2818
rect 694 2812 697 2918
rect 702 2892 705 2918
rect 718 2862 721 2898
rect 742 2881 745 2988
rect 750 2952 753 2988
rect 758 2962 761 2968
rect 802 2948 806 2951
rect 750 2922 753 2948
rect 766 2922 769 2928
rect 814 2912 817 2938
rect 742 2878 753 2881
rect 738 2868 742 2871
rect 750 2862 753 2878
rect 782 2872 785 2908
rect 702 2812 705 2858
rect 738 2848 742 2851
rect 710 2792 713 2838
rect 718 2792 721 2818
rect 694 2762 697 2788
rect 750 2761 753 2818
rect 766 2812 769 2848
rect 750 2758 761 2761
rect 594 2748 598 2751
rect 714 2748 721 2751
rect 622 2742 625 2748
rect 726 2742 729 2758
rect 738 2748 742 2751
rect 538 2728 542 2731
rect 598 2712 601 2738
rect 718 2732 721 2738
rect 742 2732 745 2738
rect 634 2728 638 2731
rect 606 2702 609 2728
rect 614 2702 617 2718
rect 590 2692 593 2698
rect 554 2688 558 2691
rect 478 2682 481 2688
rect 582 2682 585 2688
rect 638 2682 641 2688
rect 422 2672 425 2678
rect 430 2662 433 2678
rect 594 2668 598 2671
rect 442 2658 446 2661
rect 574 2662 577 2668
rect 646 2662 649 2668
rect 430 2652 433 2658
rect 478 2652 481 2659
rect 414 2648 425 2651
rect 554 2648 558 2651
rect 410 2638 414 2641
rect 354 2568 358 2571
rect 326 2542 329 2568
rect 370 2558 374 2561
rect 382 2552 385 2638
rect 374 2542 377 2548
rect 390 2542 393 2618
rect 422 2612 425 2648
rect 446 2642 449 2648
rect 566 2642 569 2658
rect 606 2652 609 2658
rect 546 2638 550 2641
rect 410 2548 414 2551
rect 330 2538 337 2541
rect 354 2538 358 2541
rect 322 2528 326 2531
rect 306 2468 310 2471
rect 222 2462 225 2468
rect 318 2462 321 2518
rect 334 2482 337 2538
rect 410 2528 414 2531
rect 334 2462 337 2478
rect 350 2472 353 2488
rect 398 2482 401 2508
rect 290 2458 294 2461
rect 182 2352 185 2458
rect 186 2348 193 2351
rect 158 2338 169 2341
rect 126 2272 129 2278
rect 118 2262 121 2268
rect 150 2262 153 2268
rect 158 2262 161 2338
rect 170 2328 174 2331
rect 166 2262 169 2288
rect 182 2282 185 2318
rect 130 2258 134 2261
rect 62 2192 65 2258
rect 174 2172 177 2268
rect 190 2262 193 2348
rect 222 2351 225 2358
rect 206 2321 209 2348
rect 198 2318 209 2321
rect 198 2292 201 2318
rect 206 2272 209 2288
rect 218 2268 222 2271
rect 194 2258 201 2261
rect 170 2168 174 2171
rect 150 2162 153 2168
rect 114 2148 118 2151
rect 6 2072 9 2138
rect 86 2072 89 2138
rect 174 2132 177 2148
rect 182 2142 185 2178
rect 190 2142 193 2148
rect 6 1942 9 2068
rect 70 2062 73 2068
rect 86 2062 89 2068
rect 114 2058 118 2061
rect 62 1982 65 1988
rect 10 1938 14 1941
rect 6 1892 9 1898
rect 14 1742 17 1938
rect 70 1882 73 2058
rect 86 1942 89 2058
rect 166 1992 169 2078
rect 190 2062 193 2068
rect 198 2062 201 2258
rect 206 2182 209 2268
rect 230 2262 233 2418
rect 238 2332 241 2338
rect 218 2258 222 2261
rect 206 2132 209 2168
rect 222 2152 225 2178
rect 238 2162 241 2328
rect 246 2292 249 2428
rect 278 2412 281 2418
rect 318 2412 321 2448
rect 390 2442 393 2458
rect 414 2452 417 2528
rect 422 2502 425 2608
rect 486 2592 489 2638
rect 438 2542 441 2548
rect 446 2542 449 2568
rect 466 2558 470 2561
rect 438 2502 441 2528
rect 454 2511 457 2548
rect 470 2532 473 2558
rect 486 2552 489 2578
rect 502 2562 505 2638
rect 490 2548 497 2551
rect 482 2538 486 2541
rect 466 2518 470 2521
rect 454 2508 465 2511
rect 328 2403 330 2407
rect 334 2403 337 2407
rect 341 2403 344 2407
rect 318 2352 321 2358
rect 306 2338 310 2341
rect 350 2332 353 2338
rect 282 2318 286 2321
rect 270 2292 273 2308
rect 286 2302 289 2318
rect 294 2312 297 2328
rect 302 2291 305 2318
rect 302 2288 313 2291
rect 282 2278 286 2281
rect 262 2272 265 2278
rect 302 2272 305 2278
rect 290 2268 294 2271
rect 310 2262 313 2288
rect 374 2262 377 2378
rect 414 2362 417 2448
rect 394 2348 401 2351
rect 398 2292 401 2348
rect 422 2312 425 2458
rect 442 2448 446 2451
rect 446 2412 449 2448
rect 454 2432 457 2458
rect 462 2422 465 2508
rect 470 2492 473 2498
rect 478 2492 481 2538
rect 470 2382 473 2448
rect 478 2442 481 2458
rect 462 2352 465 2358
rect 438 2342 441 2348
rect 454 2342 457 2348
rect 446 2292 449 2318
rect 390 2272 393 2288
rect 406 2282 409 2288
rect 394 2268 398 2271
rect 426 2268 430 2271
rect 446 2262 449 2268
rect 250 2258 254 2261
rect 290 2258 294 2261
rect 362 2258 366 2261
rect 418 2258 422 2261
rect 454 2261 457 2338
rect 470 2312 473 2338
rect 478 2332 481 2438
rect 486 2332 489 2518
rect 494 2492 497 2548
rect 534 2511 537 2547
rect 566 2542 569 2598
rect 550 2532 553 2538
rect 526 2508 537 2511
rect 526 2492 529 2508
rect 494 2472 497 2488
rect 518 2462 521 2468
rect 542 2462 545 2508
rect 558 2472 561 2478
rect 566 2472 569 2538
rect 598 2482 601 2518
rect 606 2482 609 2488
rect 594 2478 598 2481
rect 614 2472 617 2608
rect 630 2511 633 2528
rect 622 2508 633 2511
rect 574 2462 577 2468
rect 610 2458 614 2461
rect 510 2452 513 2458
rect 506 2368 510 2371
rect 526 2352 529 2448
rect 542 2362 545 2368
rect 574 2362 577 2418
rect 590 2392 593 2438
rect 622 2372 625 2508
rect 646 2492 649 2548
rect 650 2468 654 2471
rect 662 2462 665 2658
rect 670 2622 673 2718
rect 750 2692 753 2748
rect 758 2742 761 2758
rect 798 2742 801 2868
rect 806 2862 809 2888
rect 810 2748 814 2751
rect 790 2712 793 2728
rect 714 2668 718 2671
rect 726 2662 729 2668
rect 706 2638 710 2641
rect 718 2632 721 2658
rect 734 2652 737 2668
rect 742 2642 745 2678
rect 758 2672 761 2678
rect 762 2658 766 2661
rect 766 2642 769 2648
rect 774 2591 777 2698
rect 790 2672 793 2708
rect 798 2682 801 2718
rect 822 2692 825 2798
rect 830 2792 833 3148
rect 838 3112 841 3148
rect 950 3142 953 3147
rect 850 3138 854 3141
rect 894 3132 897 3138
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 861 3103 864 3107
rect 958 3082 961 3138
rect 966 3132 969 3308
rect 982 3282 985 3368
rect 990 3352 993 3358
rect 998 3342 1001 3368
rect 1010 3358 1014 3361
rect 990 3332 993 3338
rect 994 3258 998 3261
rect 1006 3212 1009 3348
rect 1022 3342 1025 3358
rect 1038 3342 1041 3368
rect 1062 3332 1065 3348
rect 1078 3262 1081 3328
rect 1118 3322 1121 3338
rect 1126 3332 1129 3358
rect 1102 3262 1105 3268
rect 1090 3258 1094 3261
rect 1078 3252 1081 3258
rect 1126 3252 1129 3318
rect 1134 3262 1137 3378
rect 1142 3342 1145 3358
rect 1174 3342 1177 3368
rect 1198 3352 1201 3358
rect 1154 3338 1158 3341
rect 1146 3328 1150 3331
rect 1142 3262 1145 3278
rect 1150 3272 1153 3308
rect 1206 3282 1209 3388
rect 1254 3372 1257 3378
rect 1262 3342 1265 3378
rect 1294 3362 1297 3368
rect 1274 3358 1278 3361
rect 1318 3352 1321 3368
rect 1098 3248 1102 3251
rect 1150 3241 1153 3268
rect 1166 3262 1169 3268
rect 1158 3252 1161 3258
rect 1174 3252 1177 3268
rect 1206 3252 1209 3259
rect 1150 3238 1161 3241
rect 1014 3132 1017 3178
rect 1022 3152 1025 3218
rect 1030 3142 1033 3148
rect 1054 3142 1057 3148
rect 1014 3122 1017 3128
rect 1022 3092 1025 3098
rect 1038 3082 1041 3118
rect 1062 3112 1065 3218
rect 1126 3172 1129 3218
rect 1134 3192 1137 3198
rect 1158 3192 1161 3238
rect 1182 3192 1185 3238
rect 1082 3148 1086 3151
rect 1078 3132 1081 3138
rect 1094 3132 1097 3168
rect 1154 3158 1158 3161
rect 1190 3152 1193 3158
rect 1206 3152 1209 3208
rect 1222 3172 1225 3178
rect 1262 3171 1265 3338
rect 1270 3312 1273 3348
rect 1326 3342 1329 3358
rect 1338 3340 1342 3343
rect 1382 3342 1385 3388
rect 1422 3382 1425 3398
rect 1446 3392 1449 3468
rect 1458 3458 1462 3461
rect 1446 3372 1449 3388
rect 1462 3362 1465 3368
rect 1318 3322 1321 3338
rect 1270 3242 1273 3308
rect 1338 3268 1342 3271
rect 1302 3262 1305 3268
rect 1270 3222 1273 3228
rect 1278 3202 1281 3258
rect 1326 3252 1329 3258
rect 1294 3242 1297 3248
rect 1310 3222 1313 3248
rect 1326 3232 1329 3248
rect 1366 3221 1369 3318
rect 1382 3282 1385 3338
rect 1406 3332 1409 3348
rect 1470 3342 1473 3468
rect 1486 3442 1489 3538
rect 1526 3528 1534 3531
rect 1494 3462 1497 3528
rect 1526 3492 1529 3528
rect 1538 3518 1542 3521
rect 1542 3492 1545 3508
rect 1506 3488 1510 3491
rect 1514 3468 1518 3471
rect 1550 3461 1553 3538
rect 1558 3522 1561 3548
rect 1566 3532 1569 3548
rect 1574 3532 1577 3548
rect 1598 3541 1601 3548
rect 1598 3538 1609 3541
rect 1590 3532 1593 3538
rect 1558 3472 1561 3508
rect 1550 3458 1561 3461
rect 1502 3412 1505 3418
rect 1494 3362 1497 3378
rect 1502 3352 1505 3358
rect 1478 3332 1481 3348
rect 1470 3321 1473 3328
rect 1486 3321 1489 3338
rect 1470 3318 1489 3321
rect 1510 3312 1513 3458
rect 1518 3442 1521 3448
rect 1534 3442 1537 3448
rect 1542 3432 1545 3448
rect 1522 3378 1526 3381
rect 1534 3372 1537 3418
rect 1550 3392 1553 3448
rect 1518 3352 1521 3368
rect 1526 3332 1529 3338
rect 1490 3288 1494 3291
rect 1390 3262 1393 3288
rect 1510 3282 1513 3308
rect 1526 3292 1529 3328
rect 1478 3272 1481 3278
rect 1542 3272 1545 3358
rect 1550 3352 1553 3368
rect 1558 3342 1561 3458
rect 1566 3452 1569 3468
rect 1574 3362 1577 3518
rect 1582 3472 1585 3518
rect 1606 3492 1609 3538
rect 1622 3512 1625 3538
rect 1630 3532 1633 3538
rect 1598 3482 1601 3488
rect 1654 3482 1657 3518
rect 1590 3472 1593 3478
rect 1670 3472 1673 3538
rect 1686 3532 1689 3598
rect 1698 3548 1702 3551
rect 1710 3492 1713 3498
rect 1718 3492 1721 3678
rect 1750 3672 1753 3678
rect 1782 3672 1785 3738
rect 1726 3652 1729 3658
rect 1790 3632 1793 3658
rect 1790 3592 1793 3618
rect 1766 3572 1769 3578
rect 1754 3568 1761 3571
rect 1758 3542 1761 3568
rect 1786 3558 1790 3561
rect 1770 3548 1774 3551
rect 1762 3538 1766 3541
rect 1750 3512 1753 3538
rect 1790 3532 1793 3538
rect 1758 3492 1761 3528
rect 1750 3472 1753 3488
rect 1774 3472 1777 3478
rect 1798 3472 1801 3848
rect 1854 3832 1857 3938
rect 1918 3922 1921 4028
rect 1926 3982 1929 4048
rect 1942 3992 1945 4058
rect 1950 3992 1953 4058
rect 1958 3952 1961 3978
rect 1946 3948 1950 3951
rect 1966 3942 1969 3988
rect 1934 3932 1937 3938
rect 1872 3903 1874 3907
rect 1878 3903 1881 3907
rect 1885 3903 1888 3907
rect 1886 3872 1889 3888
rect 1898 3868 1902 3871
rect 1874 3838 1878 3841
rect 1814 3751 1817 3768
rect 1830 3742 1833 3828
rect 1854 3772 1857 3778
rect 1886 3762 1889 3868
rect 1906 3858 1910 3861
rect 1910 3802 1913 3818
rect 1878 3752 1881 3758
rect 1846 3722 1849 3738
rect 1814 3672 1817 3688
rect 1834 3678 1838 3681
rect 1854 3662 1857 3748
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1885 3703 1888 3707
rect 1894 3672 1897 3698
rect 1910 3672 1913 3778
rect 1918 3742 1921 3918
rect 1930 3868 1934 3871
rect 1918 3682 1921 3688
rect 1926 3672 1929 3848
rect 1942 3822 1945 3858
rect 1954 3848 1958 3851
rect 1934 3752 1937 3758
rect 1942 3732 1945 3818
rect 1966 3812 1969 3868
rect 1950 3712 1953 3758
rect 1958 3752 1961 3758
rect 1974 3751 1977 4108
rect 1998 4062 2001 4088
rect 1986 4058 1990 4061
rect 1986 4038 1990 4041
rect 2006 3992 2009 4018
rect 2010 3958 2022 3961
rect 2010 3948 2014 3951
rect 2018 3938 2022 3941
rect 1986 3928 1990 3931
rect 1998 3872 2001 3878
rect 2030 3872 2033 4098
rect 2038 4082 2041 4118
rect 2054 4032 2057 4138
rect 2078 4132 2081 4158
rect 2086 4152 2089 4188
rect 2106 4158 2110 4161
rect 2142 4152 2145 4188
rect 2150 4152 2153 4308
rect 2158 4252 2161 4318
rect 2166 4262 2169 4328
rect 2230 4312 2233 4348
rect 2262 4342 2265 4398
rect 2238 4322 2241 4328
rect 2214 4272 2217 4278
rect 2222 4272 2225 4278
rect 2262 4272 2265 4338
rect 2174 4262 2177 4268
rect 2134 4142 2137 4148
rect 2114 4138 2118 4141
rect 2086 4122 2089 4138
rect 2114 4128 2118 4131
rect 2102 4072 2105 4078
rect 2126 4071 2129 4118
rect 2166 4102 2169 4258
rect 2190 4242 2193 4248
rect 2198 4231 2201 4258
rect 2254 4252 2257 4259
rect 2190 4228 2201 4231
rect 2206 4242 2209 4248
rect 2190 4212 2193 4228
rect 2198 4192 2201 4218
rect 2194 4168 2198 4171
rect 2178 4148 2182 4151
rect 2194 4148 2198 4151
rect 2206 4142 2209 4238
rect 2250 4148 2254 4151
rect 2262 4142 2265 4268
rect 2278 4252 2281 4408
rect 2326 4372 2329 4538
rect 2350 4532 2353 4548
rect 2334 4472 2337 4528
rect 2366 4482 2369 4538
rect 2374 4482 2377 4518
rect 2382 4492 2385 4528
rect 2402 4518 2406 4521
rect 2326 4362 2329 4368
rect 2286 4342 2289 4348
rect 2318 4282 2321 4288
rect 2334 4271 2337 4458
rect 2358 4422 2361 4458
rect 2366 4352 2369 4458
rect 2374 4382 2377 4478
rect 2382 4462 2385 4478
rect 2406 4462 2409 4468
rect 2386 4458 2390 4461
rect 2390 4442 2393 4458
rect 2414 4412 2417 4748
rect 2454 4742 2457 4748
rect 2478 4742 2481 4748
rect 2422 4732 2425 4738
rect 2430 4722 2433 4728
rect 2438 4722 2441 4728
rect 2426 4688 2430 4691
rect 2438 4682 2441 4708
rect 2454 4692 2457 4728
rect 2462 4682 2465 4688
rect 2462 4662 2465 4668
rect 2454 4552 2457 4558
rect 2470 4542 2473 4728
rect 2486 4662 2489 4668
rect 2478 4602 2481 4618
rect 2486 4552 2489 4658
rect 2494 4652 2497 4668
rect 2518 4662 2521 4848
rect 2538 4748 2542 4751
rect 2534 4722 2537 4728
rect 2538 4678 2542 4681
rect 2550 4671 2553 4748
rect 2558 4732 2561 4738
rect 2558 4682 2561 4688
rect 2542 4668 2553 4671
rect 2582 4672 2585 4738
rect 2590 4672 2593 4858
rect 2622 4852 2625 4858
rect 2630 4842 2633 4858
rect 2638 4762 2641 4818
rect 2610 4748 2614 4751
rect 2630 4742 2633 4748
rect 2638 4742 2641 4748
rect 2610 4738 2614 4741
rect 2602 4728 2606 4731
rect 2662 4712 2665 4718
rect 2654 4682 2657 4688
rect 2530 4658 2534 4661
rect 2518 4652 2521 4658
rect 2510 4582 2513 4618
rect 2518 4592 2521 4638
rect 2510 4552 2513 4568
rect 2534 4552 2537 4598
rect 2422 4432 2425 4468
rect 2384 4403 2386 4407
rect 2390 4403 2393 4407
rect 2397 4403 2400 4407
rect 2390 4352 2393 4378
rect 2414 4352 2417 4368
rect 2330 4268 2337 4271
rect 2334 4222 2337 4258
rect 2302 4182 2305 4188
rect 2342 4161 2345 4348
rect 2422 4342 2425 4348
rect 2370 4338 2374 4341
rect 2430 4332 2433 4388
rect 2438 4331 2441 4418
rect 2446 4392 2449 4448
rect 2454 4401 2457 4498
rect 2474 4468 2478 4471
rect 2462 4432 2465 4458
rect 2454 4398 2465 4401
rect 2446 4342 2449 4358
rect 2454 4352 2457 4378
rect 2462 4362 2465 4398
rect 2478 4372 2481 4418
rect 2494 4362 2497 4388
rect 2478 4352 2481 4358
rect 2502 4352 2505 4548
rect 2534 4472 2537 4548
rect 2526 4452 2529 4458
rect 2526 4352 2529 4448
rect 2542 4422 2545 4668
rect 2582 4662 2585 4668
rect 2590 4662 2593 4668
rect 2574 4652 2577 4658
rect 2574 4551 2577 4578
rect 2590 4562 2593 4618
rect 2558 4532 2561 4538
rect 2590 4462 2593 4558
rect 2606 4552 2609 4668
rect 2622 4652 2625 4659
rect 2638 4592 2641 4678
rect 2650 4668 2654 4671
rect 2670 4602 2673 4878
rect 2678 4832 2681 4868
rect 2702 4672 2705 4938
rect 2754 4918 2758 4921
rect 2774 4882 2777 4938
rect 2798 4932 2801 4948
rect 2874 4938 2878 4941
rect 2894 4932 2897 4968
rect 2878 4922 2881 4928
rect 2888 4903 2890 4907
rect 2894 4903 2897 4907
rect 2901 4903 2904 4907
rect 2854 4882 2857 4888
rect 2862 4862 2865 4868
rect 2786 4858 2790 4861
rect 2714 4748 2718 4751
rect 2742 4742 2745 4858
rect 2830 4772 2833 4788
rect 2894 4782 2897 4858
rect 2902 4852 2905 4858
rect 2878 4752 2881 4778
rect 2794 4748 2798 4751
rect 2854 4742 2857 4748
rect 2902 4742 2905 4748
rect 2870 4732 2873 4738
rect 2858 4728 2862 4731
rect 2898 4728 2902 4731
rect 2886 4722 2889 4728
rect 2846 4712 2849 4718
rect 2888 4703 2890 4707
rect 2894 4703 2897 4707
rect 2901 4703 2904 4707
rect 2910 4682 2913 4928
rect 2918 4882 2921 5058
rect 2942 5012 2945 5058
rect 2926 4952 2929 4968
rect 2926 4942 2929 4948
rect 2926 4822 2929 4858
rect 2934 4842 2937 4958
rect 2942 4952 2945 5008
rect 2942 4932 2945 4938
rect 2950 4842 2953 5058
rect 2962 5028 2966 5031
rect 2958 4952 2961 5018
rect 2958 4872 2961 4938
rect 2966 4932 2969 4938
rect 2966 4872 2969 4888
rect 2862 4672 2865 4678
rect 2702 4662 2705 4668
rect 2814 4662 2817 4668
rect 2870 4662 2873 4668
rect 2730 4658 2734 4661
rect 2918 4661 2921 4818
rect 2926 4752 2929 4758
rect 2958 4742 2961 4788
rect 2974 4732 2977 4918
rect 2982 4882 2985 4888
rect 2990 4872 2993 4948
rect 2986 4868 2990 4871
rect 2998 4862 3001 5028
rect 3038 5022 3041 5068
rect 3054 5052 3057 5068
rect 3066 5058 3070 5061
rect 3054 4982 3057 5048
rect 3086 5032 3089 5048
rect 3126 5042 3129 5048
rect 3006 4952 3009 4958
rect 3046 4952 3049 4978
rect 3110 4952 3113 4968
rect 3126 4962 3129 5038
rect 3118 4952 3121 4958
rect 3078 4942 3081 4947
rect 3110 4932 3113 4948
rect 3126 4932 3129 4938
rect 3142 4912 3145 5058
rect 3150 4992 3153 5068
rect 3158 5052 3161 5058
rect 3166 5042 3169 5058
rect 3174 5052 3177 5058
rect 3182 5042 3185 5048
rect 3198 5042 3201 5058
rect 3150 4952 3153 4978
rect 3018 4888 3022 4891
rect 3022 4872 3025 4878
rect 3070 4872 3073 4898
rect 3134 4882 3137 4888
rect 3030 4862 3033 4868
rect 3054 4852 3057 4868
rect 3118 4862 3121 4868
rect 3018 4848 3025 4851
rect 2982 4772 2985 4818
rect 2990 4742 2993 4748
rect 2934 4692 2937 4718
rect 2942 4692 2945 4728
rect 2982 4682 2985 4738
rect 3022 4712 3025 4848
rect 2930 4678 2934 4681
rect 2926 4662 2929 4668
rect 2918 4658 2926 4661
rect 2690 4618 2697 4621
rect 2678 4542 2681 4548
rect 2638 4512 2641 4518
rect 2614 4492 2617 4498
rect 2646 4482 2649 4518
rect 2686 4502 2689 4548
rect 2686 4462 2689 4478
rect 2550 4392 2553 4458
rect 2590 4441 2593 4458
rect 2598 4452 2601 4458
rect 2582 4438 2593 4441
rect 2538 4368 2545 4371
rect 2534 4352 2537 4368
rect 2514 4348 2518 4351
rect 2514 4338 2518 4341
rect 2438 4328 2449 4331
rect 2430 4282 2433 4328
rect 2350 4252 2353 4278
rect 2438 4272 2441 4318
rect 2446 4272 2449 4328
rect 2462 4302 2465 4318
rect 2486 4312 2489 4338
rect 2498 4318 2502 4321
rect 2462 4272 2465 4278
rect 2426 4268 2430 4271
rect 2490 4268 2494 4271
rect 2366 4262 2369 4268
rect 2438 4252 2441 4258
rect 2382 4242 2385 4248
rect 2384 4203 2386 4207
rect 2390 4203 2393 4207
rect 2397 4203 2400 4207
rect 2406 4172 2409 4218
rect 2342 4158 2353 4161
rect 2314 4148 2318 4151
rect 2338 4148 2345 4151
rect 2122 4068 2129 4071
rect 2086 4042 2089 4059
rect 2154 4058 2158 4061
rect 2174 4061 2177 4118
rect 2190 4062 2193 4138
rect 2230 4082 2233 4138
rect 2326 4132 2329 4148
rect 2342 4112 2345 4148
rect 2330 4078 2334 4081
rect 2230 4072 2233 4078
rect 2238 4062 2241 4078
rect 2342 4062 2345 4108
rect 2350 4072 2353 4158
rect 2454 4152 2457 4268
rect 2470 4262 2473 4268
rect 2510 4252 2513 4258
rect 2486 4242 2489 4248
rect 2470 4202 2473 4218
rect 2462 4152 2465 4178
rect 2510 4152 2513 4218
rect 2430 4142 2433 4147
rect 2362 4138 2366 4141
rect 2398 4122 2401 4128
rect 2490 4118 2494 4121
rect 2366 4102 2369 4108
rect 2366 4062 2369 4098
rect 2406 4072 2409 4078
rect 2174 4058 2182 4061
rect 2306 4058 2310 4061
rect 2418 4058 2422 4061
rect 2042 3958 2065 3961
rect 2042 3948 2046 3951
rect 2054 3942 2057 3948
rect 2062 3942 2065 3958
rect 2042 3938 2046 3941
rect 2078 3932 2081 3998
rect 2102 3992 2105 4038
rect 2094 3952 2097 3988
rect 2118 3962 2121 4008
rect 2126 3972 2129 4058
rect 2134 3972 2137 4058
rect 2142 4042 2145 4048
rect 2118 3952 2121 3958
rect 2126 3952 2129 3958
rect 2086 3932 2089 3948
rect 2070 3882 2073 3918
rect 2134 3882 2137 3958
rect 2166 3952 2169 3958
rect 2158 3942 2161 3948
rect 2102 3872 2105 3878
rect 2042 3868 2046 3871
rect 2086 3862 2089 3868
rect 2010 3858 2014 3861
rect 2042 3858 2046 3861
rect 2098 3858 2102 3861
rect 1990 3852 1993 3858
rect 2078 3852 2081 3858
rect 2110 3852 2113 3858
rect 2066 3848 2070 3851
rect 2126 3822 2129 3848
rect 2134 3821 2137 3878
rect 2150 3872 2153 3918
rect 2162 3888 2166 3891
rect 2150 3852 2153 3858
rect 2130 3818 2137 3821
rect 1990 3762 1993 3818
rect 2110 3812 2113 3818
rect 1970 3748 1977 3751
rect 1982 3752 1985 3758
rect 2030 3752 2033 3788
rect 2094 3752 2097 3798
rect 2126 3752 2129 3768
rect 2142 3752 2145 3818
rect 2154 3778 2158 3781
rect 2114 3748 2118 3751
rect 1962 3738 1966 3741
rect 1826 3648 1830 3651
rect 1838 3602 1841 3618
rect 1806 3512 1809 3548
rect 1814 3542 1817 3548
rect 1830 3512 1833 3538
rect 1586 3458 1590 3461
rect 1586 3448 1590 3451
rect 1582 3352 1585 3358
rect 1590 3352 1593 3408
rect 1598 3362 1601 3458
rect 1606 3372 1609 3378
rect 1558 3322 1561 3338
rect 1566 3312 1569 3328
rect 1450 3248 1454 3251
rect 1470 3242 1473 3248
rect 1478 3232 1481 3258
rect 1502 3252 1505 3258
rect 1486 3242 1489 3248
rect 1366 3218 1377 3221
rect 1254 3168 1265 3171
rect 1246 3152 1249 3158
rect 1238 3142 1241 3148
rect 1154 3138 1158 3141
rect 1178 3138 1182 3141
rect 1202 3138 1206 3141
rect 1102 3132 1105 3138
rect 1070 3102 1073 3128
rect 846 3072 849 3078
rect 942 3072 945 3078
rect 866 3059 870 3062
rect 966 3062 969 3078
rect 1038 3062 1041 3068
rect 1062 3062 1065 3068
rect 1142 3062 1145 3128
rect 1246 3122 1249 3148
rect 1254 3142 1257 3168
rect 1286 3142 1289 3147
rect 1254 3132 1257 3138
rect 1154 3068 1158 3071
rect 1174 3062 1177 3078
rect 1182 3062 1185 3068
rect 1130 3058 1134 3061
rect 1170 3058 1174 3061
rect 1006 3042 1009 3058
rect 1102 3042 1105 3048
rect 930 3038 934 3041
rect 926 2992 929 3008
rect 942 2952 945 2958
rect 1006 2952 1009 3038
rect 1070 2952 1073 2978
rect 1078 2972 1081 3028
rect 1142 3002 1145 3058
rect 1198 3052 1201 3068
rect 1226 3058 1230 3061
rect 1270 3052 1273 3138
rect 1310 3102 1313 3218
rect 1352 3203 1354 3207
rect 1358 3203 1361 3207
rect 1365 3203 1368 3207
rect 1346 3178 1350 3181
rect 1350 3142 1353 3178
rect 1374 3152 1377 3218
rect 1382 3172 1385 3178
rect 1390 3162 1393 3178
rect 1478 3172 1481 3228
rect 1414 3162 1417 3168
rect 1402 3158 1406 3161
rect 1434 3158 1438 3161
rect 1490 3158 1494 3161
rect 1278 3082 1281 3088
rect 1286 3082 1289 3098
rect 1374 3092 1377 3138
rect 1334 3072 1337 3078
rect 1326 3062 1329 3068
rect 1342 3062 1345 3068
rect 1158 2952 1161 2958
rect 858 2948 862 2951
rect 1146 2948 1150 2951
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 861 2903 864 2907
rect 870 2892 873 2918
rect 870 2862 873 2868
rect 850 2838 854 2841
rect 854 2762 857 2768
rect 862 2722 865 2818
rect 878 2752 881 2928
rect 902 2892 905 2948
rect 910 2902 913 2918
rect 894 2852 897 2868
rect 918 2852 921 2858
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 861 2703 864 2707
rect 854 2682 857 2688
rect 814 2672 817 2678
rect 870 2672 873 2738
rect 782 2632 785 2658
rect 790 2622 793 2668
rect 830 2662 833 2668
rect 838 2652 841 2658
rect 802 2648 806 2651
rect 774 2588 785 2591
rect 706 2568 710 2571
rect 766 2542 769 2547
rect 750 2532 753 2538
rect 686 2518 694 2521
rect 686 2482 689 2518
rect 678 2478 686 2481
rect 666 2458 670 2461
rect 630 2452 633 2458
rect 678 2452 681 2478
rect 702 2472 705 2478
rect 742 2472 745 2478
rect 650 2448 662 2451
rect 654 2392 657 2438
rect 702 2422 705 2458
rect 710 2442 713 2468
rect 718 2462 721 2468
rect 726 2462 729 2468
rect 750 2462 753 2468
rect 782 2462 785 2588
rect 798 2562 801 2568
rect 814 2562 817 2568
rect 822 2552 825 2618
rect 830 2582 833 2618
rect 830 2562 833 2568
rect 846 2562 849 2618
rect 830 2542 833 2548
rect 822 2532 825 2538
rect 634 2388 638 2391
rect 670 2362 673 2408
rect 742 2392 745 2458
rect 758 2432 761 2458
rect 774 2432 777 2438
rect 678 2362 681 2368
rect 506 2348 510 2351
rect 530 2348 534 2351
rect 542 2342 545 2348
rect 658 2348 662 2351
rect 574 2342 577 2347
rect 646 2342 649 2348
rect 694 2342 697 2378
rect 718 2352 721 2358
rect 726 2342 729 2378
rect 734 2342 737 2388
rect 758 2362 761 2408
rect 746 2348 750 2351
rect 766 2342 769 2348
rect 522 2338 526 2341
rect 654 2332 657 2338
rect 782 2332 785 2338
rect 554 2288 558 2291
rect 462 2282 465 2288
rect 574 2272 577 2328
rect 450 2258 457 2261
rect 238 2142 241 2158
rect 254 2102 257 2258
rect 262 2091 265 2148
rect 286 2132 289 2138
rect 258 2088 265 2091
rect 286 2082 289 2118
rect 250 2068 254 2071
rect 270 2062 273 2068
rect 222 2052 225 2058
rect 178 2048 182 2051
rect 174 1962 177 1988
rect 190 1952 193 1998
rect 122 1948 126 1951
rect 178 1948 182 1951
rect 190 1931 193 1948
rect 198 1942 201 2038
rect 222 1952 225 2048
rect 230 2022 233 2058
rect 238 2052 241 2058
rect 230 1962 233 1968
rect 250 1958 254 1961
rect 262 1952 265 2018
rect 286 1992 289 2058
rect 294 2052 297 2078
rect 302 1992 305 2258
rect 314 2248 318 2251
rect 382 2232 385 2258
rect 494 2252 497 2259
rect 442 2248 446 2251
rect 328 2203 330 2207
rect 334 2203 337 2207
rect 341 2203 344 2207
rect 358 2192 361 2218
rect 358 2172 361 2178
rect 338 2158 342 2161
rect 314 2118 318 2121
rect 322 2118 329 2121
rect 326 2072 329 2118
rect 310 2052 313 2058
rect 318 2002 321 2068
rect 342 2052 345 2098
rect 350 2092 353 2158
rect 382 2152 385 2228
rect 526 2222 529 2258
rect 574 2222 577 2268
rect 598 2262 601 2268
rect 542 2192 545 2218
rect 614 2192 617 2208
rect 654 2192 657 2328
rect 702 2322 705 2328
rect 678 2262 681 2268
rect 710 2262 713 2288
rect 726 2272 729 2298
rect 758 2272 761 2278
rect 790 2271 793 2508
rect 798 2452 801 2458
rect 806 2342 809 2528
rect 846 2522 849 2548
rect 854 2542 857 2668
rect 878 2572 881 2748
rect 886 2682 889 2828
rect 894 2802 897 2848
rect 926 2842 929 2918
rect 934 2882 937 2898
rect 982 2892 985 2948
rect 1190 2942 1193 2947
rect 1198 2942 1201 3048
rect 1302 3042 1305 3058
rect 1310 3052 1313 3058
rect 1362 3048 1366 3051
rect 1298 3018 1302 3021
rect 1286 2962 1289 2998
rect 1318 2972 1321 3018
rect 1352 3003 1354 3007
rect 1358 3003 1361 3007
rect 1365 3003 1368 3007
rect 1342 2962 1345 2968
rect 1270 2952 1273 2958
rect 1266 2948 1270 2951
rect 1098 2938 1102 2941
rect 1258 2938 1262 2941
rect 1054 2932 1057 2938
rect 1142 2932 1145 2938
rect 1310 2932 1313 2938
rect 1114 2928 1118 2931
rect 1254 2922 1257 2928
rect 1318 2922 1321 2948
rect 1330 2938 1334 2941
rect 1362 2938 1366 2941
rect 1350 2932 1353 2938
rect 1038 2912 1041 2918
rect 942 2882 945 2888
rect 1014 2882 1017 2908
rect 1086 2902 1089 2918
rect 1250 2888 1254 2891
rect 1038 2882 1041 2888
rect 1078 2882 1081 2888
rect 974 2872 977 2878
rect 962 2868 966 2871
rect 998 2862 1001 2878
rect 1014 2862 1017 2878
rect 1042 2868 1046 2871
rect 958 2812 961 2858
rect 966 2832 969 2858
rect 1094 2852 1097 2858
rect 1074 2848 1078 2851
rect 946 2758 950 2761
rect 962 2758 966 2761
rect 902 2752 905 2758
rect 934 2752 937 2758
rect 894 2742 897 2748
rect 902 2692 905 2698
rect 886 2662 889 2678
rect 910 2672 913 2738
rect 918 2732 921 2748
rect 926 2742 929 2748
rect 910 2662 913 2668
rect 918 2662 921 2728
rect 942 2682 945 2718
rect 918 2652 921 2658
rect 934 2652 937 2678
rect 950 2672 953 2748
rect 982 2742 985 2798
rect 1006 2752 1009 2758
rect 1054 2712 1057 2818
rect 1094 2802 1097 2818
rect 1102 2792 1105 2868
rect 1110 2852 1113 2858
rect 1126 2852 1129 2888
rect 1138 2868 1142 2871
rect 1150 2842 1153 2858
rect 1070 2752 1073 2788
rect 1118 2762 1121 2808
rect 1082 2758 1086 2761
rect 1122 2758 1126 2761
rect 1074 2738 1078 2741
rect 990 2663 993 2698
rect 1022 2672 1025 2678
rect 1062 2672 1065 2718
rect 1070 2682 1073 2688
rect 1078 2662 1081 2678
rect 1094 2672 1097 2758
rect 1142 2752 1145 2808
rect 1158 2802 1161 2868
rect 1174 2772 1177 2868
rect 1190 2863 1193 2868
rect 1262 2852 1265 2908
rect 1302 2902 1305 2918
rect 1326 2892 1329 2928
rect 1374 2912 1377 2948
rect 1282 2868 1286 2871
rect 1306 2868 1310 2871
rect 1286 2851 1289 2858
rect 1302 2852 1305 2858
rect 1286 2848 1294 2851
rect 1154 2758 1158 2761
rect 1138 2748 1142 2751
rect 1154 2748 1158 2751
rect 1110 2742 1113 2748
rect 1174 2742 1177 2768
rect 1190 2751 1193 2758
rect 1270 2742 1273 2768
rect 1294 2752 1297 2768
rect 1102 2732 1105 2738
rect 1126 2722 1129 2728
rect 1110 2672 1113 2718
rect 1118 2672 1121 2688
rect 902 2642 905 2648
rect 922 2638 926 2641
rect 854 2532 857 2538
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 861 2503 864 2507
rect 870 2472 873 2558
rect 910 2552 913 2558
rect 818 2468 822 2471
rect 826 2458 830 2461
rect 838 2402 841 2458
rect 846 2382 849 2468
rect 830 2352 833 2368
rect 854 2322 857 2338
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 861 2303 864 2307
rect 790 2268 798 2271
rect 802 2268 806 2271
rect 718 2262 721 2268
rect 782 2262 785 2268
rect 814 2262 817 2268
rect 822 2262 825 2268
rect 666 2258 670 2261
rect 706 2258 710 2261
rect 762 2258 766 2261
rect 686 2252 689 2258
rect 690 2178 694 2181
rect 446 2152 449 2168
rect 666 2158 670 2161
rect 686 2152 689 2158
rect 358 2122 361 2148
rect 422 2142 425 2148
rect 734 2142 737 2258
rect 790 2252 793 2258
rect 750 2222 753 2228
rect 766 2192 769 2198
rect 782 2192 785 2248
rect 790 2222 793 2248
rect 838 2242 841 2278
rect 870 2232 873 2458
rect 878 2452 881 2518
rect 890 2458 894 2461
rect 878 2402 881 2448
rect 894 2442 897 2448
rect 890 2388 894 2391
rect 902 2362 905 2528
rect 914 2468 918 2471
rect 950 2471 953 2618
rect 958 2512 961 2658
rect 970 2568 974 2571
rect 1006 2562 1009 2568
rect 986 2558 990 2561
rect 998 2558 1006 2561
rect 978 2548 982 2551
rect 974 2532 977 2538
rect 998 2482 1001 2558
rect 950 2468 958 2471
rect 986 2468 990 2471
rect 954 2458 958 2461
rect 926 2452 929 2458
rect 934 2452 937 2458
rect 950 2432 953 2438
rect 902 2322 905 2358
rect 926 2352 929 2428
rect 966 2392 969 2468
rect 1014 2462 1017 2568
rect 1022 2522 1025 2658
rect 1046 2592 1049 2648
rect 1078 2572 1081 2658
rect 1086 2652 1089 2668
rect 1086 2632 1089 2638
rect 1086 2592 1089 2628
rect 1062 2552 1065 2558
rect 1062 2542 1065 2548
rect 978 2458 982 2461
rect 1002 2458 1006 2461
rect 1022 2461 1025 2488
rect 1030 2472 1033 2538
rect 1054 2462 1057 2468
rect 1062 2462 1065 2468
rect 1022 2458 1030 2461
rect 1070 2452 1073 2548
rect 1094 2542 1097 2658
rect 1102 2642 1105 2658
rect 1102 2542 1105 2548
rect 1078 2452 1081 2508
rect 1094 2472 1097 2518
rect 990 2442 993 2448
rect 966 2372 969 2388
rect 1022 2382 1025 2448
rect 1070 2442 1073 2448
rect 1042 2438 1046 2441
rect 1058 2438 1062 2441
rect 938 2368 942 2371
rect 938 2348 942 2351
rect 938 2338 942 2341
rect 910 2332 913 2338
rect 982 2332 985 2348
rect 998 2342 1001 2378
rect 1030 2371 1033 2418
rect 1022 2368 1033 2371
rect 1022 2362 1025 2368
rect 982 2322 985 2328
rect 886 2282 889 2318
rect 918 2272 921 2318
rect 990 2302 993 2338
rect 1006 2272 1009 2348
rect 1014 2322 1017 2338
rect 890 2259 894 2262
rect 990 2262 993 2268
rect 998 2262 1001 2268
rect 954 2238 958 2241
rect 746 2188 750 2191
rect 790 2181 793 2218
rect 782 2178 793 2181
rect 966 2182 969 2258
rect 974 2212 977 2248
rect 982 2212 985 2218
rect 1014 2192 1017 2258
rect 1022 2222 1025 2348
rect 1038 2342 1041 2358
rect 1046 2262 1049 2268
rect 1054 2262 1057 2398
rect 1062 2352 1065 2358
rect 1110 2332 1113 2668
rect 1126 2662 1129 2668
rect 1134 2662 1137 2738
rect 1142 2692 1145 2698
rect 1150 2682 1153 2688
rect 1142 2662 1145 2668
rect 1142 2632 1145 2648
rect 1126 2542 1129 2558
rect 1134 2552 1137 2558
rect 1126 2462 1129 2518
rect 1134 2462 1137 2528
rect 1142 2512 1145 2628
rect 1150 2562 1153 2678
rect 1190 2672 1193 2718
rect 1254 2712 1257 2718
rect 1166 2662 1169 2668
rect 1158 2551 1161 2558
rect 1150 2548 1161 2551
rect 1150 2532 1153 2548
rect 1174 2542 1177 2668
rect 1182 2642 1185 2658
rect 1198 2652 1201 2708
rect 1206 2672 1209 2688
rect 1270 2663 1273 2688
rect 1302 2662 1305 2668
rect 1310 2662 1313 2828
rect 1318 2752 1321 2868
rect 1374 2831 1377 2858
rect 1382 2842 1385 3068
rect 1390 3062 1393 3158
rect 1454 3152 1457 3158
rect 1502 3152 1505 3228
rect 1510 3222 1513 3268
rect 1518 3252 1521 3258
rect 1534 3252 1537 3258
rect 1550 3242 1553 3268
rect 1558 3262 1561 3288
rect 1574 3271 1577 3298
rect 1582 3292 1585 3328
rect 1590 3322 1593 3348
rect 1574 3268 1582 3271
rect 1570 3248 1574 3251
rect 1538 3238 1542 3241
rect 1418 3148 1422 3151
rect 1438 3142 1441 3148
rect 1478 3142 1481 3148
rect 1550 3142 1553 3158
rect 1574 3152 1577 3168
rect 1558 3142 1561 3148
rect 1566 3142 1569 3148
rect 1466 3138 1470 3141
rect 1406 3132 1409 3138
rect 1446 3122 1449 3138
rect 1530 3128 1534 3131
rect 1462 3102 1465 3128
rect 1494 3122 1497 3128
rect 1542 3122 1545 3128
rect 1438 3082 1441 3088
rect 1478 3082 1481 3088
rect 1414 3072 1417 3078
rect 1470 3062 1473 3068
rect 1502 3062 1505 3108
rect 1402 3058 1406 3061
rect 1442 3058 1446 3061
rect 1458 3058 1462 3061
rect 1414 3051 1417 3058
rect 1410 3048 1417 3051
rect 1422 3042 1425 3058
rect 1450 3048 1454 3051
rect 1482 3048 1486 3051
rect 1438 3042 1441 3048
rect 1422 3012 1425 3038
rect 1390 2952 1393 2998
rect 1458 2988 1462 2991
rect 1510 2952 1513 3018
rect 1518 2972 1521 3118
rect 1574 3102 1577 3148
rect 1582 3112 1585 3258
rect 1590 3252 1593 3268
rect 1590 3162 1593 3178
rect 1598 3132 1601 3358
rect 1614 3312 1617 3458
rect 1630 3392 1633 3468
rect 1646 3452 1649 3459
rect 1634 3388 1641 3391
rect 1622 3332 1625 3338
rect 1638 3282 1641 3388
rect 1646 3362 1649 3368
rect 1666 3358 1670 3361
rect 1606 3262 1609 3268
rect 1606 3242 1609 3248
rect 1606 3142 1609 3148
rect 1614 3141 1617 3198
rect 1622 3152 1625 3278
rect 1646 3262 1649 3288
rect 1670 3252 1673 3348
rect 1678 3342 1681 3468
rect 1790 3462 1793 3468
rect 1838 3462 1841 3568
rect 1850 3548 1854 3551
rect 1870 3532 1873 3658
rect 1886 3612 1889 3648
rect 1894 3542 1897 3668
rect 1934 3662 1937 3678
rect 1950 3672 1953 3708
rect 1958 3692 1961 3728
rect 1974 3671 1977 3748
rect 1986 3738 1990 3741
rect 1990 3712 1993 3718
rect 2014 3692 2017 3708
rect 1966 3668 1977 3671
rect 1998 3682 2001 3688
rect 1902 3652 1905 3658
rect 1922 3648 1926 3651
rect 1966 3552 1969 3668
rect 1986 3658 1990 3661
rect 1974 3612 1977 3658
rect 1998 3572 2001 3678
rect 2022 3672 2025 3728
rect 2030 3702 2033 3748
rect 2038 3742 2041 3748
rect 2086 3742 2089 3748
rect 2114 3738 2118 3741
rect 2126 3732 2129 3738
rect 2146 3728 2150 3731
rect 2110 3702 2113 3718
rect 2038 3692 2041 3698
rect 2078 3682 2081 3698
rect 2098 3668 2102 3671
rect 2022 3662 2025 3668
rect 2110 3662 2113 3668
rect 2118 3662 2121 3698
rect 2134 3672 2137 3718
rect 2158 3672 2161 3748
rect 2154 3668 2158 3671
rect 2058 3658 2062 3661
rect 2146 3658 2150 3661
rect 2030 3562 2033 3658
rect 1982 3552 1985 3558
rect 2002 3548 2006 3551
rect 2026 3548 2030 3551
rect 1902 3542 1905 3548
rect 1974 3542 1977 3548
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1885 3503 1888 3507
rect 1902 3482 1905 3488
rect 1854 3462 1857 3478
rect 1918 3472 1921 3498
rect 1866 3468 1870 3471
rect 1970 3468 1974 3471
rect 1918 3462 1921 3468
rect 1722 3458 1726 3461
rect 1778 3458 1782 3461
rect 1810 3458 1814 3461
rect 1898 3458 1902 3461
rect 1750 3452 1753 3458
rect 1846 3452 1849 3458
rect 1790 3448 1798 3451
rect 1766 3442 1769 3448
rect 1694 3342 1697 3438
rect 1790 3392 1793 3448
rect 1822 3382 1825 3418
rect 1854 3402 1857 3458
rect 1770 3368 1774 3371
rect 1710 3351 1713 3358
rect 1726 3272 1729 3288
rect 1758 3272 1761 3288
rect 1714 3268 1718 3271
rect 1758 3262 1761 3268
rect 1766 3262 1769 3358
rect 1790 3352 1793 3378
rect 1802 3358 1806 3361
rect 1814 3352 1817 3368
rect 1934 3362 1937 3468
rect 1954 3459 1958 3462
rect 1982 3462 1985 3548
rect 2014 3542 2017 3548
rect 1990 3532 1993 3538
rect 2030 3532 2033 3538
rect 2030 3512 2033 3528
rect 2038 3492 2041 3648
rect 2086 3632 2089 3658
rect 2126 3642 2129 3658
rect 2110 3592 2113 3618
rect 2166 3562 2169 3888
rect 2174 3802 2177 4018
rect 2190 3962 2193 4058
rect 2318 4052 2321 4058
rect 2342 4052 2345 4058
rect 2430 4052 2433 4098
rect 2454 4062 2457 4078
rect 2462 4072 2465 4078
rect 2442 4058 2446 4061
rect 2298 4048 2302 4051
rect 2382 4042 2385 4048
rect 2414 4022 2417 4028
rect 2198 3952 2201 3968
rect 2186 3948 2190 3951
rect 2206 3942 2209 4018
rect 2190 3932 2193 3938
rect 2190 3791 2193 3858
rect 2214 3852 2217 4018
rect 2222 3962 2225 3968
rect 2230 3952 2233 3968
rect 2294 3951 2297 3968
rect 2246 3932 2249 3938
rect 2226 3928 2230 3931
rect 2262 3911 2265 3948
rect 2310 3942 2313 3988
rect 2334 3972 2337 3978
rect 2334 3952 2337 3958
rect 2330 3938 2334 3941
rect 2358 3932 2361 3958
rect 2254 3908 2265 3911
rect 2222 3863 2225 3878
rect 2254 3872 2257 3908
rect 2326 3892 2329 3908
rect 2286 3882 2289 3888
rect 2274 3878 2278 3881
rect 2254 3852 2257 3858
rect 2262 3852 2265 3868
rect 2186 3788 2193 3791
rect 2182 3752 2185 3788
rect 2246 3762 2249 3838
rect 2270 3752 2273 3858
rect 2302 3852 2305 3858
rect 2310 3762 2313 3858
rect 2318 3752 2321 3888
rect 2342 3822 2345 3868
rect 2350 3862 2353 3868
rect 2366 3861 2369 4018
rect 2384 4003 2386 4007
rect 2390 4003 2393 4007
rect 2397 4003 2400 4007
rect 2374 3952 2377 3978
rect 2382 3892 2385 3938
rect 2398 3932 2401 3948
rect 2422 3942 2425 3968
rect 2430 3942 2433 3948
rect 2438 3942 2441 4048
rect 2478 3992 2481 4068
rect 2498 4058 2502 4061
rect 2510 4022 2513 4148
rect 2414 3882 2417 3918
rect 2438 3882 2441 3918
rect 2414 3863 2417 3868
rect 2358 3858 2369 3861
rect 2378 3858 2382 3861
rect 2206 3712 2209 3748
rect 2246 3742 2249 3748
rect 2214 3682 2217 3728
rect 2262 3702 2265 3738
rect 2222 3662 2225 3688
rect 2246 3672 2249 3678
rect 2174 3562 2177 3578
rect 2054 3552 2057 3558
rect 2090 3548 2094 3551
rect 2062 3542 2065 3548
rect 2054 3532 2057 3538
rect 2046 3522 2049 3528
rect 2062 3502 2065 3538
rect 2102 3532 2105 3538
rect 2110 3532 2113 3558
rect 2126 3522 2129 3548
rect 2134 3542 2137 3558
rect 2142 3542 2145 3548
rect 2174 3542 2177 3548
rect 2010 3488 2014 3491
rect 2038 3462 2041 3468
rect 2070 3463 2073 3518
rect 2086 3512 2089 3518
rect 1830 3352 1833 3358
rect 1918 3352 1921 3358
rect 1778 3338 1782 3341
rect 1778 3268 1782 3271
rect 1670 3221 1673 3248
rect 1702 3232 1705 3248
rect 1670 3218 1681 3221
rect 1670 3192 1673 3208
rect 1646 3158 1654 3161
rect 1634 3148 1638 3151
rect 1614 3138 1622 3141
rect 1634 3138 1638 3141
rect 1546 3078 1550 3081
rect 1558 3062 1561 3078
rect 1574 3062 1577 3088
rect 1526 3032 1529 3058
rect 1466 2948 1470 2951
rect 1390 2892 1393 2948
rect 1422 2942 1425 2948
rect 1402 2938 1406 2941
rect 1406 2872 1409 2918
rect 1422 2882 1425 2938
rect 1438 2882 1441 2928
rect 1486 2902 1489 2938
rect 1534 2932 1537 3058
rect 1582 3032 1585 3088
rect 1590 3052 1593 3078
rect 1598 3062 1601 3068
rect 1606 3062 1609 3098
rect 1574 2942 1577 3018
rect 1582 2992 1585 3028
rect 1598 3011 1601 3058
rect 1606 3042 1609 3058
rect 1606 3022 1609 3028
rect 1598 3008 1609 3011
rect 1606 2992 1609 3008
rect 1614 3002 1617 3138
rect 1630 3062 1633 3128
rect 1646 3092 1649 3158
rect 1666 3148 1670 3151
rect 1666 3138 1670 3141
rect 1654 3132 1657 3138
rect 1678 3131 1681 3218
rect 1734 3202 1737 3258
rect 1698 3188 1702 3191
rect 1766 3191 1769 3258
rect 1782 3192 1785 3258
rect 1790 3202 1793 3348
rect 1822 3312 1825 3338
rect 1842 3328 1846 3331
rect 1822 3272 1825 3308
rect 1830 3272 1833 3278
rect 1810 3258 1822 3261
rect 1846 3252 1849 3258
rect 1806 3212 1809 3248
rect 1822 3222 1825 3228
rect 1766 3188 1777 3191
rect 1694 3182 1697 3188
rect 1774 3172 1777 3188
rect 1690 3158 1694 3161
rect 1670 3128 1681 3131
rect 1658 3078 1662 3081
rect 1622 3052 1625 3058
rect 1622 2952 1625 3038
rect 1630 2992 1633 3058
rect 1638 2971 1641 3068
rect 1654 3002 1657 3068
rect 1670 3062 1673 3128
rect 1710 3092 1713 3158
rect 1806 3152 1809 3158
rect 1746 3148 1750 3151
rect 1774 3142 1777 3148
rect 1846 3142 1849 3148
rect 1854 3142 1857 3338
rect 1894 3322 1897 3348
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1885 3303 1888 3307
rect 1894 3272 1897 3288
rect 1910 3272 1913 3278
rect 1870 3242 1873 3268
rect 1870 3222 1873 3238
rect 1862 3212 1865 3218
rect 1902 3162 1905 3258
rect 1918 3252 1921 3288
rect 1934 3272 1937 3358
rect 1950 3342 1953 3368
rect 1982 3362 1985 3458
rect 2038 3442 2041 3448
rect 2086 3392 2089 3508
rect 2110 3501 2113 3518
rect 2142 3501 2145 3538
rect 2150 3532 2153 3538
rect 2110 3498 2121 3501
rect 2102 3422 2105 3458
rect 1958 3352 1961 3358
rect 1966 3342 1969 3348
rect 1974 3322 1977 3328
rect 1958 3252 1961 3258
rect 1934 3182 1937 3188
rect 1982 3161 1985 3358
rect 2014 3352 2017 3368
rect 2030 3362 2033 3368
rect 2062 3358 2070 3361
rect 2054 3352 2057 3358
rect 1994 3348 1998 3351
rect 2042 3338 2046 3341
rect 2006 3332 2009 3338
rect 2030 3282 2033 3288
rect 2010 3218 2014 3221
rect 2014 3182 2017 3188
rect 1974 3158 1985 3161
rect 1974 3152 1977 3158
rect 1990 3152 1993 3158
rect 1942 3142 1945 3148
rect 1982 3142 1985 3148
rect 1998 3142 2001 3178
rect 1806 3132 1809 3138
rect 1794 3128 1798 3131
rect 2014 3122 2017 3128
rect 1798 3112 1801 3118
rect 2022 3111 2025 3218
rect 2030 3192 2033 3258
rect 2038 3252 2041 3268
rect 2046 3262 2049 3278
rect 2046 3232 2049 3238
rect 2062 3192 2065 3358
rect 2078 3342 2081 3348
rect 2102 3342 2105 3348
rect 2102 3272 2105 3308
rect 2094 3242 2097 3268
rect 2110 3262 2113 3378
rect 2118 3372 2121 3498
rect 2134 3498 2145 3501
rect 2134 3492 2137 3498
rect 2146 3488 2150 3491
rect 2142 3432 2145 3448
rect 2158 3402 2161 3468
rect 2170 3458 2174 3461
rect 2142 3362 2145 3368
rect 2126 3342 2129 3348
rect 2134 3322 2137 3358
rect 2166 3352 2169 3408
rect 2162 3338 2166 3341
rect 2070 3222 2073 3238
rect 2110 3232 2113 3238
rect 2042 3178 2049 3181
rect 2046 3152 2049 3178
rect 2038 3148 2046 3151
rect 2014 3108 2025 3111
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1885 3103 1888 3107
rect 1822 3092 1825 3098
rect 1934 3092 1937 3098
rect 1722 3078 1726 3081
rect 1930 3078 1934 3081
rect 1846 3072 1849 3078
rect 1890 3068 1894 3071
rect 1694 3062 1697 3068
rect 1638 2968 1646 2971
rect 1646 2962 1649 2968
rect 1670 2952 1673 3058
rect 1678 3032 1681 3058
rect 1702 3052 1705 3068
rect 1686 3022 1689 3048
rect 1726 3042 1729 3048
rect 1682 2968 1686 2971
rect 1586 2948 1590 2951
rect 1722 2948 1726 2951
rect 1662 2942 1665 2948
rect 1390 2852 1393 2858
rect 1422 2832 1425 2878
rect 1486 2872 1489 2898
rect 1506 2878 1510 2881
rect 1438 2852 1441 2868
rect 1454 2863 1457 2868
rect 1526 2862 1529 2928
rect 1582 2882 1585 2888
rect 1598 2872 1601 2898
rect 1622 2862 1625 2868
rect 1558 2852 1561 2858
rect 1566 2842 1569 2858
rect 1374 2828 1385 2831
rect 1352 2803 1354 2807
rect 1358 2803 1361 2807
rect 1365 2803 1368 2807
rect 1382 2792 1385 2828
rect 1422 2812 1425 2818
rect 1350 2762 1353 2768
rect 1374 2732 1377 2738
rect 1330 2688 1334 2691
rect 1354 2668 1358 2671
rect 1326 2662 1329 2668
rect 1182 2552 1185 2638
rect 1194 2548 1198 2551
rect 1246 2542 1249 2658
rect 1302 2622 1305 2658
rect 1334 2651 1337 2668
rect 1366 2662 1369 2728
rect 1382 2672 1385 2748
rect 1390 2672 1393 2698
rect 1330 2648 1337 2651
rect 1350 2642 1353 2658
rect 1294 2562 1297 2568
rect 1310 2562 1313 2568
rect 1262 2542 1265 2548
rect 1318 2542 1321 2618
rect 1342 2552 1345 2638
rect 1352 2603 1354 2607
rect 1358 2603 1361 2607
rect 1365 2603 1368 2607
rect 1362 2558 1374 2561
rect 1386 2558 1390 2561
rect 1330 2548 1334 2551
rect 1162 2538 1166 2541
rect 1186 2538 1190 2541
rect 1210 2538 1214 2541
rect 1150 2502 1153 2528
rect 1174 2492 1177 2498
rect 1122 2368 1126 2371
rect 1130 2358 1134 2361
rect 1130 2348 1134 2351
rect 1142 2342 1145 2458
rect 1182 2442 1185 2468
rect 1190 2462 1193 2538
rect 1182 2362 1185 2368
rect 1190 2362 1193 2418
rect 1154 2358 1166 2361
rect 1186 2348 1190 2351
rect 1130 2338 1134 2341
rect 1102 2272 1105 2278
rect 1142 2272 1145 2338
rect 1158 2302 1161 2338
rect 1166 2332 1169 2348
rect 1198 2341 1201 2468
rect 1206 2452 1209 2498
rect 1214 2472 1217 2518
rect 1218 2458 1222 2461
rect 1210 2358 1214 2361
rect 1210 2348 1214 2351
rect 1194 2338 1201 2341
rect 1230 2342 1233 2538
rect 1254 2532 1257 2538
rect 1238 2462 1241 2468
rect 1238 2442 1241 2448
rect 1246 2442 1249 2468
rect 1254 2462 1257 2528
rect 1278 2491 1281 2538
rect 1278 2488 1289 2491
rect 1286 2472 1289 2488
rect 1302 2463 1305 2468
rect 1254 2442 1257 2448
rect 1270 2442 1273 2448
rect 1230 2332 1233 2338
rect 1198 2282 1201 2288
rect 1206 2272 1209 2278
rect 1082 2268 1086 2271
rect 1062 2262 1065 2268
rect 1038 2222 1041 2258
rect 774 2162 777 2168
rect 782 2151 785 2178
rect 1046 2172 1049 2258
rect 850 2158 854 2161
rect 774 2148 785 2151
rect 554 2138 558 2141
rect 666 2138 670 2141
rect 354 2038 358 2041
rect 328 2003 330 2007
rect 334 2003 337 2007
rect 341 2003 344 2007
rect 338 1988 342 1991
rect 286 1962 289 1968
rect 254 1942 257 1948
rect 222 1932 225 1938
rect 190 1928 201 1931
rect 102 1882 105 1888
rect 118 1862 121 1908
rect 142 1872 145 1908
rect 182 1882 185 1888
rect 126 1862 129 1868
rect 150 1862 153 1868
rect 190 1862 193 1868
rect 70 1852 73 1859
rect 62 1792 65 1818
rect 142 1742 145 1748
rect 10 1738 14 1741
rect 74 1738 78 1741
rect 62 1672 65 1728
rect 14 1542 17 1668
rect 50 1658 54 1661
rect 38 1542 41 1548
rect 14 1472 17 1538
rect 14 1392 17 1468
rect 50 1458 54 1461
rect 78 1371 81 1738
rect 158 1732 161 1738
rect 94 1692 97 1708
rect 102 1662 105 1668
rect 118 1662 121 1688
rect 106 1648 110 1651
rect 126 1642 129 1668
rect 134 1652 137 1708
rect 158 1672 161 1718
rect 190 1692 193 1748
rect 198 1722 201 1928
rect 206 1802 209 1928
rect 250 1888 254 1891
rect 262 1882 265 1948
rect 270 1892 273 1958
rect 278 1952 281 1958
rect 322 1948 326 1951
rect 302 1931 305 1948
rect 366 1942 369 2138
rect 462 2082 465 2098
rect 386 2078 390 2081
rect 314 1938 321 1941
rect 338 1938 342 1941
rect 302 1928 313 1931
rect 282 1918 286 1921
rect 310 1892 313 1928
rect 318 1922 321 1938
rect 318 1882 321 1888
rect 282 1878 286 1881
rect 374 1872 377 1948
rect 382 1912 385 2068
rect 398 2062 401 2068
rect 470 2062 473 2138
rect 486 1992 489 2138
rect 638 2112 641 2118
rect 530 2088 534 2091
rect 542 2082 545 2098
rect 550 2082 553 2088
rect 558 2082 561 2088
rect 566 2082 569 2098
rect 574 2092 577 2098
rect 526 2062 529 2078
rect 582 2062 585 2078
rect 606 2072 609 2078
rect 606 2062 609 2068
rect 494 2052 497 2059
rect 614 2052 617 2058
rect 634 2048 638 2051
rect 662 2032 665 2068
rect 710 2042 713 2128
rect 726 2062 729 2088
rect 674 2038 678 2041
rect 434 1968 438 1971
rect 422 1962 425 1968
rect 470 1952 473 1978
rect 734 1972 737 2068
rect 750 2032 753 2138
rect 758 2102 761 2138
rect 766 2042 769 2048
rect 754 1988 758 1991
rect 626 1968 630 1971
rect 758 1962 761 1968
rect 654 1952 657 1958
rect 774 1952 777 2148
rect 790 2132 793 2138
rect 798 2112 801 2138
rect 790 2072 793 2078
rect 806 2062 809 2148
rect 822 2142 825 2158
rect 846 2122 849 2148
rect 854 2142 857 2148
rect 862 2142 865 2168
rect 934 2152 937 2158
rect 1018 2148 1022 2151
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 861 2103 864 2107
rect 834 2088 838 2091
rect 822 2072 825 2078
rect 794 2058 798 2061
rect 818 2058 822 2061
rect 826 2048 830 2051
rect 798 2042 801 2048
rect 814 2042 817 2048
rect 782 1972 785 2018
rect 394 1948 398 1951
rect 398 1932 401 1938
rect 422 1912 425 1928
rect 382 1891 385 1908
rect 398 1892 401 1908
rect 382 1888 393 1891
rect 254 1852 257 1858
rect 238 1792 241 1798
rect 262 1792 265 1868
rect 286 1812 289 1868
rect 334 1862 337 1868
rect 382 1862 385 1878
rect 390 1862 393 1888
rect 430 1862 433 1918
rect 454 1912 457 1928
rect 470 1901 473 1948
rect 762 1948 766 1951
rect 502 1922 505 1947
rect 574 1942 577 1948
rect 646 1942 649 1948
rect 590 1932 593 1938
rect 670 1932 673 1938
rect 694 1932 697 1948
rect 622 1928 630 1931
rect 642 1928 646 1931
rect 462 1898 473 1901
rect 462 1882 465 1898
rect 622 1892 625 1928
rect 602 1888 606 1891
rect 634 1878 638 1881
rect 746 1878 750 1881
rect 510 1872 513 1878
rect 614 1872 617 1878
rect 702 1872 705 1878
rect 766 1872 769 1918
rect 690 1868 694 1871
rect 462 1863 465 1868
rect 346 1858 350 1861
rect 378 1858 382 1861
rect 542 1862 545 1868
rect 718 1862 721 1868
rect 506 1858 510 1861
rect 610 1858 614 1861
rect 682 1858 686 1861
rect 698 1858 702 1861
rect 282 1748 286 1751
rect 254 1742 257 1748
rect 166 1672 169 1678
rect 154 1658 158 1661
rect 142 1652 145 1658
rect 174 1642 177 1658
rect 190 1622 193 1658
rect 206 1651 209 1728
rect 238 1672 241 1728
rect 254 1702 257 1738
rect 294 1712 297 1858
rect 358 1841 361 1858
rect 494 1842 497 1858
rect 358 1838 369 1841
rect 328 1803 330 1807
rect 334 1803 337 1807
rect 341 1803 344 1807
rect 334 1712 337 1718
rect 342 1701 345 1728
rect 334 1698 345 1701
rect 254 1681 257 1698
rect 334 1692 337 1698
rect 358 1692 361 1748
rect 254 1678 265 1681
rect 218 1668 222 1671
rect 202 1648 209 1651
rect 214 1652 217 1658
rect 190 1592 193 1618
rect 98 1568 102 1571
rect 134 1562 137 1568
rect 138 1558 142 1561
rect 102 1552 105 1558
rect 130 1548 134 1551
rect 118 1542 121 1548
rect 106 1538 110 1541
rect 94 1482 97 1488
rect 102 1452 105 1468
rect 118 1462 121 1508
rect 126 1502 129 1538
rect 126 1472 129 1498
rect 110 1452 113 1458
rect 70 1368 81 1371
rect 70 1342 73 1368
rect 110 1352 113 1358
rect 70 1332 73 1338
rect 86 1322 89 1338
rect 14 1272 17 1318
rect 106 1268 110 1271
rect 14 1142 17 1268
rect 38 1262 41 1268
rect 118 1262 121 1458
rect 126 1342 129 1468
rect 134 1452 137 1478
rect 142 1462 145 1468
rect 150 1462 153 1548
rect 158 1472 161 1538
rect 166 1532 169 1558
rect 206 1552 209 1638
rect 222 1592 225 1658
rect 254 1652 257 1659
rect 254 1562 257 1568
rect 242 1558 246 1561
rect 218 1548 222 1551
rect 250 1548 254 1551
rect 174 1522 177 1528
rect 206 1521 209 1548
rect 214 1531 217 1538
rect 214 1528 222 1531
rect 206 1518 217 1521
rect 190 1481 193 1518
rect 190 1478 198 1481
rect 166 1472 169 1478
rect 158 1462 161 1468
rect 198 1462 201 1468
rect 186 1458 190 1461
rect 150 1292 153 1458
rect 170 1448 174 1451
rect 170 1368 174 1371
rect 206 1362 209 1368
rect 194 1348 198 1351
rect 170 1338 174 1341
rect 182 1302 185 1348
rect 214 1322 217 1518
rect 238 1462 241 1498
rect 246 1462 249 1538
rect 262 1462 265 1678
rect 334 1652 337 1668
rect 346 1658 350 1661
rect 270 1572 273 1578
rect 310 1552 313 1588
rect 318 1582 321 1618
rect 328 1603 330 1607
rect 334 1603 337 1607
rect 341 1603 344 1607
rect 330 1548 334 1551
rect 278 1542 281 1548
rect 222 1352 225 1358
rect 182 1282 185 1288
rect 222 1282 225 1348
rect 230 1342 233 1458
rect 246 1392 249 1438
rect 278 1362 281 1538
rect 310 1492 313 1528
rect 326 1502 329 1538
rect 342 1532 345 1548
rect 366 1532 369 1838
rect 430 1782 433 1788
rect 378 1758 382 1761
rect 374 1742 377 1748
rect 398 1742 401 1768
rect 418 1758 422 1761
rect 434 1748 438 1751
rect 418 1738 422 1741
rect 382 1692 385 1718
rect 374 1652 377 1658
rect 382 1612 385 1688
rect 390 1682 393 1708
rect 398 1692 401 1718
rect 398 1672 401 1688
rect 406 1682 409 1718
rect 438 1702 441 1738
rect 398 1622 401 1658
rect 422 1652 425 1678
rect 438 1672 441 1698
rect 406 1582 409 1618
rect 374 1552 377 1558
rect 382 1552 385 1558
rect 398 1552 401 1568
rect 422 1562 425 1578
rect 414 1552 417 1558
rect 430 1551 433 1608
rect 438 1592 441 1648
rect 454 1642 457 1758
rect 518 1752 521 1828
rect 526 1802 529 1858
rect 550 1832 553 1858
rect 570 1848 574 1851
rect 582 1782 585 1858
rect 598 1842 601 1848
rect 510 1742 513 1748
rect 478 1702 481 1718
rect 462 1652 465 1658
rect 478 1552 481 1648
rect 430 1548 438 1551
rect 342 1512 345 1528
rect 390 1522 393 1538
rect 350 1492 353 1498
rect 298 1488 302 1491
rect 302 1472 305 1478
rect 310 1392 313 1458
rect 278 1352 281 1358
rect 310 1352 313 1358
rect 266 1348 270 1351
rect 318 1342 321 1488
rect 374 1472 377 1478
rect 382 1472 385 1488
rect 414 1482 417 1518
rect 390 1462 393 1468
rect 430 1462 433 1548
rect 510 1542 513 1738
rect 526 1692 529 1778
rect 586 1758 590 1761
rect 542 1751 545 1758
rect 586 1748 590 1751
rect 578 1738 582 1741
rect 558 1732 561 1738
rect 518 1682 521 1688
rect 542 1670 545 1678
rect 558 1672 561 1688
rect 562 1668 566 1671
rect 550 1642 553 1668
rect 582 1652 585 1658
rect 590 1652 593 1698
rect 598 1672 601 1758
rect 614 1732 617 1738
rect 646 1682 649 1858
rect 654 1752 657 1818
rect 670 1812 673 1858
rect 710 1852 713 1858
rect 710 1792 713 1808
rect 718 1751 721 1858
rect 726 1812 729 1868
rect 742 1762 745 1818
rect 750 1812 753 1868
rect 762 1858 766 1861
rect 766 1792 769 1838
rect 774 1812 777 1948
rect 790 1942 793 1968
rect 814 1962 817 1998
rect 802 1948 806 1951
rect 782 1852 785 1908
rect 798 1772 801 1948
rect 806 1932 809 1938
rect 830 1892 833 1978
rect 862 1972 865 2068
rect 870 2062 873 2138
rect 934 2092 937 2138
rect 1006 2132 1009 2138
rect 878 2082 881 2088
rect 938 2078 942 2081
rect 878 2072 881 2078
rect 926 2072 929 2078
rect 1006 2072 1009 2128
rect 910 2062 913 2068
rect 954 2058 958 2061
rect 870 1942 873 1948
rect 862 1932 865 1938
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 861 1903 864 1907
rect 838 1882 841 1898
rect 878 1872 881 2058
rect 926 2052 929 2058
rect 886 2002 889 2018
rect 902 2012 905 2038
rect 902 1992 905 2008
rect 938 1958 942 1961
rect 934 1882 937 1928
rect 810 1868 814 1871
rect 878 1862 881 1868
rect 942 1862 945 1868
rect 810 1858 814 1861
rect 822 1842 825 1858
rect 846 1852 849 1858
rect 854 1832 857 1858
rect 710 1748 721 1751
rect 730 1748 734 1751
rect 662 1672 665 1738
rect 610 1668 614 1671
rect 642 1668 646 1671
rect 610 1658 614 1661
rect 614 1648 622 1651
rect 574 1592 577 1628
rect 518 1552 521 1578
rect 590 1552 593 1638
rect 614 1632 617 1648
rect 622 1592 625 1598
rect 638 1582 641 1618
rect 646 1612 649 1658
rect 686 1632 689 1658
rect 598 1552 601 1578
rect 606 1562 609 1578
rect 626 1548 630 1551
rect 450 1538 454 1541
rect 438 1472 441 1528
rect 462 1492 465 1518
rect 478 1492 481 1528
rect 446 1472 449 1478
rect 346 1458 350 1461
rect 362 1458 366 1461
rect 430 1452 433 1458
rect 438 1452 441 1468
rect 502 1462 505 1468
rect 450 1458 454 1461
rect 350 1442 353 1448
rect 328 1403 330 1407
rect 334 1403 337 1407
rect 341 1403 344 1407
rect 234 1338 238 1341
rect 274 1338 278 1341
rect 130 1268 134 1271
rect 158 1262 161 1268
rect 130 1258 134 1261
rect 102 1252 105 1258
rect 138 1248 142 1251
rect 94 1242 97 1248
rect 150 1221 153 1258
rect 158 1232 161 1258
rect 190 1252 193 1278
rect 206 1262 209 1268
rect 238 1262 241 1318
rect 246 1262 249 1298
rect 170 1238 174 1241
rect 150 1218 161 1221
rect 158 1182 161 1218
rect 150 1172 153 1178
rect 94 1162 97 1168
rect 102 1162 105 1168
rect 130 1158 134 1161
rect 158 1152 161 1178
rect 50 1148 54 1151
rect 98 1148 102 1151
rect 122 1148 126 1151
rect 166 1142 169 1158
rect 130 1138 134 1141
rect 14 1072 17 1138
rect 158 1132 161 1138
rect 38 1062 41 1078
rect 62 1072 65 1078
rect 38 952 41 958
rect 30 882 33 928
rect 42 858 46 861
rect 62 752 65 858
rect 78 832 81 1118
rect 118 1072 121 1078
rect 126 1062 129 1078
rect 150 1062 153 1088
rect 174 1082 177 1238
rect 214 1182 217 1218
rect 182 1162 185 1168
rect 190 1162 193 1168
rect 214 1152 217 1178
rect 230 1172 233 1178
rect 202 1148 206 1151
rect 238 1151 241 1258
rect 254 1252 257 1258
rect 250 1158 257 1161
rect 238 1148 246 1151
rect 226 1138 230 1141
rect 214 1122 217 1138
rect 182 1112 185 1118
rect 158 1062 161 1078
rect 174 1062 177 1068
rect 190 1063 193 1118
rect 254 1092 257 1158
rect 262 1142 265 1338
rect 270 1262 273 1268
rect 290 1258 294 1261
rect 278 1242 281 1258
rect 328 1203 330 1207
rect 334 1203 337 1207
rect 341 1203 344 1207
rect 262 1122 265 1138
rect 262 1072 265 1118
rect 270 1102 273 1118
rect 114 1058 118 1061
rect 146 1058 150 1061
rect 190 1058 193 1059
rect 266 1058 270 1061
rect 98 968 102 971
rect 134 962 137 968
rect 114 958 118 961
rect 114 948 121 951
rect 106 938 110 941
rect 118 912 121 948
rect 158 951 161 998
rect 198 972 201 978
rect 182 962 185 968
rect 154 948 161 951
rect 150 922 153 948
rect 158 902 161 938
rect 166 932 169 958
rect 206 951 209 1018
rect 222 992 225 1028
rect 254 972 257 1018
rect 202 948 209 951
rect 226 948 230 951
rect 98 888 102 891
rect 150 882 153 888
rect 158 872 161 898
rect 102 852 105 858
rect 110 842 113 868
rect 166 862 169 918
rect 174 882 177 918
rect 186 868 190 871
rect 198 862 201 948
rect 238 942 241 958
rect 262 952 265 958
rect 250 948 254 951
rect 270 942 273 958
rect 278 952 281 1148
rect 286 1052 289 1118
rect 302 1102 305 1138
rect 294 1072 297 1078
rect 302 1062 305 1098
rect 326 1072 329 1178
rect 342 1092 345 1148
rect 350 1142 353 1258
rect 366 1092 369 1438
rect 406 1402 409 1448
rect 430 1422 433 1428
rect 378 1347 382 1350
rect 398 1342 401 1348
rect 414 1342 417 1348
rect 398 1272 401 1338
rect 430 1292 433 1408
rect 454 1382 457 1418
rect 470 1392 473 1448
rect 478 1412 481 1448
rect 494 1392 497 1458
rect 478 1332 481 1338
rect 486 1332 489 1388
rect 502 1362 505 1378
rect 486 1292 489 1328
rect 450 1288 454 1291
rect 438 1272 441 1278
rect 494 1272 497 1348
rect 510 1332 513 1468
rect 558 1362 561 1548
rect 586 1538 590 1541
rect 606 1538 614 1541
rect 578 1518 582 1521
rect 566 1482 569 1488
rect 582 1472 585 1508
rect 590 1462 593 1518
rect 606 1492 609 1538
rect 638 1492 641 1558
rect 654 1552 657 1618
rect 686 1592 689 1608
rect 670 1552 673 1558
rect 702 1552 705 1588
rect 710 1572 713 1748
rect 750 1742 753 1748
rect 718 1712 721 1738
rect 758 1731 761 1758
rect 798 1752 801 1768
rect 786 1748 790 1751
rect 830 1742 833 1818
rect 902 1812 905 1858
rect 950 1762 953 2038
rect 966 1951 969 2018
rect 962 1948 969 1951
rect 982 1952 985 1958
rect 990 1952 993 1998
rect 958 1922 961 1948
rect 998 1942 1001 1948
rect 966 1932 969 1938
rect 1006 1932 1009 2068
rect 1018 2058 1022 2061
rect 1054 1952 1057 2258
rect 1086 2182 1089 2258
rect 1118 2252 1121 2268
rect 1138 2259 1142 2262
rect 1214 2262 1217 2268
rect 1230 2262 1233 2328
rect 1246 2302 1249 2438
rect 1254 2352 1257 2358
rect 1262 2272 1265 2278
rect 1270 2262 1273 2408
rect 1318 2391 1321 2498
rect 1326 2462 1329 2548
rect 1398 2542 1401 2788
rect 1406 2782 1409 2808
rect 1406 2772 1409 2778
rect 1438 2752 1441 2838
rect 1518 2812 1521 2818
rect 1534 2792 1537 2828
rect 1550 2791 1553 2818
rect 1574 2792 1577 2818
rect 1550 2788 1561 2791
rect 1450 2768 1454 2771
rect 1474 2758 1478 2761
rect 1414 2748 1422 2751
rect 1478 2748 1486 2751
rect 1406 2682 1409 2718
rect 1414 2672 1417 2748
rect 1430 2712 1433 2738
rect 1438 2732 1441 2738
rect 1406 2662 1409 2668
rect 1338 2538 1342 2541
rect 1366 2532 1369 2538
rect 1406 2492 1409 2648
rect 1414 2632 1417 2668
rect 1462 2662 1465 2748
rect 1478 2692 1481 2748
rect 1490 2738 1494 2741
rect 1502 2732 1505 2758
rect 1542 2752 1545 2758
rect 1506 2718 1510 2721
rect 1518 2682 1521 2748
rect 1550 2742 1553 2778
rect 1558 2762 1561 2788
rect 1638 2772 1641 2858
rect 1670 2812 1673 2948
rect 1766 2942 1769 3058
rect 1782 3032 1785 3058
rect 1822 3032 1825 3048
rect 1798 2982 1801 2988
rect 1826 2948 1830 2951
rect 1782 2942 1785 2948
rect 1678 2832 1681 2938
rect 1702 2862 1705 2868
rect 1710 2862 1713 2898
rect 1742 2862 1745 2928
rect 1766 2892 1769 2938
rect 1814 2932 1817 2938
rect 1750 2862 1753 2868
rect 1734 2852 1737 2858
rect 1690 2848 1694 2851
rect 1574 2762 1577 2768
rect 1638 2752 1641 2768
rect 1562 2748 1566 2751
rect 1574 2742 1577 2748
rect 1542 2732 1545 2738
rect 1526 2692 1529 2728
rect 1582 2692 1585 2718
rect 1450 2658 1454 2661
rect 1422 2642 1425 2658
rect 1442 2648 1446 2651
rect 1422 2612 1425 2638
rect 1470 2622 1473 2668
rect 1506 2659 1510 2662
rect 1430 2552 1433 2558
rect 1418 2548 1422 2551
rect 1366 2482 1369 2488
rect 1414 2472 1417 2478
rect 1394 2468 1398 2471
rect 1406 2452 1409 2458
rect 1354 2448 1358 2451
rect 1352 2403 1354 2407
rect 1358 2403 1361 2407
rect 1365 2403 1368 2407
rect 1382 2398 1390 2401
rect 1382 2392 1385 2398
rect 1314 2388 1321 2391
rect 1318 2352 1321 2378
rect 1326 2342 1329 2388
rect 1378 2348 1382 2351
rect 1390 2342 1393 2378
rect 1342 2332 1345 2338
rect 1382 2292 1385 2328
rect 1398 2321 1401 2408
rect 1422 2352 1425 2548
rect 1446 2532 1449 2538
rect 1438 2462 1441 2518
rect 1430 2412 1433 2458
rect 1438 2352 1441 2428
rect 1446 2352 1449 2468
rect 1454 2442 1457 2548
rect 1478 2542 1481 2628
rect 1510 2552 1513 2638
rect 1518 2572 1521 2668
rect 1526 2632 1529 2688
rect 1574 2682 1577 2688
rect 1590 2662 1593 2708
rect 1606 2672 1609 2728
rect 1614 2692 1617 2748
rect 1646 2682 1649 2688
rect 1622 2672 1625 2678
rect 1654 2672 1657 2708
rect 1598 2662 1601 2668
rect 1606 2662 1609 2668
rect 1566 2642 1569 2648
rect 1542 2592 1545 2618
rect 1526 2568 1534 2571
rect 1526 2562 1529 2568
rect 1554 2558 1558 2561
rect 1566 2552 1569 2608
rect 1582 2572 1585 2628
rect 1590 2612 1593 2658
rect 1598 2552 1601 2658
rect 1630 2652 1633 2658
rect 1662 2631 1665 2688
rect 1654 2628 1665 2631
rect 1678 2652 1681 2738
rect 1686 2682 1689 2748
rect 1702 2732 1705 2738
rect 1710 2682 1713 2738
rect 1686 2662 1689 2668
rect 1702 2662 1705 2668
rect 1710 2662 1713 2668
rect 1698 2658 1702 2661
rect 1614 2552 1617 2558
rect 1622 2552 1625 2558
rect 1654 2552 1657 2628
rect 1666 2618 1670 2621
rect 1530 2548 1534 2551
rect 1586 2548 1590 2551
rect 1482 2538 1486 2541
rect 1562 2538 1566 2541
rect 1462 2452 1465 2508
rect 1486 2502 1489 2528
rect 1470 2462 1473 2468
rect 1474 2438 1478 2441
rect 1454 2392 1457 2428
rect 1486 2392 1489 2398
rect 1390 2318 1401 2321
rect 1294 2282 1297 2288
rect 1390 2282 1393 2318
rect 1282 2278 1286 2281
rect 1338 2278 1342 2281
rect 1278 2262 1281 2278
rect 1258 2258 1262 2261
rect 1206 2182 1209 2188
rect 1090 2148 1094 2151
rect 1102 2148 1110 2151
rect 1070 2142 1073 2148
rect 1074 2138 1081 2141
rect 1062 2102 1065 2118
rect 1066 2088 1070 2091
rect 1078 2072 1081 2138
rect 1086 2102 1089 2128
rect 1086 2070 1089 2098
rect 1102 2092 1105 2148
rect 1110 2142 1113 2148
rect 1110 2062 1113 2078
rect 1126 2072 1129 2178
rect 1214 2152 1217 2218
rect 1238 2192 1241 2248
rect 1162 2148 1166 2151
rect 1230 2142 1233 2148
rect 1246 2142 1249 2258
rect 1286 2242 1289 2258
rect 1278 2162 1281 2218
rect 1142 2122 1145 2128
rect 1158 2082 1161 2088
rect 1222 2072 1225 2118
rect 1122 2068 1126 2071
rect 1194 2068 1198 2071
rect 1210 2068 1214 2071
rect 1142 2062 1145 2068
rect 1130 2058 1134 2061
rect 1122 1988 1126 1991
rect 1118 1978 1134 1981
rect 1118 1952 1121 1978
rect 1126 1952 1129 1968
rect 1066 1948 1070 1951
rect 958 1802 961 1918
rect 1022 1902 1025 1948
rect 1018 1888 1022 1891
rect 1026 1868 1030 1871
rect 1038 1822 1041 1938
rect 1070 1872 1073 1888
rect 1062 1862 1065 1868
rect 1078 1862 1081 1898
rect 1050 1858 1054 1861
rect 914 1758 918 1761
rect 1038 1752 1041 1818
rect 850 1747 854 1750
rect 970 1748 974 1751
rect 1018 1748 1022 1751
rect 938 1738 942 1741
rect 754 1728 761 1731
rect 766 1722 769 1728
rect 746 1688 750 1691
rect 750 1672 753 1678
rect 750 1662 753 1668
rect 758 1642 761 1658
rect 782 1652 785 1688
rect 726 1591 729 1638
rect 762 1628 766 1631
rect 718 1588 729 1591
rect 798 1612 801 1658
rect 646 1542 649 1548
rect 654 1542 657 1548
rect 662 1542 665 1548
rect 718 1542 721 1588
rect 654 1492 657 1528
rect 614 1472 617 1478
rect 654 1472 657 1488
rect 678 1462 681 1488
rect 618 1458 622 1461
rect 530 1358 534 1361
rect 558 1352 561 1358
rect 522 1348 526 1351
rect 590 1351 593 1418
rect 534 1342 537 1348
rect 622 1342 625 1348
rect 418 1268 422 1271
rect 502 1262 505 1318
rect 526 1312 529 1338
rect 558 1332 561 1338
rect 598 1272 601 1278
rect 418 1258 422 1261
rect 374 1252 377 1258
rect 438 1162 441 1168
rect 454 1162 457 1168
rect 426 1158 430 1161
rect 406 1152 409 1158
rect 374 1092 377 1098
rect 294 1052 297 1058
rect 286 962 289 1048
rect 318 1042 321 1048
rect 326 1022 329 1068
rect 334 1062 337 1088
rect 390 1062 393 1148
rect 422 1142 425 1148
rect 486 1142 489 1258
rect 494 1142 497 1158
rect 398 1132 401 1138
rect 414 1072 417 1138
rect 430 1122 433 1138
rect 434 1078 438 1081
rect 374 1052 377 1058
rect 302 962 305 1018
rect 328 1003 330 1007
rect 334 1003 337 1007
rect 341 1003 344 1007
rect 322 968 326 971
rect 310 942 313 968
rect 282 938 286 941
rect 206 922 209 938
rect 214 892 217 938
rect 222 892 225 938
rect 238 862 241 888
rect 246 872 249 878
rect 122 858 126 861
rect 134 842 137 858
rect 214 852 217 858
rect 34 748 38 751
rect 10 738 14 741
rect 34 738 38 741
rect 62 672 65 678
rect 38 662 41 668
rect 70 662 73 668
rect 78 662 81 828
rect 118 752 121 768
rect 166 762 169 818
rect 154 748 158 751
rect 102 742 105 748
rect 118 742 121 748
rect 182 722 185 848
rect 222 841 225 848
rect 214 838 225 841
rect 202 758 206 761
rect 206 742 209 748
rect 194 718 198 721
rect 174 692 177 708
rect 182 682 185 718
rect 214 692 217 838
rect 226 748 230 751
rect 230 732 233 738
rect 230 702 233 728
rect 222 682 225 688
rect 126 672 129 678
rect 134 672 137 678
rect 230 672 233 698
rect 58 658 62 661
rect 14 462 17 658
rect 46 652 49 658
rect 78 642 81 658
rect 30 551 33 618
rect 30 482 33 528
rect 46 462 49 488
rect 6 342 9 348
rect 6 262 9 308
rect 38 292 41 318
rect 22 282 25 288
rect 54 262 57 638
rect 78 552 81 618
rect 94 592 97 668
rect 102 652 105 668
rect 122 658 126 661
rect 134 592 137 668
rect 158 662 161 668
rect 174 642 177 648
rect 190 602 193 618
rect 198 612 201 658
rect 186 588 190 591
rect 206 562 209 668
rect 246 661 249 788
rect 262 772 265 868
rect 262 742 265 768
rect 278 752 281 938
rect 270 722 273 748
rect 262 672 265 678
rect 294 672 297 898
rect 302 862 305 918
rect 334 892 337 958
rect 350 952 353 958
rect 366 952 369 1048
rect 346 948 350 951
rect 326 842 329 858
rect 350 812 353 818
rect 328 803 330 807
rect 334 803 337 807
rect 341 803 344 807
rect 266 668 270 671
rect 302 662 305 668
rect 242 658 249 661
rect 274 658 278 661
rect 238 572 241 618
rect 126 551 129 558
rect 230 542 233 548
rect 62 532 65 538
rect 110 532 113 538
rect 206 532 209 538
rect 118 462 121 468
rect 126 462 129 508
rect 186 488 190 491
rect 238 482 241 538
rect 246 512 249 658
rect 254 642 257 648
rect 270 632 273 638
rect 286 592 289 638
rect 318 552 321 778
rect 358 762 361 938
rect 374 932 377 1008
rect 398 991 401 1068
rect 430 1063 433 1068
rect 430 1058 433 1059
rect 454 992 457 1118
rect 486 1082 489 1138
rect 494 1092 497 1138
rect 510 1132 513 1148
rect 526 1082 529 1088
rect 538 1058 542 1061
rect 398 988 409 991
rect 398 962 401 968
rect 394 948 398 951
rect 382 882 385 928
rect 398 922 401 928
rect 406 912 409 988
rect 414 952 417 958
rect 438 952 441 978
rect 470 952 473 958
rect 550 952 553 1238
rect 574 1232 577 1258
rect 562 1158 566 1161
rect 606 1152 609 1158
rect 614 1152 617 1278
rect 638 1252 641 1448
rect 654 1392 657 1398
rect 718 1352 721 1538
rect 734 1472 737 1488
rect 750 1462 753 1498
rect 758 1492 761 1548
rect 774 1462 777 1478
rect 790 1472 793 1478
rect 786 1458 790 1461
rect 754 1378 758 1381
rect 758 1368 766 1371
rect 758 1352 761 1368
rect 766 1352 769 1358
rect 698 1348 702 1351
rect 670 1342 673 1348
rect 718 1342 721 1348
rect 750 1338 758 1341
rect 750 1302 753 1338
rect 774 1322 777 1458
rect 782 1352 785 1418
rect 790 1372 793 1378
rect 738 1288 742 1291
rect 662 1262 665 1268
rect 702 1262 705 1278
rect 750 1272 753 1298
rect 770 1278 774 1281
rect 750 1262 753 1268
rect 758 1262 761 1268
rect 782 1262 785 1348
rect 790 1282 793 1368
rect 798 1351 801 1608
rect 806 1422 809 1738
rect 830 1732 833 1738
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 861 1703 864 1707
rect 902 1692 905 1738
rect 926 1722 929 1738
rect 914 1718 918 1721
rect 894 1682 897 1688
rect 870 1672 873 1678
rect 814 1632 817 1668
rect 842 1648 846 1651
rect 878 1642 881 1658
rect 838 1592 841 1628
rect 818 1548 822 1551
rect 878 1532 881 1538
rect 814 1502 817 1518
rect 814 1362 817 1498
rect 826 1488 830 1491
rect 838 1471 841 1518
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 861 1503 864 1507
rect 830 1468 841 1471
rect 798 1348 806 1351
rect 830 1342 833 1468
rect 846 1462 849 1488
rect 894 1482 897 1668
rect 910 1662 913 1668
rect 906 1548 910 1551
rect 918 1492 921 1528
rect 926 1482 929 1668
rect 942 1572 945 1668
rect 950 1662 953 1678
rect 958 1592 961 1608
rect 914 1468 918 1471
rect 870 1462 873 1468
rect 838 1442 841 1458
rect 902 1451 905 1458
rect 902 1448 913 1451
rect 838 1422 841 1438
rect 886 1432 889 1438
rect 910 1362 913 1448
rect 870 1342 873 1348
rect 798 1282 801 1288
rect 806 1282 809 1288
rect 830 1282 833 1338
rect 846 1332 849 1338
rect 926 1331 929 1478
rect 942 1472 945 1568
rect 966 1382 969 1748
rect 1054 1742 1057 1858
rect 1074 1768 1078 1771
rect 1086 1762 1089 1928
rect 1094 1862 1097 1868
rect 1102 1862 1105 1878
rect 1110 1872 1113 1898
rect 1118 1862 1121 1938
rect 1126 1922 1129 1938
rect 1134 1932 1137 1948
rect 1134 1892 1137 1908
rect 1142 1882 1145 2058
rect 1166 2012 1169 2068
rect 1178 2058 1182 2061
rect 1218 2058 1222 2061
rect 1190 2042 1193 2048
rect 1178 2028 1182 2031
rect 1230 2022 1233 2138
rect 1270 2132 1273 2148
rect 1270 2092 1273 2118
rect 1242 2078 1246 2081
rect 1238 2052 1241 2068
rect 1246 2062 1249 2068
rect 1254 2062 1257 2078
rect 1294 2072 1297 2258
rect 1310 2112 1313 2258
rect 1318 2252 1321 2258
rect 1342 2242 1345 2278
rect 1350 2231 1353 2268
rect 1366 2262 1369 2278
rect 1398 2272 1401 2308
rect 1406 2302 1409 2318
rect 1406 2262 1409 2278
rect 1342 2228 1353 2231
rect 1310 2062 1313 2068
rect 1318 2062 1321 2178
rect 1342 2122 1345 2228
rect 1352 2203 1354 2207
rect 1358 2203 1361 2207
rect 1365 2203 1368 2207
rect 1374 2152 1377 2208
rect 1422 2202 1425 2348
rect 1430 2342 1433 2348
rect 1446 2272 1449 2338
rect 1462 2332 1465 2348
rect 1478 2342 1481 2348
rect 1494 2342 1497 2498
rect 1526 2492 1529 2498
rect 1506 2468 1510 2471
rect 1518 2461 1521 2488
rect 1514 2458 1521 2461
rect 1534 2472 1537 2538
rect 1550 2532 1553 2538
rect 1590 2532 1593 2538
rect 1558 2492 1561 2508
rect 1502 2362 1505 2408
rect 1510 2392 1513 2448
rect 1502 2352 1505 2358
rect 1518 2342 1521 2398
rect 1526 2362 1529 2418
rect 1534 2402 1537 2468
rect 1546 2458 1550 2461
rect 1578 2458 1582 2461
rect 1550 2352 1553 2458
rect 1558 2352 1561 2368
rect 1590 2352 1593 2518
rect 1598 2502 1601 2548
rect 1630 2542 1633 2548
rect 1662 2542 1665 2548
rect 1618 2468 1622 2471
rect 1606 2462 1609 2468
rect 1630 2462 1633 2518
rect 1638 2462 1641 2518
rect 1678 2512 1681 2648
rect 1694 2551 1697 2558
rect 1646 2482 1649 2488
rect 1598 2362 1601 2418
rect 1614 2372 1617 2458
rect 1630 2392 1633 2458
rect 1646 2442 1649 2448
rect 1662 2441 1665 2468
rect 1686 2452 1689 2458
rect 1710 2442 1713 2658
rect 1718 2552 1721 2768
rect 1726 2692 1729 2808
rect 1734 2782 1737 2848
rect 1758 2802 1761 2868
rect 1774 2862 1777 2918
rect 1798 2902 1801 2918
rect 1822 2902 1825 2918
rect 1798 2872 1801 2878
rect 1782 2862 1785 2868
rect 1830 2852 1833 2859
rect 1778 2848 1782 2851
rect 1742 2772 1745 2798
rect 1758 2762 1761 2788
rect 1806 2752 1809 2818
rect 1750 2748 1769 2751
rect 1734 2742 1737 2748
rect 1750 2732 1753 2748
rect 1766 2742 1769 2748
rect 1758 2732 1761 2738
rect 1774 2722 1777 2748
rect 1734 2682 1737 2698
rect 1742 2651 1745 2718
rect 1782 2692 1785 2738
rect 1790 2692 1793 2748
rect 1802 2738 1806 2741
rect 1814 2692 1817 2798
rect 1822 2792 1825 2808
rect 1838 2792 1841 3058
rect 1854 3052 1857 3068
rect 1918 3062 1921 3068
rect 1866 3058 1870 3061
rect 1878 3052 1881 3058
rect 1894 3051 1897 3058
rect 1890 3048 1897 3051
rect 1902 3052 1905 3058
rect 1886 2952 1889 3028
rect 1910 2952 1913 2978
rect 1862 2892 1865 2938
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1885 2903 1888 2907
rect 1910 2902 1913 2948
rect 1942 2922 1945 2928
rect 1862 2862 1865 2888
rect 1894 2872 1897 2888
rect 1926 2791 1929 2818
rect 1934 2812 1937 2858
rect 1926 2788 1937 2791
rect 1830 2742 1833 2748
rect 1886 2742 1889 2748
rect 1750 2682 1753 2688
rect 1750 2668 1774 2671
rect 1750 2662 1753 2668
rect 1782 2662 1785 2678
rect 1794 2658 1798 2661
rect 1742 2648 1750 2651
rect 1718 2542 1721 2548
rect 1654 2438 1665 2441
rect 1482 2338 1489 2341
rect 1434 2268 1441 2271
rect 1438 2262 1441 2268
rect 1430 2252 1433 2258
rect 1406 2152 1409 2158
rect 1430 2152 1433 2218
rect 1446 2182 1449 2268
rect 1454 2262 1457 2298
rect 1474 2288 1478 2291
rect 1486 2282 1489 2338
rect 1582 2332 1585 2338
rect 1534 2322 1537 2328
rect 1502 2282 1505 2308
rect 1566 2292 1569 2328
rect 1598 2322 1601 2348
rect 1606 2332 1609 2358
rect 1634 2348 1638 2351
rect 1622 2342 1625 2348
rect 1634 2338 1638 2341
rect 1614 2331 1617 2338
rect 1646 2331 1649 2338
rect 1614 2328 1649 2331
rect 1614 2312 1617 2318
rect 1462 2262 1465 2268
rect 1478 2262 1481 2278
rect 1534 2272 1537 2278
rect 1562 2268 1566 2271
rect 1486 2221 1489 2258
rect 1482 2218 1489 2221
rect 1502 2212 1505 2268
rect 1518 2262 1521 2268
rect 1522 2258 1526 2261
rect 1558 2242 1561 2258
rect 1542 2222 1545 2238
rect 1570 2218 1574 2221
rect 1614 2192 1617 2308
rect 1654 2282 1657 2438
rect 1686 2392 1689 2438
rect 1710 2392 1713 2398
rect 1726 2362 1729 2648
rect 1758 2632 1761 2658
rect 1766 2632 1769 2658
rect 1750 2462 1753 2598
rect 1758 2592 1761 2628
rect 1806 2612 1809 2658
rect 1822 2652 1825 2678
rect 1838 2672 1841 2738
rect 1858 2728 1862 2731
rect 1902 2722 1905 2728
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1885 2703 1888 2707
rect 1934 2692 1937 2788
rect 1950 2752 1953 3108
rect 1998 3063 2001 3068
rect 1958 2992 1961 3018
rect 1966 2982 1969 3058
rect 1990 2992 1993 3018
rect 2006 2952 2009 2958
rect 2014 2952 2017 3108
rect 2030 3101 2033 3118
rect 2038 3112 2041 3148
rect 2030 3098 2041 3101
rect 2022 3091 2025 3098
rect 2022 3088 2033 3091
rect 2030 3082 2033 3088
rect 1970 2948 1974 2951
rect 1974 2872 1977 2948
rect 1998 2942 2001 2948
rect 1982 2922 1985 2928
rect 2022 2922 2025 2958
rect 2038 2951 2041 3098
rect 2054 3092 2057 3138
rect 2062 3092 2065 3148
rect 2070 3112 2073 3168
rect 2078 3162 2081 3168
rect 2098 3148 2102 3151
rect 2086 3142 2089 3148
rect 2118 3132 2121 3318
rect 2134 3282 2137 3288
rect 2142 3172 2145 3318
rect 2174 3312 2177 3458
rect 2182 3332 2185 3658
rect 2270 3632 2273 3748
rect 2318 3742 2321 3748
rect 2282 3738 2286 3741
rect 2326 3732 2329 3748
rect 2334 3742 2337 3758
rect 2342 3732 2345 3818
rect 2358 3781 2361 3858
rect 2370 3848 2374 3851
rect 2438 3832 2441 3878
rect 2446 3862 2449 3868
rect 2384 3803 2386 3807
rect 2390 3803 2393 3807
rect 2397 3803 2400 3807
rect 2350 3778 2361 3781
rect 2350 3732 2353 3778
rect 2358 3752 2361 3768
rect 2358 3742 2361 3748
rect 2366 3742 2369 3798
rect 2306 3728 2310 3731
rect 2278 3692 2281 3728
rect 2286 3692 2289 3718
rect 2294 3662 2297 3668
rect 2322 3658 2326 3661
rect 2230 3552 2233 3598
rect 2218 3548 2222 3551
rect 2190 3522 2193 3548
rect 2206 3542 2209 3548
rect 2238 3542 2241 3568
rect 2326 3562 2329 3588
rect 2250 3558 2254 3561
rect 2250 3548 2254 3551
rect 2266 3548 2270 3551
rect 2198 3482 2201 3538
rect 2214 3502 2217 3518
rect 2278 3512 2281 3558
rect 2306 3548 2310 3551
rect 2294 3502 2297 3548
rect 2334 3542 2337 3718
rect 2342 3602 2345 3718
rect 2374 3711 2377 3718
rect 2366 3708 2377 3711
rect 2350 3552 2353 3558
rect 2358 3552 2361 3608
rect 2302 3522 2305 3538
rect 2326 3532 2329 3540
rect 2334 3492 2337 3508
rect 2342 3492 2345 3548
rect 2358 3492 2361 3528
rect 2366 3492 2369 3708
rect 2374 3692 2377 3698
rect 2390 3652 2393 3778
rect 2470 3752 2473 3928
rect 2486 3892 2489 3958
rect 2502 3942 2505 3947
rect 2518 3932 2521 4268
rect 2526 4182 2529 4348
rect 2542 4272 2545 4368
rect 2558 4352 2561 4408
rect 2570 4378 2574 4381
rect 2582 4372 2585 4438
rect 2566 4352 2569 4368
rect 2550 4292 2553 4308
rect 2558 4292 2561 4348
rect 2566 4282 2569 4348
rect 2570 4258 2574 4261
rect 2534 4252 2537 4258
rect 2590 4232 2593 4408
rect 2606 4352 2609 4358
rect 2582 4212 2585 4218
rect 2550 4142 2553 4188
rect 2590 4152 2593 4228
rect 2598 4162 2601 4168
rect 2630 4151 2633 4458
rect 2662 4432 2665 4458
rect 2694 4442 2697 4618
rect 2702 4482 2705 4598
rect 2742 4532 2745 4588
rect 2758 4552 2761 4568
rect 2786 4558 2790 4561
rect 2766 4552 2769 4558
rect 2798 4552 2801 4558
rect 2778 4548 2782 4551
rect 2806 4542 2809 4658
rect 2838 4552 2841 4658
rect 2846 4652 2849 4658
rect 2854 4652 2857 4658
rect 2846 4552 2849 4628
rect 2814 4542 2817 4548
rect 2742 4522 2745 4528
rect 2714 4468 2718 4471
rect 2726 4471 2729 4488
rect 2738 4478 2742 4481
rect 2726 4468 2734 4471
rect 2702 4462 2705 4468
rect 2662 4372 2665 4418
rect 2686 4381 2689 4418
rect 2710 4392 2713 4468
rect 2750 4462 2753 4518
rect 2790 4470 2793 4508
rect 2798 4472 2801 4538
rect 2830 4502 2833 4518
rect 2810 4488 2814 4491
rect 2762 4448 2766 4451
rect 2734 4422 2737 4428
rect 2766 4422 2769 4448
rect 2678 4378 2689 4381
rect 2718 4382 2721 4418
rect 2670 4362 2673 4378
rect 2638 4351 2641 4358
rect 2638 4272 2641 4328
rect 2678 4292 2681 4378
rect 2686 4362 2689 4368
rect 2698 4358 2702 4361
rect 2718 4352 2721 4378
rect 2750 4352 2753 4418
rect 2758 4362 2761 4388
rect 2774 4372 2777 4418
rect 2798 4372 2801 4468
rect 2822 4462 2825 4488
rect 2834 4468 2838 4471
rect 2846 4462 2849 4488
rect 2854 4472 2857 4648
rect 2874 4558 2878 4561
rect 2910 4532 2913 4618
rect 2950 4612 2953 4658
rect 2954 4548 2958 4551
rect 2982 4542 2985 4678
rect 2994 4658 2998 4661
rect 3014 4552 3017 4628
rect 3030 4572 3033 4818
rect 3050 4758 3054 4761
rect 3046 4632 3049 4758
rect 3066 4748 3070 4751
rect 3066 4738 3070 4741
rect 3070 4662 3073 4668
rect 3046 4562 3049 4618
rect 3030 4542 3033 4548
rect 2866 4528 2870 4531
rect 3002 4528 3006 4531
rect 2888 4503 2890 4507
rect 2894 4503 2897 4507
rect 2901 4503 2904 4507
rect 2890 4488 2894 4491
rect 2910 4482 2913 4528
rect 3006 4492 3009 4518
rect 3046 4511 3049 4547
rect 3038 4508 3049 4511
rect 2834 4458 2838 4461
rect 2806 4432 2809 4448
rect 2738 4348 2742 4351
rect 2802 4348 2806 4351
rect 2694 4312 2697 4338
rect 2638 4192 2641 4258
rect 2662 4172 2665 4218
rect 2702 4212 2705 4348
rect 2710 4342 2713 4348
rect 2766 4342 2769 4348
rect 2722 4338 2726 4341
rect 2734 4322 2737 4338
rect 2758 4332 2761 4338
rect 2774 4322 2777 4348
rect 2710 4252 2713 4258
rect 2630 4148 2638 4151
rect 2642 4148 2646 4151
rect 2558 4132 2561 4148
rect 2614 4142 2617 4148
rect 2622 4142 2625 4148
rect 2526 4102 2529 4118
rect 2534 4112 2537 4128
rect 2630 4122 2633 4138
rect 2678 4122 2681 4148
rect 2694 4142 2697 4148
rect 2534 3962 2537 3968
rect 2550 3952 2553 4098
rect 2558 4072 2561 4088
rect 2566 4072 2569 4118
rect 2566 4061 2569 4068
rect 2558 4058 2569 4061
rect 2574 4062 2577 4118
rect 2598 4082 2601 4118
rect 2622 4072 2625 4098
rect 2630 4092 2633 4118
rect 2638 4092 2641 4118
rect 2686 4102 2689 4138
rect 2702 4072 2705 4208
rect 2718 4142 2721 4168
rect 2726 4142 2729 4308
rect 2770 4288 2774 4291
rect 2774 4272 2777 4278
rect 2750 4202 2753 4238
rect 2774 4232 2777 4258
rect 2782 4242 2785 4338
rect 2790 4292 2793 4348
rect 2814 4342 2817 4438
rect 2854 4392 2857 4468
rect 2878 4462 2881 4468
rect 2974 4462 2977 4468
rect 3022 4462 3025 4468
rect 2870 4382 2873 4458
rect 2834 4348 2838 4351
rect 2798 4332 2801 4338
rect 2822 4322 2825 4328
rect 2830 4322 2833 4328
rect 2802 4278 2806 4281
rect 2798 4232 2801 4268
rect 2814 4262 2817 4268
rect 2838 4252 2841 4278
rect 2814 4242 2817 4248
rect 2754 4168 2758 4171
rect 2742 4152 2745 4158
rect 2774 4152 2777 4178
rect 2786 4158 2790 4161
rect 2690 4068 2694 4071
rect 2586 4058 2590 4061
rect 2534 3942 2537 3948
rect 2558 3942 2561 4058
rect 2574 4052 2577 4058
rect 2598 4052 2601 4068
rect 2486 3852 2489 3878
rect 2502 3872 2505 3928
rect 2558 3922 2561 3938
rect 2566 3922 2569 3948
rect 2582 3942 2585 3978
rect 2622 3952 2625 3958
rect 2582 3932 2585 3938
rect 2566 3912 2569 3918
rect 2574 3902 2577 3918
rect 2510 3872 2513 3888
rect 2550 3862 2553 3878
rect 2574 3862 2577 3868
rect 2482 3838 2486 3841
rect 2502 3812 2505 3858
rect 2502 3762 2505 3798
rect 2566 3762 2569 3838
rect 2478 3752 2481 3758
rect 2506 3748 2510 3751
rect 2410 3728 2414 3731
rect 2422 3692 2425 3728
rect 2402 3688 2406 3691
rect 2430 3682 2433 3748
rect 2446 3742 2449 3748
rect 2558 3742 2561 3748
rect 2486 3732 2489 3738
rect 2494 3712 2497 3718
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2397 3603 2400 3607
rect 2374 3522 2377 3548
rect 2374 3492 2377 3518
rect 2398 3492 2401 3538
rect 2198 3462 2201 3478
rect 2214 3472 2217 3478
rect 2326 3472 2329 3478
rect 2342 3472 2345 3488
rect 2414 3482 2417 3668
rect 2446 3662 2449 3668
rect 2438 3652 2441 3658
rect 2422 3612 2425 3648
rect 2438 3552 2441 3628
rect 2454 3592 2457 3668
rect 2462 3662 2465 3698
rect 2494 3671 2497 3678
rect 2486 3668 2497 3671
rect 2486 3662 2489 3668
rect 2494 3652 2497 3658
rect 2478 3582 2481 3648
rect 2446 3522 2449 3538
rect 2350 3472 2353 3478
rect 2206 3462 2209 3468
rect 2286 3442 2289 3458
rect 2194 3438 2198 3441
rect 2246 3422 2249 3438
rect 2310 3422 2313 3468
rect 2246 3342 2249 3418
rect 2326 3402 2329 3468
rect 2346 3448 2350 3451
rect 2366 3412 2369 3448
rect 2258 3347 2262 3350
rect 2198 3322 2201 3338
rect 2202 3318 2206 3321
rect 2166 3152 2169 3298
rect 2182 3242 2185 3318
rect 2146 3148 2150 3151
rect 2050 3068 2054 3071
rect 2050 3058 2054 3061
rect 2062 3052 2065 3088
rect 2070 3072 2073 3108
rect 2070 3062 2073 3068
rect 2054 2962 2057 2968
rect 2034 2948 2041 2951
rect 2070 2942 2073 2998
rect 2078 2992 2081 3058
rect 2074 2938 2078 2941
rect 2086 2932 2089 3128
rect 2094 3082 2097 3118
rect 2126 3062 2129 3068
rect 2134 3062 2137 3108
rect 2146 3068 2150 3071
rect 2182 3062 2185 3088
rect 2114 3058 2118 3061
rect 2094 3022 2097 3058
rect 2134 3042 2137 3058
rect 2166 3042 2169 3048
rect 2106 3028 2110 3031
rect 2102 2952 2105 2958
rect 2066 2928 2070 2931
rect 1966 2752 1969 2868
rect 1998 2862 2001 2898
rect 2034 2888 2038 2891
rect 2038 2862 2041 2878
rect 2050 2868 2057 2871
rect 1974 2842 1977 2858
rect 2054 2852 2057 2868
rect 2070 2862 2073 2868
rect 2070 2852 2073 2858
rect 2078 2852 2081 2928
rect 2094 2892 2097 2918
rect 2086 2882 2089 2888
rect 1942 2732 1945 2748
rect 2006 2742 2009 2778
rect 2038 2762 2041 2768
rect 1998 2682 2001 2718
rect 1834 2668 1838 2671
rect 1862 2662 1865 2668
rect 1834 2658 1838 2661
rect 1822 2632 1825 2648
rect 1830 2602 1833 2658
rect 1870 2651 1873 2668
rect 1858 2648 1873 2651
rect 1878 2612 1881 2678
rect 2014 2672 2017 2748
rect 2030 2712 2033 2758
rect 2038 2742 2041 2748
rect 2046 2702 2049 2718
rect 2054 2682 2057 2848
rect 2062 2832 2065 2838
rect 2070 2751 2073 2838
rect 2094 2812 2097 2848
rect 2102 2802 2105 2888
rect 2110 2872 2113 2918
rect 2110 2852 2113 2858
rect 2118 2852 2121 2908
rect 2094 2761 2097 2798
rect 2118 2792 2121 2828
rect 2126 2781 2129 3018
rect 2142 2872 2145 2878
rect 2150 2872 2153 2888
rect 2158 2862 2161 3018
rect 2182 3002 2185 3058
rect 2174 2942 2177 2947
rect 2174 2902 2177 2928
rect 2174 2892 2177 2898
rect 2182 2882 2185 2888
rect 2138 2858 2142 2861
rect 2190 2852 2193 3318
rect 2246 3302 2249 3338
rect 2294 3322 2297 3328
rect 2234 3288 2238 3291
rect 2198 3263 2201 3288
rect 2214 3272 2217 3278
rect 2254 3272 2257 3288
rect 2262 3272 2265 3308
rect 2290 3288 2294 3291
rect 2246 3252 2249 3258
rect 2230 3232 2233 3248
rect 2230 3152 2233 3168
rect 2222 3142 2225 3148
rect 2198 3012 2201 3018
rect 2246 2992 2249 3248
rect 2262 3161 2265 3268
rect 2270 3262 2273 3288
rect 2286 3242 2289 3248
rect 2294 3222 2297 3268
rect 2302 3262 2305 3378
rect 2310 3342 2313 3348
rect 2318 3342 2321 3348
rect 2330 3338 2334 3341
rect 2302 3242 2305 3248
rect 2254 3158 2265 3161
rect 2254 3152 2257 3158
rect 2302 3152 2305 3168
rect 2310 3152 2313 3338
rect 2342 3312 2345 3348
rect 2334 3152 2337 3268
rect 2358 3162 2361 3258
rect 2374 3222 2377 3438
rect 2438 3422 2441 3458
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2397 3403 2400 3407
rect 2422 3352 2425 3398
rect 2398 3332 2401 3348
rect 2382 3262 2385 3288
rect 2390 3282 2393 3328
rect 2438 3302 2441 3418
rect 2446 3402 2449 3518
rect 2462 3462 2465 3488
rect 2502 3482 2505 3738
rect 2518 3672 2521 3708
rect 2526 3682 2529 3718
rect 2542 3702 2545 3728
rect 2550 3672 2553 3698
rect 2558 3682 2561 3738
rect 2566 3702 2569 3758
rect 2574 3752 2577 3848
rect 2582 3752 2585 3808
rect 2582 3742 2585 3748
rect 2590 3742 2593 3908
rect 2598 3862 2601 3938
rect 2638 3932 2641 4018
rect 2646 3952 2649 3968
rect 2582 3672 2585 3698
rect 2598 3672 2601 3738
rect 2606 3702 2609 3818
rect 2622 3792 2625 3888
rect 2638 3872 2641 3908
rect 2662 3892 2665 4058
rect 2694 4052 2697 4058
rect 2710 4051 2713 4140
rect 2726 4132 2729 4138
rect 2734 4122 2737 4148
rect 2750 4072 2753 4148
rect 2786 4138 2790 4141
rect 2722 4058 2726 4061
rect 2710 4048 2721 4051
rect 2694 3992 2697 4048
rect 2710 3962 2713 4018
rect 2694 3892 2697 3948
rect 2702 3922 2705 3928
rect 2646 3872 2649 3878
rect 2702 3872 2705 3918
rect 2666 3868 2670 3871
rect 2678 3862 2681 3868
rect 2666 3858 2670 3861
rect 2630 3842 2633 3848
rect 2626 3788 2633 3791
rect 2630 3762 2633 3788
rect 2630 3752 2633 3758
rect 2530 3648 2534 3651
rect 2526 3642 2529 3648
rect 2534 3592 2537 3598
rect 2510 3582 2513 3588
rect 2542 3572 2545 3658
rect 2574 3652 2577 3658
rect 2514 3548 2518 3551
rect 2550 3542 2553 3558
rect 2558 3551 2561 3618
rect 2574 3592 2577 3648
rect 2590 3632 2593 3668
rect 2622 3662 2625 3748
rect 2638 3742 2641 3858
rect 2646 3842 2649 3848
rect 2662 3752 2665 3858
rect 2710 3842 2713 3858
rect 2718 3822 2721 4048
rect 2734 4012 2737 4058
rect 2742 3912 2745 4048
rect 2750 3942 2753 3968
rect 2726 3892 2729 3908
rect 2742 3882 2745 3888
rect 2734 3872 2737 3878
rect 2694 3762 2697 3818
rect 2670 3752 2673 3758
rect 2702 3752 2705 3768
rect 2758 3762 2761 4118
rect 2766 4072 2769 4118
rect 2798 4112 2801 4228
rect 2854 4202 2857 4338
rect 2870 4332 2873 4378
rect 2958 4372 2961 4458
rect 2938 4348 2945 4351
rect 2894 4342 2897 4348
rect 2888 4303 2890 4307
rect 2894 4303 2897 4307
rect 2901 4303 2904 4307
rect 2934 4292 2937 4318
rect 2874 4278 2878 4281
rect 2918 4272 2921 4278
rect 2862 4212 2865 4258
rect 2870 4232 2873 4268
rect 2910 4242 2913 4258
rect 2926 4242 2929 4248
rect 2934 4242 2937 4248
rect 2818 4168 2822 4171
rect 2810 4158 2814 4161
rect 2854 4152 2857 4198
rect 2810 4148 2814 4151
rect 2814 4112 2817 4138
rect 2870 4132 2873 4228
rect 2878 4152 2881 4158
rect 2934 4152 2937 4218
rect 2942 4192 2945 4348
rect 2982 4332 2985 4378
rect 3014 4352 3017 4358
rect 3030 4352 3033 4508
rect 3038 4492 3041 4508
rect 3054 4462 3057 4648
rect 3078 4642 3081 4858
rect 3086 4652 3089 4858
rect 3150 4782 3153 4948
rect 3166 4942 3169 5018
rect 3206 5002 3209 5068
rect 3262 5062 3265 5068
rect 3366 5062 3369 5068
rect 3446 5062 3449 5068
rect 3470 5062 3473 5068
rect 3766 5063 3769 5068
rect 3538 5058 3542 5061
rect 3578 5058 3582 5061
rect 3946 5058 3950 5061
rect 3342 5052 3345 5058
rect 3214 5042 3217 5048
rect 3426 5038 3430 5041
rect 3194 4948 3198 4951
rect 3206 4942 3209 4998
rect 3166 4882 3169 4938
rect 3214 4872 3217 5008
rect 3230 4972 3233 4978
rect 3250 4968 3254 4971
rect 3262 4952 3265 5038
rect 3494 5012 3497 5058
rect 3400 5003 3402 5007
rect 3406 5003 3409 5007
rect 3413 5003 3416 5007
rect 3290 4968 3294 4971
rect 3302 4952 3305 4958
rect 3274 4948 3278 4951
rect 3262 4942 3265 4948
rect 3230 4901 3233 4928
rect 3222 4898 3233 4901
rect 3166 4863 3169 4868
rect 3198 4821 3201 4858
rect 3198 4818 3209 4821
rect 3094 4752 3097 4758
rect 3206 4752 3209 4818
rect 3102 4702 3105 4748
rect 3110 4692 3113 4718
rect 3150 4692 3153 4718
rect 3158 4692 3161 4738
rect 3174 4711 3177 4747
rect 3174 4708 3185 4711
rect 3182 4692 3185 4708
rect 3062 4482 3065 4558
rect 3094 4481 3097 4688
rect 3150 4682 3153 4688
rect 3146 4668 3150 4671
rect 3118 4662 3121 4668
rect 3102 4512 3105 4658
rect 3110 4642 3113 4658
rect 3158 4551 3161 4688
rect 3190 4662 3193 4668
rect 3154 4548 3161 4551
rect 3150 4542 3153 4548
rect 3110 4482 3113 4518
rect 3118 4482 3121 4518
rect 3094 4478 3102 4481
rect 3078 4472 3081 4478
rect 3098 4468 3102 4471
rect 3114 4468 3118 4471
rect 3134 4462 3137 4528
rect 3166 4502 3169 4658
rect 3198 4652 3201 4658
rect 3206 4652 3209 4708
rect 3198 4552 3201 4648
rect 3214 4552 3217 4868
rect 3222 4662 3225 4898
rect 3230 4882 3233 4888
rect 3246 4872 3249 4938
rect 3254 4872 3257 4938
rect 3278 4872 3281 4928
rect 3286 4892 3289 4948
rect 3310 4942 3313 4988
rect 3282 4868 3286 4871
rect 3246 4862 3249 4868
rect 3302 4862 3305 4868
rect 3274 4858 3278 4861
rect 3238 4682 3241 4718
rect 3230 4672 3233 4678
rect 3246 4662 3249 4858
rect 3262 4852 3265 4858
rect 3254 4662 3257 4668
rect 3262 4662 3265 4838
rect 3270 4742 3273 4828
rect 3302 4792 3305 4858
rect 3310 4832 3313 4938
rect 3318 4882 3321 4918
rect 3270 4732 3273 4738
rect 3286 4692 3289 4748
rect 3306 4747 3310 4750
rect 3302 4692 3305 4728
rect 3318 4691 3321 4878
rect 3326 4832 3329 4868
rect 3334 4862 3337 4958
rect 3350 4952 3353 4978
rect 3434 4968 3438 4971
rect 3370 4948 3374 4951
rect 3382 4862 3385 4938
rect 3414 4902 3417 4918
rect 3398 4862 3401 4868
rect 3438 4862 3441 4888
rect 3350 4842 3353 4848
rect 3374 4752 3377 4818
rect 3382 4772 3385 4858
rect 3400 4803 3402 4807
rect 3406 4803 3409 4807
rect 3413 4803 3416 4807
rect 3414 4751 3417 4758
rect 3362 4718 3366 4721
rect 3318 4688 3329 4691
rect 3326 4682 3329 4688
rect 3350 4682 3353 4718
rect 3318 4672 3321 4678
rect 3350 4672 3353 4678
rect 3270 4662 3273 4668
rect 3366 4662 3369 4678
rect 3378 4668 3382 4671
rect 3398 4662 3401 4688
rect 3422 4672 3425 4678
rect 3222 4562 3225 4618
rect 3254 4612 3257 4618
rect 3262 4582 3265 4658
rect 3330 4648 3334 4651
rect 3342 4622 3345 4658
rect 3382 4652 3385 4658
rect 3406 4642 3409 4668
rect 3362 4638 3366 4641
rect 3294 4562 3297 4568
rect 3322 4558 3326 4561
rect 3282 4548 3289 4551
rect 3182 4542 3185 4547
rect 3214 4512 3217 4548
rect 3222 4502 3225 4538
rect 3230 4532 3233 4538
rect 3246 4482 3249 4528
rect 3262 4522 3265 4538
rect 3270 4502 3273 4548
rect 3154 4478 3158 4481
rect 3178 4468 3182 4471
rect 3218 4468 3222 4471
rect 3150 4462 3153 4468
rect 3074 4458 3078 4461
rect 3122 4458 3126 4461
rect 3046 4402 3049 4458
rect 3054 4452 3057 4458
rect 3078 4442 3081 4448
rect 3070 4351 3073 4358
rect 2974 4282 2977 4318
rect 2982 4292 2985 4328
rect 3038 4322 3041 4348
rect 3054 4332 3057 4338
rect 2950 4252 2953 4258
rect 2974 4161 2977 4278
rect 2982 4272 2985 4278
rect 2990 4262 2993 4308
rect 3014 4272 3017 4278
rect 3006 4262 3009 4268
rect 3010 4248 3014 4251
rect 3022 4212 3025 4258
rect 3030 4252 3033 4258
rect 3038 4252 3041 4288
rect 3054 4272 3057 4328
rect 3070 4263 3073 4268
rect 2970 4158 2977 4161
rect 2982 4152 2985 4208
rect 3050 4188 3054 4191
rect 3022 4172 3025 4178
rect 3086 4162 3089 4398
rect 3094 4222 3097 4438
rect 3102 4342 3105 4418
rect 3134 4402 3137 4458
rect 3158 4451 3161 4468
rect 3194 4458 3198 4461
rect 3226 4458 3230 4461
rect 3206 4452 3209 4458
rect 3150 4448 3161 4451
rect 3178 4448 3190 4451
rect 3150 4392 3153 4448
rect 3222 4442 3225 4448
rect 3238 4432 3241 4458
rect 3254 4442 3257 4448
rect 3286 4442 3289 4548
rect 3358 4551 3361 4558
rect 3318 4542 3321 4548
rect 3342 4542 3345 4548
rect 3326 4532 3329 4538
rect 3334 4472 3337 4488
rect 3374 4472 3377 4518
rect 3382 4472 3385 4478
rect 3310 4462 3313 4468
rect 3350 4452 3353 4458
rect 3358 4452 3361 4458
rect 3366 4442 3369 4458
rect 3130 4378 3134 4381
rect 3150 4352 3153 4388
rect 3166 4362 3169 4418
rect 3138 4338 3142 4341
rect 3042 4158 3046 4161
rect 3022 4142 3025 4148
rect 3086 4142 3089 4148
rect 3102 4142 3105 4148
rect 3110 4142 3113 4158
rect 3118 4152 3121 4318
rect 3130 4288 3134 4291
rect 3150 4252 3153 4348
rect 3166 4282 3169 4318
rect 3174 4292 3177 4318
rect 3182 4262 3185 4268
rect 3166 4242 3169 4258
rect 3182 4182 3185 4248
rect 3150 4152 3153 4158
rect 3130 4148 3134 4151
rect 2774 4072 2777 4098
rect 2766 4052 2769 4058
rect 2774 4022 2777 4068
rect 2782 4062 2785 4068
rect 2798 4052 2801 4078
rect 2830 4072 2833 4088
rect 2822 4042 2825 4048
rect 2830 4032 2833 4058
rect 2846 3972 2849 4068
rect 2862 4052 2865 4059
rect 2870 4052 2873 4128
rect 2888 4103 2890 4107
rect 2894 4103 2897 4107
rect 2901 4103 2904 4107
rect 2918 4092 2921 4138
rect 2930 4088 2934 4091
rect 2926 4082 2929 4088
rect 2894 4062 2897 4068
rect 2946 4058 2950 4061
rect 2826 3958 2830 3961
rect 2862 3961 2865 4028
rect 2894 3992 2897 4048
rect 2942 3972 2945 3978
rect 2858 3958 2865 3961
rect 2766 3951 2769 3958
rect 2810 3948 2814 3951
rect 2850 3948 2854 3951
rect 2742 3752 2745 3758
rect 2766 3752 2769 3788
rect 2782 3752 2785 3948
rect 2838 3942 2841 3948
rect 2798 3932 2801 3938
rect 2862 3921 2865 3958
rect 2922 3948 2926 3951
rect 2878 3942 2881 3948
rect 2966 3942 2969 4058
rect 2990 4022 2993 4138
rect 2998 4092 3001 4128
rect 3022 4112 3025 4138
rect 3078 4132 3081 4138
rect 3118 4092 3121 4148
rect 3154 4138 3158 4141
rect 3190 4122 3193 4428
rect 3330 4347 3334 4350
rect 3202 4268 3206 4271
rect 3214 4152 3217 4338
rect 3238 4322 3241 4347
rect 3350 4342 3353 4348
rect 3254 4332 3257 4338
rect 3274 4318 3278 4321
rect 3254 4292 3257 4318
rect 3222 4282 3225 4288
rect 3222 4262 3225 4278
rect 3262 4262 3265 4268
rect 3270 4262 3273 4268
rect 3234 4258 3238 4261
rect 3238 4142 3241 4148
rect 3246 4142 3249 4248
rect 3286 4221 3289 4318
rect 3302 4282 3305 4338
rect 3366 4322 3369 4358
rect 3374 4352 3377 4468
rect 3382 4452 3385 4458
rect 3390 4452 3393 4618
rect 3400 4603 3402 4607
rect 3406 4603 3409 4607
rect 3413 4603 3416 4607
rect 3418 4568 3422 4571
rect 3398 4462 3401 4508
rect 3406 4472 3409 4528
rect 3422 4472 3425 4548
rect 3410 4468 3414 4471
rect 3382 4372 3385 4378
rect 3390 4361 3393 4438
rect 3398 4432 3401 4458
rect 3400 4403 3402 4407
rect 3406 4403 3409 4407
rect 3413 4403 3416 4407
rect 3382 4358 3393 4361
rect 3414 4362 3417 4368
rect 3382 4352 3385 4358
rect 3402 4348 3406 4351
rect 3390 4342 3393 4348
rect 3314 4258 3318 4261
rect 3286 4218 3297 4221
rect 3278 4152 3281 4218
rect 3006 4062 3009 4078
rect 3118 4072 3121 4078
rect 3190 4072 3193 4118
rect 3018 4068 3022 4071
rect 3050 4068 3054 4071
rect 3094 4062 3097 4068
rect 3102 4062 3105 4068
rect 3022 4052 3025 4058
rect 3070 4052 3073 4058
rect 3038 4012 3041 4018
rect 3006 3952 3009 3978
rect 3046 3942 3049 3968
rect 3070 3962 3073 4048
rect 3134 4042 3137 4059
rect 3094 4032 3097 4038
rect 3118 3992 3121 4018
rect 3098 3978 3102 3981
rect 3070 3952 3073 3958
rect 3090 3948 3094 3951
rect 3130 3948 3134 3951
rect 3142 3942 3145 3978
rect 3150 3962 3153 4038
rect 3198 3961 3201 4098
rect 3206 3992 3209 4108
rect 3222 4072 3225 4078
rect 3230 4062 3233 4078
rect 3218 4058 3222 4061
rect 3222 3982 3225 3988
rect 3218 3978 3222 3981
rect 3190 3958 3201 3961
rect 3150 3952 3153 3958
rect 3182 3952 3185 3958
rect 3162 3948 3166 3951
rect 3190 3942 3193 3958
rect 2870 3932 2873 3938
rect 2862 3918 2873 3921
rect 2822 3872 2825 3888
rect 2838 3872 2841 3878
rect 2846 3872 2849 3878
rect 2806 3852 2809 3859
rect 2802 3768 2806 3771
rect 2822 3762 2825 3768
rect 2694 3742 2697 3748
rect 2726 3742 2729 3748
rect 2690 3738 2694 3741
rect 2706 3738 2710 3741
rect 2654 3702 2657 3718
rect 2662 3692 2665 3728
rect 2710 3711 2713 3718
rect 2710 3708 2718 3711
rect 2650 3688 2657 3691
rect 2630 3662 2633 3688
rect 2654 3682 2657 3688
rect 2694 3672 2697 3708
rect 2598 3582 2601 3658
rect 2638 3642 2641 3658
rect 2650 3648 2654 3651
rect 2558 3548 2566 3551
rect 2574 3542 2577 3558
rect 2582 3542 2585 3578
rect 2606 3562 2609 3628
rect 2594 3558 2598 3561
rect 2590 3521 2593 3548
rect 2614 3542 2617 3618
rect 2638 3572 2641 3638
rect 2662 3632 2665 3648
rect 2678 3592 2681 3658
rect 2686 3602 2689 3668
rect 2706 3658 2710 3661
rect 2714 3658 2718 3661
rect 2702 3642 2705 3648
rect 2718 3632 2721 3648
rect 2686 3562 2689 3568
rect 2642 3558 2646 3561
rect 2650 3548 2654 3551
rect 2590 3518 2601 3521
rect 2518 3482 2521 3488
rect 2534 3472 2537 3518
rect 2562 3458 2566 3461
rect 2502 3442 2505 3458
rect 2510 3412 2513 3458
rect 2474 3348 2478 3351
rect 2486 3342 2489 3348
rect 2466 3338 2470 3341
rect 2462 3292 2465 3308
rect 2438 3272 2441 3278
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2397 3203 2400 3207
rect 2262 3142 2265 3148
rect 2262 3062 2265 3138
rect 2270 3042 2273 3148
rect 2278 3142 2281 3148
rect 2314 3138 2326 3141
rect 2330 3138 2334 3141
rect 2342 3131 2345 3158
rect 2406 3142 2409 3268
rect 2470 3262 2473 3268
rect 2478 3262 2481 3338
rect 2498 3328 2502 3331
rect 2510 3292 2513 3298
rect 2494 3282 2497 3288
rect 2518 3262 2521 3348
rect 2550 3342 2553 3448
rect 2582 3422 2585 3458
rect 2582 3352 2585 3418
rect 2330 3128 2345 3131
rect 2294 3122 2297 3128
rect 2322 3118 2326 3121
rect 2286 3102 2289 3118
rect 2294 3072 2297 3078
rect 2310 3072 2313 3088
rect 2342 3072 2345 3078
rect 2278 3052 2281 3059
rect 2270 3002 2273 3038
rect 2238 2952 2241 2988
rect 2246 2952 2249 2978
rect 2302 2952 2305 3038
rect 2210 2948 2214 2951
rect 2258 2948 2262 2951
rect 2210 2938 2214 2941
rect 2270 2892 2273 2918
rect 2214 2862 2217 2888
rect 2278 2872 2281 2878
rect 2178 2848 2182 2851
rect 2118 2778 2129 2781
rect 2094 2758 2105 2761
rect 2066 2748 2073 2751
rect 2094 2742 2097 2748
rect 2070 2732 2073 2738
rect 2042 2678 2046 2681
rect 1898 2558 1902 2561
rect 1766 2552 1769 2558
rect 1766 2501 1769 2548
rect 1778 2528 1782 2531
rect 1758 2498 1769 2501
rect 1758 2472 1761 2498
rect 1774 2482 1777 2518
rect 1798 2492 1801 2548
rect 1786 2468 1790 2471
rect 1814 2462 1817 2468
rect 1786 2458 1790 2461
rect 1738 2418 1742 2421
rect 1774 2412 1777 2418
rect 1746 2358 1750 2361
rect 1662 2342 1665 2358
rect 1670 2352 1673 2358
rect 1766 2352 1769 2398
rect 1806 2392 1809 2448
rect 1822 2412 1825 2548
rect 1910 2542 1913 2668
rect 1926 2663 1929 2668
rect 1998 2662 2001 2668
rect 2030 2662 2033 2678
rect 2058 2658 2062 2661
rect 1918 2572 1921 2618
rect 1990 2612 1993 2618
rect 1926 2552 1929 2608
rect 2022 2592 2025 2658
rect 1974 2551 1977 2558
rect 2046 2552 2049 2658
rect 2070 2652 2073 2678
rect 2078 2662 2081 2718
rect 2078 2642 2081 2648
rect 2086 2642 2089 2728
rect 2102 2672 2105 2758
rect 2118 2742 2121 2778
rect 2126 2752 2129 2768
rect 2134 2752 2137 2838
rect 2214 2821 2217 2858
rect 2246 2852 2249 2859
rect 2206 2818 2217 2821
rect 2158 2772 2161 2818
rect 2206 2792 2209 2818
rect 2214 2812 2217 2818
rect 2146 2768 2150 2771
rect 2174 2762 2177 2768
rect 2146 2748 2150 2751
rect 2138 2738 2142 2741
rect 2110 2672 2113 2678
rect 2142 2672 2145 2718
rect 2166 2682 2169 2758
rect 2194 2738 2198 2741
rect 2178 2718 2182 2721
rect 2190 2692 2193 2708
rect 2182 2682 2185 2688
rect 2206 2672 2209 2768
rect 2214 2672 2217 2798
rect 2286 2772 2289 2928
rect 2302 2902 2305 2948
rect 2318 2932 2321 2958
rect 2334 2952 2337 2988
rect 2342 2952 2345 2958
rect 2350 2952 2353 3008
rect 2294 2852 2297 2868
rect 2270 2752 2273 2758
rect 2294 2752 2297 2758
rect 2130 2668 2134 2671
rect 2094 2662 2097 2668
rect 2114 2658 2118 2661
rect 2150 2658 2158 2661
rect 2226 2658 2230 2661
rect 2150 2652 2153 2658
rect 2162 2648 2166 2651
rect 2094 2602 2097 2618
rect 2070 2562 2073 2598
rect 2126 2592 2129 2628
rect 2134 2622 2137 2648
rect 2002 2548 2006 2551
rect 1834 2538 1838 2541
rect 1918 2532 1921 2538
rect 1942 2532 1945 2538
rect 1894 2522 1897 2528
rect 1830 2482 1833 2518
rect 1894 2512 1897 2518
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1885 2503 1888 2507
rect 1882 2468 1886 2471
rect 1850 2458 1854 2461
rect 1830 2402 1833 2458
rect 1838 2442 1841 2448
rect 1862 2422 1865 2468
rect 1890 2458 1894 2461
rect 1854 2412 1857 2418
rect 1778 2358 1782 2361
rect 1798 2352 1801 2358
rect 1830 2352 1833 2398
rect 1886 2362 1889 2368
rect 1714 2348 1718 2351
rect 1754 2348 1758 2351
rect 1786 2348 1790 2351
rect 1842 2348 1846 2351
rect 1882 2348 1886 2351
rect 1678 2322 1681 2348
rect 1702 2332 1705 2338
rect 1758 2332 1761 2348
rect 1798 2342 1801 2348
rect 1894 2342 1897 2418
rect 1834 2338 1838 2341
rect 1766 2332 1769 2338
rect 1694 2322 1697 2328
rect 1750 2322 1753 2328
rect 1662 2312 1665 2318
rect 1734 2292 1737 2298
rect 1630 2262 1633 2278
rect 1654 2272 1657 2278
rect 1674 2268 1678 2271
rect 1698 2268 1702 2271
rect 1682 2258 1694 2261
rect 1678 2242 1681 2258
rect 1726 2252 1729 2268
rect 1742 2262 1745 2318
rect 1774 2272 1777 2278
rect 1758 2262 1761 2268
rect 1790 2263 1793 2298
rect 1746 2258 1750 2261
rect 1822 2262 1825 2328
rect 1902 2322 1905 2528
rect 1918 2482 1921 2508
rect 1914 2448 1918 2451
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1885 2303 1888 2307
rect 1862 2272 1865 2278
rect 1682 2218 1686 2221
rect 1678 2192 1681 2208
rect 1694 2192 1697 2248
rect 1354 2148 1358 2151
rect 1394 2148 1398 2151
rect 1366 2142 1369 2148
rect 1414 2142 1417 2148
rect 1374 2132 1377 2138
rect 1334 2082 1337 2088
rect 1330 2068 1334 2071
rect 1358 2062 1361 2108
rect 1390 2092 1393 2118
rect 1366 2082 1369 2088
rect 1398 2082 1401 2128
rect 1422 2092 1425 2148
rect 1438 2092 1441 2158
rect 1478 2152 1481 2168
rect 1454 2142 1457 2148
rect 1454 2072 1457 2108
rect 1402 2068 1406 2071
rect 1442 2068 1446 2071
rect 1466 2068 1473 2071
rect 1366 2062 1369 2068
rect 1378 2058 1382 2061
rect 1426 2058 1430 2061
rect 1206 1992 1209 2018
rect 1158 1972 1161 1988
rect 1158 1962 1161 1968
rect 1214 1962 1217 1978
rect 1126 1872 1129 1878
rect 1150 1862 1153 1898
rect 1158 1862 1161 1868
rect 1130 1858 1134 1861
rect 1130 1848 1134 1851
rect 1094 1802 1097 1848
rect 1106 1768 1110 1771
rect 1086 1752 1089 1758
rect 1094 1742 1097 1748
rect 1074 1738 1078 1741
rect 974 1702 977 1738
rect 990 1732 993 1738
rect 1014 1692 1017 1698
rect 1110 1682 1113 1768
rect 1142 1752 1145 1808
rect 1174 1802 1177 1948
rect 1190 1942 1193 1948
rect 1198 1942 1201 1948
rect 1214 1942 1217 1948
rect 1246 1942 1249 1947
rect 1182 1932 1185 1938
rect 1246 1911 1249 1928
rect 1238 1908 1249 1911
rect 1190 1822 1193 1868
rect 1202 1858 1206 1861
rect 1238 1842 1241 1908
rect 1262 1872 1265 1948
rect 1278 1922 1281 2058
rect 1294 2032 1297 2058
rect 1358 2042 1361 2058
rect 1352 2003 1354 2007
rect 1358 2003 1361 2007
rect 1365 2003 1368 2007
rect 1338 1978 1342 1981
rect 1318 1952 1321 1958
rect 1374 1952 1377 1958
rect 1334 1922 1337 1948
rect 1346 1938 1350 1941
rect 1390 1941 1393 2038
rect 1406 2032 1409 2048
rect 1422 2012 1425 2028
rect 1422 1972 1425 2008
rect 1398 1952 1401 1968
rect 1422 1962 1425 1968
rect 1438 1962 1441 2048
rect 1446 2042 1449 2068
rect 1462 1992 1465 2058
rect 1470 2002 1473 2068
rect 1486 2052 1489 2178
rect 1554 2168 1558 2171
rect 1682 2168 1686 2171
rect 1566 2162 1569 2168
rect 1590 2152 1593 2168
rect 1702 2162 1705 2168
rect 1710 2162 1713 2218
rect 1694 2152 1697 2158
rect 1726 2152 1729 2178
rect 1734 2161 1737 2198
rect 1742 2182 1745 2258
rect 1746 2168 1750 2171
rect 1734 2158 1745 2161
rect 1554 2148 1558 2151
rect 1570 2148 1574 2151
rect 1642 2148 1646 2151
rect 1606 2142 1609 2148
rect 1734 2142 1737 2148
rect 1538 2138 1542 2141
rect 1574 2122 1577 2138
rect 1602 2128 1606 2131
rect 1658 2128 1662 2131
rect 1538 2118 1542 2121
rect 1598 2092 1601 2108
rect 1582 2082 1585 2088
rect 1606 2082 1609 2098
rect 1630 2082 1633 2128
rect 1654 2082 1657 2118
rect 1610 2078 1614 2081
rect 1626 2078 1630 2081
rect 1494 2072 1497 2078
rect 1558 2072 1561 2078
rect 1646 2072 1649 2078
rect 1566 2062 1569 2068
rect 1514 2058 1518 2061
rect 1554 2058 1558 2061
rect 1574 2052 1577 2068
rect 1630 2062 1633 2068
rect 1654 2062 1657 2078
rect 1670 2062 1673 2128
rect 1710 2092 1713 2128
rect 1718 2111 1721 2138
rect 1718 2108 1726 2111
rect 1734 2102 1737 2138
rect 1598 2058 1606 2061
rect 1666 2058 1670 2061
rect 1518 2002 1521 2018
rect 1534 2012 1537 2048
rect 1410 1958 1417 1961
rect 1414 1952 1417 1958
rect 1390 1938 1398 1941
rect 1270 1862 1273 1878
rect 1278 1862 1281 1868
rect 1310 1862 1313 1918
rect 1366 1902 1369 1938
rect 1398 1931 1401 1938
rect 1398 1928 1409 1931
rect 1358 1892 1361 1898
rect 1318 1872 1321 1878
rect 1294 1842 1297 1848
rect 1258 1838 1262 1841
rect 1238 1822 1241 1838
rect 1158 1752 1161 1798
rect 1130 1748 1134 1751
rect 1158 1742 1161 1748
rect 1174 1742 1177 1748
rect 1182 1742 1185 1768
rect 1138 1738 1142 1741
rect 1190 1731 1193 1818
rect 1206 1752 1209 1768
rect 1238 1742 1241 1818
rect 1310 1802 1313 1858
rect 1326 1852 1329 1868
rect 1334 1862 1337 1868
rect 1350 1852 1353 1878
rect 1374 1852 1377 1868
rect 1390 1862 1393 1918
rect 1266 1748 1270 1751
rect 1182 1728 1193 1731
rect 1222 1732 1225 1738
rect 1182 1682 1185 1728
rect 1138 1678 1142 1681
rect 1046 1662 1049 1668
rect 1078 1663 1081 1668
rect 1110 1662 1113 1668
rect 1126 1662 1129 1668
rect 1006 1642 1009 1648
rect 1110 1641 1113 1648
rect 1102 1638 1113 1641
rect 1014 1582 1017 1618
rect 1054 1602 1057 1628
rect 1046 1552 1049 1568
rect 1054 1552 1057 1598
rect 1102 1592 1105 1638
rect 1126 1598 1134 1601
rect 1126 1592 1129 1598
rect 1086 1572 1089 1578
rect 1134 1572 1137 1578
rect 1118 1562 1121 1568
rect 1018 1548 1022 1551
rect 1098 1548 1102 1551
rect 982 1542 985 1548
rect 990 1542 993 1548
rect 1078 1542 1081 1548
rect 978 1458 982 1461
rect 1006 1442 1009 1448
rect 1014 1442 1017 1538
rect 1030 1422 1033 1518
rect 1102 1512 1105 1548
rect 1114 1538 1118 1541
rect 1126 1492 1129 1548
rect 1142 1522 1145 1668
rect 1190 1662 1193 1718
rect 1254 1682 1257 1728
rect 1286 1692 1289 1778
rect 1334 1771 1337 1818
rect 1342 1812 1345 1838
rect 1350 1832 1353 1848
rect 1352 1803 1354 1807
rect 1358 1803 1361 1807
rect 1365 1803 1368 1807
rect 1334 1768 1345 1771
rect 1318 1758 1334 1761
rect 1318 1752 1321 1758
rect 1330 1748 1334 1751
rect 1330 1738 1334 1741
rect 1318 1722 1321 1728
rect 1330 1688 1334 1691
rect 1298 1678 1302 1681
rect 1274 1668 1278 1671
rect 1330 1668 1334 1671
rect 1266 1658 1270 1661
rect 1150 1571 1153 1618
rect 1278 1612 1281 1658
rect 1302 1622 1305 1668
rect 1342 1662 1345 1768
rect 1374 1732 1377 1758
rect 1398 1752 1401 1918
rect 1406 1862 1409 1928
rect 1422 1922 1425 1948
rect 1434 1938 1438 1941
rect 1406 1852 1409 1858
rect 1422 1832 1425 1858
rect 1430 1762 1433 1868
rect 1426 1748 1430 1751
rect 1402 1738 1406 1741
rect 1422 1732 1425 1738
rect 1366 1672 1369 1678
rect 1358 1662 1361 1668
rect 1374 1662 1377 1728
rect 1406 1712 1409 1728
rect 1434 1718 1441 1721
rect 1414 1702 1417 1718
rect 1406 1672 1409 1678
rect 1390 1662 1393 1668
rect 1310 1652 1313 1658
rect 1166 1572 1169 1578
rect 1150 1568 1161 1571
rect 1150 1532 1153 1558
rect 1158 1542 1161 1568
rect 1182 1552 1185 1588
rect 1342 1572 1345 1618
rect 1390 1612 1393 1658
rect 1414 1652 1417 1698
rect 1438 1682 1441 1718
rect 1422 1672 1425 1678
rect 1426 1658 1430 1661
rect 1352 1603 1354 1607
rect 1358 1603 1361 1607
rect 1365 1603 1368 1607
rect 1406 1592 1409 1598
rect 1314 1558 1318 1561
rect 1358 1552 1361 1558
rect 1170 1548 1174 1551
rect 1338 1548 1342 1551
rect 1246 1542 1249 1548
rect 1170 1538 1174 1541
rect 1094 1472 1097 1478
rect 1046 1462 1049 1468
rect 1102 1462 1105 1468
rect 1066 1458 1070 1461
rect 1114 1458 1118 1461
rect 1054 1442 1057 1458
rect 1142 1452 1145 1468
rect 1170 1458 1174 1461
rect 1078 1442 1081 1448
rect 1126 1432 1129 1448
rect 1078 1392 1081 1408
rect 946 1348 950 1351
rect 974 1342 977 1348
rect 954 1338 958 1341
rect 918 1328 929 1331
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 861 1303 864 1307
rect 882 1288 886 1291
rect 870 1272 873 1288
rect 890 1268 894 1271
rect 906 1268 910 1271
rect 822 1262 825 1268
rect 778 1258 782 1261
rect 842 1258 846 1261
rect 638 1192 641 1228
rect 646 1222 649 1228
rect 646 1152 649 1218
rect 578 1148 582 1151
rect 634 1148 638 1151
rect 582 1132 585 1138
rect 422 942 425 948
rect 426 938 433 941
rect 398 852 401 858
rect 406 772 409 908
rect 422 862 425 878
rect 430 852 433 938
rect 462 932 465 948
rect 486 912 489 938
rect 510 932 513 948
rect 446 872 449 908
rect 486 882 489 888
rect 462 862 465 868
rect 470 852 473 858
rect 354 748 358 751
rect 366 712 369 748
rect 374 742 377 748
rect 386 718 390 721
rect 366 672 369 698
rect 362 658 366 661
rect 374 652 377 678
rect 390 672 393 678
rect 390 652 393 658
rect 334 622 337 638
rect 328 603 330 607
rect 334 603 337 607
rect 341 603 344 607
rect 358 582 361 618
rect 306 548 310 551
rect 338 548 342 551
rect 354 548 358 551
rect 398 551 401 568
rect 306 538 310 541
rect 382 532 385 538
rect 166 462 169 478
rect 174 462 177 468
rect 246 462 249 498
rect 326 492 329 498
rect 306 488 310 491
rect 342 482 345 488
rect 322 468 326 471
rect 374 462 377 468
rect 306 458 310 461
rect 62 392 65 458
rect 150 452 153 458
rect 198 452 201 458
rect 126 418 134 421
rect 126 352 129 418
rect 182 392 185 448
rect 382 442 385 468
rect 198 392 201 428
rect 328 403 330 407
rect 334 403 337 407
rect 341 403 344 407
rect 210 358 214 361
rect 350 352 353 368
rect 330 348 334 351
rect 86 342 89 348
rect 206 342 209 348
rect 66 338 70 341
rect 194 338 198 341
rect 70 272 73 308
rect 94 262 97 308
rect 110 282 113 298
rect 142 263 145 268
rect 10 138 14 141
rect 54 112 57 258
rect 62 252 65 258
rect 86 152 89 218
rect 150 172 153 268
rect 102 151 105 158
rect 150 142 153 168
rect 10 88 14 91
rect 62 72 65 118
rect 70 63 73 78
rect 86 72 89 138
rect 102 82 105 88
rect 126 72 129 78
rect 118 62 121 68
rect 150 62 153 68
rect 158 62 161 278
rect 166 192 169 298
rect 190 292 193 338
rect 210 288 214 291
rect 222 272 225 348
rect 246 281 249 338
rect 254 322 257 348
rect 310 342 313 348
rect 362 338 366 341
rect 242 278 249 281
rect 214 252 217 258
rect 206 152 209 188
rect 166 62 169 148
rect 182 132 185 138
rect 222 102 225 268
rect 254 262 257 268
rect 238 192 241 218
rect 262 192 265 328
rect 294 272 297 338
rect 314 328 318 331
rect 358 312 361 338
rect 366 322 369 328
rect 302 262 305 278
rect 366 272 369 308
rect 382 292 385 328
rect 282 258 286 261
rect 270 172 273 218
rect 294 151 297 168
rect 318 152 321 268
rect 342 262 345 268
rect 390 262 393 408
rect 398 352 401 458
rect 406 452 409 768
rect 414 752 417 778
rect 422 752 425 838
rect 494 832 497 858
rect 486 752 489 808
rect 502 792 505 848
rect 518 792 521 858
rect 506 758 510 761
rect 450 748 454 751
rect 466 748 470 751
rect 422 742 425 748
rect 526 742 529 938
rect 542 862 545 868
rect 550 862 553 948
rect 558 892 561 1098
rect 594 1088 598 1091
rect 646 1082 649 1088
rect 610 1068 614 1071
rect 630 1062 633 1068
rect 618 1058 622 1061
rect 598 1052 601 1058
rect 566 972 569 978
rect 574 952 577 1048
rect 630 992 633 1058
rect 646 982 649 1058
rect 654 1052 657 1148
rect 662 1131 665 1248
rect 726 1231 729 1238
rect 726 1228 737 1231
rect 722 1158 726 1161
rect 670 1142 673 1158
rect 722 1148 726 1151
rect 662 1128 673 1131
rect 670 1092 673 1128
rect 678 1082 681 1148
rect 698 1138 702 1141
rect 694 1122 697 1128
rect 678 1072 681 1078
rect 662 1052 665 1068
rect 686 1052 689 1088
rect 702 1072 705 1108
rect 602 948 606 951
rect 574 912 577 948
rect 582 942 585 948
rect 646 932 649 978
rect 654 952 657 958
rect 594 928 598 931
rect 626 928 630 931
rect 586 868 590 871
rect 578 858 582 861
rect 554 848 558 851
rect 534 791 537 818
rect 598 791 601 878
rect 606 872 609 898
rect 610 868 614 871
rect 618 858 622 861
rect 630 852 633 898
rect 638 872 641 918
rect 630 802 633 848
rect 614 792 617 798
rect 534 788 545 791
rect 598 788 606 791
rect 542 751 545 788
rect 570 748 574 751
rect 422 462 425 738
rect 462 732 465 738
rect 470 722 473 728
rect 430 662 433 718
rect 478 712 481 728
rect 486 702 489 738
rect 494 692 497 718
rect 482 688 486 691
rect 446 662 449 678
rect 510 662 513 708
rect 534 672 537 678
rect 446 472 449 658
rect 490 648 494 651
rect 458 588 462 591
rect 486 462 489 608
rect 494 592 497 638
rect 518 612 521 668
rect 558 662 561 698
rect 610 688 614 691
rect 622 662 625 768
rect 646 762 649 888
rect 654 862 657 908
rect 662 902 665 928
rect 662 872 665 878
rect 670 871 673 988
rect 686 972 689 978
rect 702 962 705 1038
rect 718 992 721 1138
rect 734 1082 737 1228
rect 758 1152 761 1258
rect 806 1192 809 1258
rect 902 1252 905 1258
rect 918 1252 921 1328
rect 926 1292 929 1308
rect 954 1268 958 1271
rect 942 1262 945 1268
rect 966 1262 969 1268
rect 894 1248 902 1251
rect 886 1222 889 1248
rect 814 1172 817 1218
rect 830 1202 833 1218
rect 838 1192 841 1208
rect 822 1152 825 1158
rect 810 1148 814 1151
rect 758 1142 761 1148
rect 782 1132 785 1148
rect 742 1062 745 1118
rect 774 1102 777 1128
rect 798 1092 801 1098
rect 814 1092 817 1128
rect 814 1072 817 1088
rect 798 992 801 1038
rect 814 992 817 1028
rect 682 948 686 951
rect 734 951 737 958
rect 694 941 697 948
rect 686 938 697 941
rect 686 892 689 938
rect 718 892 721 938
rect 714 878 718 881
rect 670 868 678 871
rect 678 862 681 868
rect 658 858 665 861
rect 646 752 649 758
rect 654 752 657 818
rect 662 782 665 858
rect 706 858 710 861
rect 670 852 673 858
rect 710 752 713 818
rect 710 732 713 738
rect 638 692 641 698
rect 718 692 721 848
rect 750 792 753 988
rect 814 952 817 958
rect 766 882 769 928
rect 782 862 785 878
rect 758 842 761 858
rect 726 722 729 728
rect 734 692 737 758
rect 754 748 758 751
rect 766 742 769 748
rect 774 742 777 748
rect 754 738 758 741
rect 782 732 785 858
rect 798 832 801 858
rect 798 752 801 828
rect 806 741 809 938
rect 822 902 825 1148
rect 830 1142 833 1168
rect 842 1148 846 1151
rect 854 1141 857 1158
rect 838 1138 857 1141
rect 878 1142 881 1188
rect 830 1062 833 1068
rect 838 1022 841 1138
rect 886 1132 889 1148
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 861 1103 864 1107
rect 834 958 838 961
rect 848 903 850 907
rect 854 903 857 907
rect 861 903 864 907
rect 814 862 817 888
rect 826 868 830 871
rect 822 802 825 858
rect 862 852 865 858
rect 830 842 833 848
rect 846 792 849 838
rect 870 762 873 938
rect 878 882 881 1068
rect 894 1012 897 1248
rect 926 1212 929 1248
rect 950 1222 953 1258
rect 918 1172 921 1178
rect 902 1162 905 1168
rect 910 1142 913 1158
rect 922 1148 926 1151
rect 942 1132 945 1158
rect 902 1062 905 1118
rect 942 1092 945 1128
rect 958 1092 961 1208
rect 966 1152 969 1258
rect 974 1152 977 1318
rect 982 1312 985 1348
rect 1014 1342 1017 1368
rect 982 1292 985 1298
rect 990 1282 993 1318
rect 982 1212 985 1248
rect 994 1218 998 1221
rect 982 1092 985 1158
rect 990 1152 993 1218
rect 998 1132 1001 1148
rect 1006 1132 1009 1340
rect 1022 1292 1025 1358
rect 1014 1262 1017 1268
rect 1014 1192 1017 1208
rect 1022 1172 1025 1238
rect 1030 1152 1033 1388
rect 1102 1372 1105 1398
rect 1114 1388 1118 1391
rect 1038 1362 1041 1368
rect 1046 1352 1049 1358
rect 1086 1352 1089 1368
rect 1054 1342 1057 1348
rect 1042 1338 1046 1341
rect 1038 1272 1041 1328
rect 1062 1322 1065 1348
rect 1118 1342 1121 1368
rect 1134 1362 1137 1418
rect 1150 1362 1153 1388
rect 1158 1362 1161 1388
rect 1134 1352 1137 1358
rect 1142 1352 1145 1358
rect 1174 1352 1177 1378
rect 1206 1362 1209 1538
rect 1214 1442 1217 1498
rect 1222 1452 1225 1538
rect 1246 1462 1249 1468
rect 1286 1462 1289 1548
rect 1326 1542 1329 1548
rect 1294 1482 1297 1528
rect 1266 1458 1270 1461
rect 1254 1452 1257 1458
rect 1294 1452 1297 1478
rect 1310 1472 1313 1488
rect 1330 1468 1334 1471
rect 1330 1458 1334 1461
rect 1234 1448 1238 1451
rect 1198 1352 1201 1358
rect 1222 1352 1225 1448
rect 1230 1392 1233 1408
rect 1254 1352 1257 1438
rect 1298 1428 1302 1431
rect 1318 1392 1321 1458
rect 1350 1452 1353 1458
rect 1366 1452 1369 1548
rect 1390 1492 1393 1558
rect 1398 1482 1401 1578
rect 1406 1552 1409 1558
rect 1414 1542 1417 1558
rect 1338 1428 1342 1431
rect 1352 1403 1354 1407
rect 1358 1403 1361 1407
rect 1365 1403 1368 1407
rect 1346 1388 1350 1391
rect 1318 1372 1321 1388
rect 1374 1382 1377 1458
rect 1162 1348 1166 1351
rect 1238 1342 1241 1348
rect 1246 1342 1249 1348
rect 1306 1338 1310 1341
rect 1118 1332 1121 1338
rect 1126 1321 1129 1338
rect 1286 1332 1289 1338
rect 1118 1318 1129 1321
rect 1046 1272 1049 1278
rect 1046 1192 1049 1268
rect 1054 1222 1057 1258
rect 1070 1252 1073 1298
rect 1098 1268 1102 1271
rect 1086 1262 1089 1268
rect 1046 1162 1049 1188
rect 1062 1152 1065 1218
rect 1094 1202 1097 1258
rect 1102 1192 1105 1268
rect 1118 1232 1121 1318
rect 1198 1302 1201 1328
rect 1270 1312 1273 1318
rect 1198 1292 1201 1298
rect 1302 1272 1305 1328
rect 1334 1322 1337 1348
rect 1138 1259 1142 1262
rect 1214 1262 1217 1268
rect 1310 1262 1313 1308
rect 1318 1262 1321 1268
rect 1350 1262 1353 1318
rect 1358 1282 1361 1338
rect 1382 1302 1385 1468
rect 1390 1282 1393 1298
rect 1398 1282 1401 1388
rect 1406 1312 1409 1458
rect 1422 1392 1425 1658
rect 1446 1592 1449 1958
rect 1454 1942 1457 1968
rect 1526 1951 1529 1978
rect 1558 1962 1561 1968
rect 1566 1952 1569 1978
rect 1574 1952 1577 2048
rect 1598 1992 1601 2058
rect 1686 2032 1689 2038
rect 1582 1952 1585 1988
rect 1614 1972 1617 2028
rect 1694 2012 1697 2058
rect 1726 2042 1729 2048
rect 1614 1962 1617 1968
rect 1726 1952 1729 1998
rect 1742 1952 1745 2158
rect 1758 1992 1761 2248
rect 1798 2112 1801 2148
rect 1822 2142 1825 2258
rect 1862 2242 1865 2268
rect 1894 2262 1897 2308
rect 1910 2292 1913 2338
rect 1926 2291 1929 2528
rect 1934 2471 1937 2518
rect 1934 2468 1945 2471
rect 1942 2462 1945 2468
rect 1934 2452 1937 2458
rect 1966 2442 1969 2448
rect 1966 2362 1969 2398
rect 1934 2352 1937 2358
rect 1918 2288 1929 2291
rect 1934 2292 1937 2318
rect 1958 2292 1961 2358
rect 1974 2342 1977 2528
rect 2014 2492 2017 2498
rect 1998 2482 2001 2488
rect 2038 2482 2041 2518
rect 2046 2492 2049 2538
rect 1986 2468 1990 2471
rect 2018 2468 2022 2471
rect 2030 2462 2033 2468
rect 2062 2462 2065 2488
rect 2054 2452 2057 2458
rect 2054 2422 2057 2448
rect 1982 2351 1985 2398
rect 2022 2392 2025 2398
rect 2070 2362 2073 2558
rect 2086 2542 2089 2558
rect 2110 2552 2113 2558
rect 2182 2552 2185 2658
rect 2238 2652 2241 2748
rect 2278 2742 2281 2748
rect 2310 2742 2313 2808
rect 2318 2791 2321 2918
rect 2326 2902 2329 2938
rect 2334 2861 2337 2948
rect 2342 2942 2345 2948
rect 2350 2892 2353 2908
rect 2330 2858 2337 2861
rect 2342 2862 2345 2878
rect 2342 2832 2345 2848
rect 2318 2788 2329 2791
rect 2326 2751 2329 2788
rect 2266 2738 2270 2741
rect 2246 2672 2249 2698
rect 2286 2671 2289 2738
rect 2282 2668 2289 2671
rect 2274 2658 2281 2661
rect 2190 2632 2193 2648
rect 2238 2612 2241 2648
rect 2138 2548 2142 2551
rect 2102 2522 2105 2528
rect 2126 2522 2129 2528
rect 2094 2512 2097 2518
rect 2094 2492 2097 2498
rect 2190 2492 2193 2608
rect 2238 2592 2241 2598
rect 2254 2572 2257 2618
rect 2078 2362 2081 2478
rect 2118 2472 2121 2478
rect 2102 2452 2105 2468
rect 2114 2458 2118 2461
rect 2146 2458 2153 2461
rect 2162 2458 2166 2461
rect 2126 2452 2129 2458
rect 2134 2442 2137 2458
rect 2142 2442 2145 2448
rect 2150 2441 2153 2458
rect 2178 2448 2182 2451
rect 2150 2438 2158 2441
rect 2170 2418 2174 2421
rect 2118 2392 2121 2408
rect 2022 2352 2025 2358
rect 2046 2352 2049 2358
rect 1974 2332 1977 2338
rect 1974 2322 1977 2328
rect 1910 2282 1913 2288
rect 1918 2282 1921 2288
rect 1966 2282 1969 2288
rect 1990 2282 1993 2288
rect 1894 2202 1897 2258
rect 1910 2172 1913 2258
rect 1838 2162 1841 2168
rect 1890 2158 1894 2161
rect 1846 2152 1849 2158
rect 1910 2152 1913 2158
rect 1858 2148 1862 2151
rect 1886 2132 1889 2148
rect 1902 2142 1905 2148
rect 1626 1948 1630 1951
rect 1706 1948 1710 1951
rect 1746 1948 1753 1951
rect 1582 1942 1585 1948
rect 1462 1822 1465 1868
rect 1470 1862 1473 1918
rect 1510 1842 1513 1938
rect 1590 1931 1593 1938
rect 1582 1928 1593 1931
rect 1598 1932 1601 1948
rect 1526 1892 1529 1898
rect 1542 1892 1545 1928
rect 1554 1878 1558 1881
rect 1570 1878 1574 1881
rect 1582 1871 1585 1928
rect 1574 1868 1585 1871
rect 1606 1872 1609 1948
rect 1654 1942 1657 1948
rect 1626 1938 1630 1941
rect 1670 1932 1673 1948
rect 1694 1942 1697 1948
rect 1706 1938 1710 1941
rect 1730 1938 1734 1941
rect 1698 1928 1702 1931
rect 1638 1922 1641 1928
rect 1670 1902 1673 1928
rect 1714 1918 1718 1921
rect 1714 1888 1718 1891
rect 1614 1882 1617 1888
rect 1558 1862 1561 1868
rect 1574 1862 1577 1868
rect 1530 1858 1534 1861
rect 1586 1858 1590 1861
rect 1462 1752 1465 1818
rect 1542 1792 1545 1858
rect 1558 1772 1561 1858
rect 1606 1852 1609 1858
rect 1590 1792 1593 1838
rect 1478 1692 1481 1748
rect 1510 1672 1513 1758
rect 1490 1668 1494 1671
rect 1462 1662 1465 1668
rect 1510 1662 1513 1668
rect 1494 1652 1497 1658
rect 1462 1552 1465 1558
rect 1478 1552 1481 1558
rect 1430 1432 1433 1548
rect 1454 1532 1457 1548
rect 1466 1538 1470 1541
rect 1486 1492 1489 1608
rect 1494 1562 1497 1568
rect 1506 1558 1510 1561
rect 1518 1542 1521 1698
rect 1526 1612 1529 1758
rect 1558 1752 1561 1758
rect 1546 1748 1550 1751
rect 1546 1738 1550 1741
rect 1578 1738 1582 1741
rect 1550 1562 1553 1598
rect 1558 1572 1561 1718
rect 1578 1668 1582 1671
rect 1578 1659 1582 1662
rect 1574 1562 1577 1568
rect 1538 1548 1545 1551
rect 1578 1548 1582 1551
rect 1530 1538 1534 1541
rect 1494 1532 1497 1538
rect 1518 1532 1521 1538
rect 1478 1482 1481 1488
rect 1510 1481 1513 1518
rect 1542 1512 1545 1548
rect 1614 1542 1617 1818
rect 1622 1742 1625 1878
rect 1726 1872 1729 1878
rect 1666 1858 1670 1861
rect 1678 1822 1681 1868
rect 1742 1862 1745 1868
rect 1714 1848 1718 1851
rect 1654 1742 1657 1748
rect 1622 1702 1625 1738
rect 1630 1712 1633 1718
rect 1670 1682 1673 1808
rect 1694 1762 1697 1848
rect 1750 1842 1753 1948
rect 1714 1758 1718 1761
rect 1726 1752 1729 1768
rect 1734 1752 1737 1768
rect 1754 1758 1758 1761
rect 1710 1742 1713 1748
rect 1766 1742 1769 2078
rect 1774 1981 1777 2068
rect 1790 2063 1793 2088
rect 1806 2072 1809 2128
rect 1838 2062 1841 2128
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1885 2103 1888 2107
rect 1858 2088 1862 2091
rect 1874 2068 1878 2071
rect 1890 2068 1894 2071
rect 1846 2062 1849 2068
rect 1902 2062 1905 2098
rect 1910 2092 1913 2138
rect 1918 2082 1921 2268
rect 1926 2202 1929 2278
rect 1938 2258 1942 2261
rect 1926 2142 1929 2198
rect 1950 2192 1953 2258
rect 1958 2192 1961 2268
rect 1974 2262 1977 2278
rect 2002 2268 2006 2271
rect 1990 2212 1993 2258
rect 1974 2162 1977 2188
rect 1958 2152 1961 2158
rect 1982 2152 1985 2168
rect 1934 2112 1937 2148
rect 1954 2138 1958 2141
rect 1942 2132 1945 2138
rect 1966 2092 1969 2098
rect 1926 2071 1929 2078
rect 1922 2068 1929 2071
rect 1966 2062 1969 2088
rect 1974 2072 1977 2108
rect 1982 2082 1985 2108
rect 1978 2068 1982 2071
rect 1838 2052 1841 2058
rect 1826 2048 1830 2051
rect 1854 2042 1857 2048
rect 1842 2038 1846 2041
rect 1786 1988 1790 1991
rect 1774 1978 1785 1981
rect 1774 1962 1777 1968
rect 1774 1902 1777 1958
rect 1774 1862 1777 1868
rect 1782 1752 1785 1978
rect 1790 1882 1793 1938
rect 1798 1932 1801 1968
rect 1814 1952 1817 2028
rect 1854 1988 1862 1991
rect 1826 1968 1830 1971
rect 1838 1962 1841 1988
rect 1854 1952 1857 1988
rect 1870 1972 1873 2058
rect 1918 2052 1921 2058
rect 1942 2052 1945 2058
rect 1926 2042 1929 2048
rect 1950 2042 1953 2048
rect 1982 2042 1985 2048
rect 1970 2038 1974 2041
rect 1902 1961 1905 1988
rect 1902 1958 1910 1961
rect 1870 1952 1873 1958
rect 1814 1822 1817 1838
rect 1798 1772 1801 1818
rect 1798 1752 1801 1758
rect 1714 1738 1718 1741
rect 1678 1732 1681 1738
rect 1742 1721 1745 1738
rect 1738 1718 1745 1721
rect 1686 1692 1689 1708
rect 1658 1668 1662 1671
rect 1670 1662 1673 1678
rect 1634 1658 1638 1661
rect 1622 1652 1625 1658
rect 1646 1562 1649 1658
rect 1662 1572 1665 1658
rect 1682 1648 1686 1651
rect 1694 1641 1697 1648
rect 1686 1638 1697 1641
rect 1702 1642 1705 1718
rect 1710 1662 1713 1688
rect 1718 1672 1721 1688
rect 1714 1648 1718 1651
rect 1686 1612 1689 1638
rect 1678 1592 1681 1598
rect 1694 1592 1697 1608
rect 1622 1552 1625 1558
rect 1662 1542 1665 1568
rect 1510 1478 1521 1481
rect 1438 1432 1441 1458
rect 1446 1452 1449 1458
rect 1454 1452 1457 1458
rect 1430 1392 1433 1418
rect 1462 1412 1465 1468
rect 1502 1462 1505 1468
rect 1510 1392 1513 1468
rect 1486 1351 1489 1388
rect 1422 1342 1425 1348
rect 1470 1342 1473 1348
rect 1518 1342 1521 1478
rect 1526 1412 1529 1458
rect 1534 1402 1537 1418
rect 1422 1328 1430 1331
rect 1414 1292 1417 1308
rect 1358 1272 1361 1278
rect 1242 1258 1246 1261
rect 1302 1258 1310 1261
rect 1094 1162 1097 1168
rect 1070 1152 1073 1158
rect 1022 1092 1025 1148
rect 1062 1122 1065 1148
rect 1102 1142 1105 1148
rect 1074 1138 1078 1141
rect 1118 1132 1121 1168
rect 1150 1151 1153 1158
rect 1166 1142 1169 1258
rect 1294 1242 1297 1248
rect 1218 1168 1222 1171
rect 1086 1082 1089 1098
rect 966 1072 969 1078
rect 990 1072 993 1078
rect 1006 1071 1009 1078
rect 1002 1068 1009 1071
rect 1038 1062 1041 1078
rect 1062 1062 1065 1078
rect 1102 1072 1105 1078
rect 1070 1062 1073 1068
rect 1010 1058 1014 1061
rect 1042 1058 1046 1061
rect 1030 1052 1033 1058
rect 966 1042 969 1048
rect 1022 1041 1025 1048
rect 1022 1038 1033 1041
rect 918 952 921 1018
rect 950 1002 953 1038
rect 998 992 1001 1038
rect 1030 992 1033 1038
rect 1050 1028 1054 1031
rect 958 962 961 968
rect 906 948 910 951
rect 886 922 889 948
rect 930 938 934 941
rect 898 928 902 931
rect 942 931 945 958
rect 974 952 977 958
rect 982 952 985 968
rect 1026 958 1030 961
rect 1062 952 1065 1058
rect 1118 1032 1121 1059
rect 962 948 966 951
rect 962 938 966 941
rect 934 928 945 931
rect 886 862 889 898
rect 894 872 897 918
rect 918 882 921 898
rect 926 862 929 928
rect 934 892 937 928
rect 958 872 961 878
rect 938 868 942 871
rect 902 852 905 858
rect 902 812 905 848
rect 914 828 918 831
rect 854 752 857 758
rect 818 748 822 751
rect 798 738 809 741
rect 670 682 673 688
rect 630 662 633 668
rect 650 658 654 661
rect 542 592 545 608
rect 538 558 542 561
rect 498 548 502 551
rect 582 551 585 578
rect 502 482 505 528
rect 518 492 521 538
rect 542 472 545 498
rect 550 482 553 528
rect 566 522 569 538
rect 566 472 569 518
rect 494 462 497 468
rect 518 462 521 468
rect 530 458 534 461
rect 406 372 409 448
rect 406 352 409 358
rect 398 342 401 348
rect 402 288 406 291
rect 414 262 417 378
rect 438 332 441 368
rect 454 362 457 458
rect 478 391 481 418
rect 478 388 489 391
rect 486 351 489 388
rect 454 342 457 348
rect 422 272 425 318
rect 438 292 441 328
rect 438 262 441 268
rect 446 262 449 278
rect 454 272 457 338
rect 470 292 473 348
rect 486 312 489 328
rect 502 282 505 318
rect 486 262 489 268
rect 328 203 330 207
rect 334 203 337 207
rect 341 203 344 207
rect 390 192 393 258
rect 414 252 417 258
rect 454 252 457 258
rect 174 72 177 98
rect 190 62 193 68
rect 198 62 201 98
rect 214 82 217 88
rect 230 72 233 138
rect 278 72 281 138
rect 306 88 310 91
rect 342 72 345 168
rect 430 162 433 218
rect 394 148 398 151
rect 434 148 438 151
rect 406 142 409 148
rect 450 138 454 141
rect 130 58 134 61
rect 414 62 417 118
rect 446 102 449 128
rect 422 92 425 98
rect 454 82 457 118
rect 462 62 465 158
rect 518 152 521 268
rect 534 192 537 258
rect 542 171 545 468
rect 550 452 553 458
rect 550 392 553 398
rect 566 342 569 468
rect 586 459 590 462
rect 582 342 585 347
rect 566 272 569 278
rect 606 262 609 278
rect 614 262 617 628
rect 630 502 633 658
rect 646 622 649 638
rect 646 592 649 618
rect 662 592 665 648
rect 670 562 673 668
rect 678 642 681 678
rect 726 672 729 688
rect 758 682 761 728
rect 706 658 710 661
rect 714 648 718 651
rect 666 558 670 561
rect 734 552 737 678
rect 758 672 761 678
rect 782 662 785 718
rect 742 612 745 648
rect 798 632 801 738
rect 818 728 822 731
rect 830 712 833 748
rect 806 592 809 708
rect 838 692 841 728
rect 848 703 850 707
rect 854 703 857 707
rect 861 703 864 707
rect 878 692 881 718
rect 878 682 881 688
rect 886 672 889 738
rect 878 668 886 671
rect 866 658 870 661
rect 770 578 774 581
rect 646 492 649 528
rect 654 481 657 538
rect 662 492 665 548
rect 646 478 657 481
rect 646 392 649 478
rect 686 472 689 498
rect 694 492 697 508
rect 702 482 705 518
rect 710 512 713 548
rect 734 472 737 548
rect 766 492 769 568
rect 818 558 822 561
rect 838 552 841 628
rect 846 552 849 608
rect 854 562 857 568
rect 862 552 865 618
rect 870 572 873 578
rect 794 548 798 551
rect 806 542 809 548
rect 794 538 798 541
rect 786 518 790 521
rect 674 468 678 471
rect 682 458 686 461
rect 654 372 657 438
rect 678 382 681 458
rect 702 352 705 468
rect 742 462 745 488
rect 774 472 777 478
rect 722 458 729 461
rect 726 382 729 458
rect 766 458 774 461
rect 742 452 745 458
rect 750 452 753 458
rect 766 442 769 458
rect 758 392 761 438
rect 766 392 769 438
rect 746 388 750 391
rect 750 372 753 378
rect 710 342 713 348
rect 638 262 641 328
rect 646 312 649 318
rect 662 282 665 338
rect 758 332 761 388
rect 798 362 801 518
rect 814 462 817 478
rect 806 392 809 418
rect 822 362 825 458
rect 830 442 833 538
rect 848 503 850 507
rect 854 503 857 507
rect 861 503 864 507
rect 850 488 854 491
rect 878 432 881 668
rect 886 542 889 648
rect 894 562 897 568
rect 902 552 905 638
rect 910 592 913 808
rect 926 732 929 838
rect 942 792 945 858
rect 974 792 977 918
rect 982 862 985 888
rect 922 558 926 561
rect 890 538 894 541
rect 890 468 894 471
rect 902 402 905 538
rect 934 532 937 758
rect 942 692 945 718
rect 958 692 961 758
rect 982 752 985 798
rect 998 752 1001 758
rect 1006 752 1009 948
rect 1038 942 1041 948
rect 1046 942 1049 948
rect 1038 892 1041 938
rect 1046 902 1049 938
rect 1046 872 1049 878
rect 1046 782 1049 868
rect 1054 862 1057 948
rect 1078 942 1081 958
rect 1094 952 1097 988
rect 1118 952 1121 958
rect 1130 948 1134 951
rect 1070 892 1073 918
rect 1094 862 1097 948
rect 1102 942 1105 948
rect 1102 872 1105 938
rect 1110 931 1113 938
rect 1110 928 1118 931
rect 1142 881 1145 958
rect 1134 878 1145 881
rect 1118 872 1121 878
rect 1058 858 1062 861
rect 1094 852 1097 858
rect 1078 832 1081 848
rect 982 732 985 738
rect 990 732 993 738
rect 970 668 974 671
rect 1014 662 1017 778
rect 1002 658 1006 661
rect 946 548 950 551
rect 958 532 961 638
rect 1014 632 1017 658
rect 982 552 985 568
rect 974 542 977 548
rect 934 492 937 528
rect 910 463 913 478
rect 942 462 945 498
rect 966 482 969 518
rect 982 462 985 468
rect 942 452 945 458
rect 950 452 953 458
rect 942 422 945 438
rect 934 392 937 398
rect 746 288 750 291
rect 662 272 665 278
rect 770 268 774 271
rect 562 258 569 261
rect 566 192 569 258
rect 614 251 617 258
rect 606 248 617 251
rect 638 252 641 258
rect 598 222 601 238
rect 590 218 598 221
rect 542 168 553 171
rect 550 152 553 168
rect 570 148 574 151
rect 518 122 521 148
rect 542 132 545 148
rect 550 142 553 148
rect 590 132 593 218
rect 606 192 609 248
rect 630 152 633 218
rect 526 91 529 128
rect 542 112 545 128
rect 598 122 601 128
rect 610 118 614 121
rect 522 88 529 91
rect 550 82 553 118
rect 558 62 561 78
rect 646 62 649 248
rect 666 148 670 151
rect 678 142 681 268
rect 686 262 689 268
rect 798 262 801 358
rect 838 352 841 388
rect 910 362 913 368
rect 942 352 945 418
rect 958 392 961 418
rect 814 342 817 348
rect 990 342 993 618
rect 1022 582 1025 758
rect 1038 742 1041 758
rect 1054 752 1057 818
rect 1074 747 1078 750
rect 1054 722 1057 738
rect 1082 688 1086 691
rect 1094 682 1097 848
rect 1118 772 1121 838
rect 1134 832 1137 878
rect 1150 872 1153 1128
rect 1182 1092 1185 1098
rect 1198 1072 1201 1168
rect 1290 1158 1294 1161
rect 1222 1152 1225 1158
rect 1222 1142 1225 1148
rect 1222 1062 1225 1068
rect 1190 992 1193 1028
rect 1238 1002 1241 1118
rect 1254 1112 1257 1158
rect 1302 1152 1305 1258
rect 1338 1248 1342 1251
rect 1350 1232 1353 1258
rect 1358 1252 1361 1258
rect 1352 1203 1354 1207
rect 1358 1203 1361 1207
rect 1365 1203 1368 1207
rect 1330 1188 1334 1191
rect 1310 1152 1313 1188
rect 1318 1152 1321 1158
rect 1350 1152 1353 1168
rect 1270 1132 1273 1138
rect 1294 1122 1297 1148
rect 1306 1138 1313 1141
rect 1266 1038 1270 1041
rect 1278 992 1281 1108
rect 1310 1062 1313 1138
rect 1318 1072 1321 1078
rect 1334 1062 1337 1148
rect 1298 1058 1302 1061
rect 1310 1052 1313 1058
rect 1290 1048 1294 1051
rect 1158 942 1161 968
rect 1166 952 1169 958
rect 1174 952 1177 958
rect 1222 952 1225 988
rect 1238 962 1241 988
rect 1254 958 1262 961
rect 1198 922 1201 948
rect 1206 938 1214 941
rect 1218 938 1222 941
rect 1198 882 1201 888
rect 1206 872 1209 938
rect 1246 932 1249 938
rect 1142 862 1145 868
rect 1214 852 1217 858
rect 1134 792 1137 828
rect 1058 668 1062 671
rect 1046 662 1049 668
rect 1058 658 1062 661
rect 998 452 1001 518
rect 1006 492 1009 578
rect 1014 552 1017 558
rect 1038 552 1041 618
rect 1070 592 1073 678
rect 1118 662 1121 768
rect 1146 758 1150 761
rect 1166 752 1169 828
rect 1222 792 1225 898
rect 1230 852 1233 888
rect 1242 868 1246 871
rect 1254 862 1257 958
rect 1262 952 1265 958
rect 1270 942 1273 948
rect 1270 872 1273 888
rect 1262 862 1265 868
rect 1286 852 1289 1008
rect 1334 952 1337 1058
rect 1318 942 1321 948
rect 1334 892 1337 938
rect 1238 822 1241 848
rect 1190 762 1193 778
rect 1190 752 1193 758
rect 1198 752 1201 758
rect 1206 732 1209 758
rect 1238 752 1241 818
rect 1246 792 1249 848
rect 1226 748 1230 751
rect 1262 742 1265 778
rect 1278 761 1281 818
rect 1286 782 1289 848
rect 1302 842 1305 868
rect 1326 862 1329 878
rect 1334 872 1337 888
rect 1342 861 1345 1148
rect 1374 1142 1377 1198
rect 1382 1192 1385 1268
rect 1390 1152 1393 1278
rect 1406 1272 1409 1278
rect 1398 1262 1401 1268
rect 1414 1262 1417 1268
rect 1402 1158 1406 1161
rect 1414 1152 1417 1228
rect 1406 1142 1409 1148
rect 1422 1082 1425 1328
rect 1526 1282 1529 1288
rect 1542 1281 1545 1508
rect 1550 1462 1553 1468
rect 1558 1462 1561 1538
rect 1582 1522 1585 1538
rect 1594 1488 1598 1491
rect 1622 1482 1625 1538
rect 1702 1502 1705 1638
rect 1726 1602 1729 1678
rect 1734 1612 1737 1718
rect 1750 1682 1753 1718
rect 1766 1682 1769 1688
rect 1782 1662 1785 1748
rect 1814 1742 1817 1818
rect 1838 1802 1841 1938
rect 1854 1872 1857 1948
rect 1870 1932 1873 1948
rect 1886 1942 1889 1958
rect 1934 1952 1937 2028
rect 1942 1952 1945 2008
rect 1990 1992 1993 2178
rect 1998 2092 2001 2258
rect 2006 2222 2009 2268
rect 2014 2052 2017 2338
rect 2038 2272 2041 2318
rect 2022 2262 2025 2268
rect 2022 2242 2025 2248
rect 2030 2132 2033 2148
rect 2038 2142 2041 2268
rect 2054 2263 2057 2268
rect 2038 2072 2041 2138
rect 2062 2062 2065 2348
rect 2078 2342 2081 2348
rect 2070 2322 2073 2338
rect 2070 2252 2073 2318
rect 2074 2248 2081 2251
rect 2078 2072 2081 2248
rect 2102 2242 2105 2318
rect 2110 2291 2113 2358
rect 2118 2348 2126 2351
rect 2118 2302 2121 2348
rect 2134 2342 2137 2378
rect 2158 2362 2161 2398
rect 2166 2392 2169 2398
rect 2138 2338 2145 2341
rect 2126 2332 2129 2338
rect 2142 2292 2145 2338
rect 2166 2332 2169 2368
rect 2182 2351 2185 2378
rect 2190 2362 2193 2418
rect 2198 2392 2201 2568
rect 2250 2548 2254 2551
rect 2262 2551 2265 2658
rect 2278 2592 2281 2658
rect 2298 2658 2305 2661
rect 2286 2652 2289 2658
rect 2258 2548 2265 2551
rect 2290 2568 2294 2571
rect 2214 2542 2217 2548
rect 2222 2542 2225 2548
rect 2206 2532 2209 2538
rect 2270 2532 2273 2568
rect 2218 2458 2222 2461
rect 2182 2348 2190 2351
rect 2198 2342 2201 2388
rect 2178 2338 2182 2341
rect 2110 2288 2118 2291
rect 2118 2192 2121 2278
rect 2150 2262 2153 2308
rect 2158 2292 2161 2318
rect 2174 2292 2177 2298
rect 2130 2258 2134 2261
rect 2150 2192 2153 2248
rect 2086 2112 2089 2118
rect 2082 2058 2086 2061
rect 2030 2042 2033 2058
rect 1894 1942 1897 1948
rect 1974 1942 1977 1948
rect 1898 1928 1902 1931
rect 1922 1928 1926 1931
rect 1954 1928 1958 1931
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1885 1903 1888 1907
rect 1926 1902 1929 1918
rect 1990 1882 1993 1948
rect 1998 1942 2001 1968
rect 2006 1952 2009 2008
rect 2030 1992 2033 2028
rect 2066 1968 2070 1971
rect 2078 1962 2081 1968
rect 2054 1952 2057 1958
rect 2082 1948 2086 1951
rect 2014 1942 2017 1948
rect 1850 1858 1854 1861
rect 1830 1742 1833 1747
rect 1794 1738 1798 1741
rect 1806 1662 1809 1688
rect 1814 1672 1817 1738
rect 1558 1432 1561 1448
rect 1566 1432 1569 1468
rect 1574 1462 1577 1468
rect 1630 1462 1633 1468
rect 1590 1432 1593 1448
rect 1558 1421 1561 1428
rect 1558 1418 1569 1421
rect 1566 1392 1569 1418
rect 1638 1392 1641 1498
rect 1690 1488 1694 1491
rect 1694 1472 1697 1478
rect 1710 1472 1713 1578
rect 1718 1562 1721 1568
rect 1734 1562 1737 1568
rect 1722 1548 1726 1551
rect 1742 1542 1745 1658
rect 1750 1602 1753 1658
rect 1762 1648 1766 1651
rect 1718 1532 1721 1538
rect 1734 1522 1737 1528
rect 1750 1502 1753 1548
rect 1758 1492 1761 1608
rect 1782 1562 1785 1568
rect 1798 1562 1801 1598
rect 1770 1558 1774 1561
rect 1766 1542 1769 1548
rect 1774 1532 1777 1538
rect 1782 1512 1785 1548
rect 1726 1472 1729 1478
rect 1738 1468 1742 1471
rect 1754 1468 1761 1471
rect 1702 1451 1705 1458
rect 1698 1448 1705 1451
rect 1630 1372 1633 1388
rect 1602 1358 1606 1361
rect 1618 1358 1622 1361
rect 1582 1352 1585 1358
rect 1686 1352 1689 1358
rect 1598 1342 1601 1348
rect 1614 1342 1617 1348
rect 1638 1342 1641 1348
rect 1702 1342 1705 1348
rect 1718 1342 1721 1347
rect 1570 1338 1574 1341
rect 1658 1338 1662 1341
rect 1582 1292 1585 1328
rect 1606 1312 1609 1338
rect 1614 1322 1617 1338
rect 1650 1328 1654 1331
rect 1538 1278 1545 1281
rect 1430 1252 1433 1258
rect 1430 1152 1433 1158
rect 1366 1072 1369 1078
rect 1386 1068 1390 1071
rect 1352 1003 1354 1007
rect 1358 1003 1361 1007
rect 1365 1003 1368 1007
rect 1334 858 1345 861
rect 1374 942 1377 1058
rect 1390 1052 1393 1058
rect 1406 1042 1409 1068
rect 1422 1063 1425 1068
rect 1430 1052 1433 1118
rect 1278 758 1286 761
rect 1294 752 1297 788
rect 1326 762 1329 768
rect 1334 752 1337 858
rect 1374 832 1377 938
rect 1406 882 1409 1008
rect 1414 952 1417 958
rect 1422 952 1425 988
rect 1430 952 1433 1038
rect 1430 942 1433 948
rect 1422 872 1425 878
rect 1352 803 1354 807
rect 1358 803 1361 807
rect 1365 803 1368 807
rect 1386 788 1390 791
rect 1406 752 1409 798
rect 1414 752 1417 858
rect 1422 752 1425 758
rect 1230 732 1233 738
rect 1142 692 1145 728
rect 1174 672 1177 718
rect 1182 692 1185 728
rect 1194 668 1198 671
rect 1142 663 1145 668
rect 1206 662 1209 678
rect 1230 662 1233 718
rect 1238 662 1241 728
rect 1218 658 1222 661
rect 1174 592 1177 638
rect 1058 588 1062 591
rect 1238 582 1241 658
rect 1046 562 1049 568
rect 1230 552 1233 558
rect 1090 548 1094 551
rect 1022 522 1025 548
rect 1030 542 1033 548
rect 1150 542 1153 548
rect 1050 528 1054 531
rect 1110 472 1113 538
rect 1118 522 1121 528
rect 1038 462 1041 468
rect 1126 462 1129 468
rect 1134 462 1137 538
rect 1154 528 1158 531
rect 1230 522 1233 538
rect 1150 482 1153 488
rect 1210 478 1214 481
rect 1058 458 1062 461
rect 1186 459 1190 462
rect 1102 452 1105 458
rect 998 352 1001 448
rect 1006 352 1009 358
rect 1014 342 1017 428
rect 848 303 850 307
rect 854 303 857 307
rect 861 303 864 307
rect 822 272 825 298
rect 886 292 889 318
rect 882 278 886 281
rect 806 262 809 268
rect 862 262 865 268
rect 818 258 822 261
rect 718 192 721 218
rect 658 78 662 81
rect 670 62 673 128
rect 694 72 697 168
rect 718 152 721 168
rect 726 158 734 161
rect 702 92 705 118
rect 710 102 713 138
rect 726 122 729 158
rect 738 138 742 141
rect 686 62 689 68
rect 246 52 249 59
rect 370 58 374 61
rect 634 58 638 61
rect 674 58 678 61
rect 646 52 649 58
rect 626 48 630 51
rect 710 42 713 78
rect 718 72 721 88
rect 798 82 801 118
rect 830 92 833 118
rect 838 82 841 168
rect 854 151 857 218
rect 848 103 850 107
rect 854 103 857 107
rect 861 103 864 107
rect 798 72 801 78
rect 846 72 849 78
rect 878 72 881 268
rect 894 242 897 338
rect 926 312 929 338
rect 886 152 889 158
rect 902 152 905 238
rect 918 192 921 278
rect 926 262 929 308
rect 942 252 945 338
rect 950 322 953 328
rect 982 302 985 318
rect 950 263 953 298
rect 990 291 993 318
rect 986 288 993 291
rect 1014 162 1017 338
rect 1046 282 1049 288
rect 1038 262 1041 268
rect 958 132 961 148
rect 1014 142 1017 158
rect 950 122 953 128
rect 926 72 929 78
rect 950 72 953 118
rect 1006 92 1009 98
rect 898 68 902 71
rect 814 62 817 68
rect 782 52 785 59
rect 822 42 825 68
rect 878 62 881 68
rect 910 62 913 68
rect 966 62 969 78
rect 1014 62 1017 108
rect 1022 72 1025 238
rect 1046 152 1049 258
rect 1062 152 1065 428
rect 1206 352 1209 358
rect 1194 348 1198 351
rect 1118 342 1121 348
rect 1202 338 1206 341
rect 1070 302 1073 318
rect 1070 292 1073 298
rect 1078 262 1081 338
rect 1094 312 1097 338
rect 1126 282 1129 318
rect 1214 301 1217 458
rect 1230 442 1233 518
rect 1238 352 1241 558
rect 1254 402 1257 728
rect 1270 702 1273 748
rect 1270 663 1273 668
rect 1278 592 1281 748
rect 1342 742 1345 748
rect 1306 728 1310 731
rect 1286 712 1289 718
rect 1286 672 1289 688
rect 1302 562 1305 718
rect 1282 548 1286 551
rect 1270 542 1273 548
rect 1294 522 1297 558
rect 1306 548 1310 551
rect 1302 532 1305 538
rect 1262 492 1265 518
rect 1326 512 1329 558
rect 1334 552 1337 728
rect 1350 692 1353 718
rect 1366 652 1369 748
rect 1398 712 1401 748
rect 1374 662 1377 668
rect 1382 652 1385 658
rect 1352 603 1354 607
rect 1358 603 1361 607
rect 1365 603 1368 607
rect 1346 558 1350 561
rect 1366 552 1369 568
rect 1390 552 1393 678
rect 1398 582 1401 618
rect 1398 562 1401 568
rect 1378 548 1382 551
rect 1294 492 1297 508
rect 1334 502 1337 538
rect 1270 472 1273 478
rect 1302 472 1305 498
rect 1302 462 1305 468
rect 1334 462 1337 468
rect 1314 458 1318 461
rect 1254 352 1257 398
rect 1270 362 1273 458
rect 1294 442 1297 448
rect 1226 348 1230 351
rect 1210 298 1217 301
rect 1206 282 1209 298
rect 1098 268 1102 271
rect 1086 242 1089 268
rect 1174 262 1177 268
rect 1214 262 1217 288
rect 1238 272 1241 348
rect 1246 332 1249 338
rect 1270 292 1273 358
rect 1302 342 1305 388
rect 1318 352 1321 418
rect 1342 402 1345 508
rect 1358 482 1361 488
rect 1374 432 1377 538
rect 1414 472 1417 748
rect 1430 712 1433 938
rect 1430 592 1433 678
rect 1430 551 1433 578
rect 1430 472 1433 528
rect 1406 452 1409 459
rect 1352 403 1354 407
rect 1358 403 1361 407
rect 1365 403 1368 407
rect 1334 362 1337 368
rect 1342 352 1345 398
rect 1378 368 1382 371
rect 1350 362 1353 368
rect 1330 348 1334 351
rect 1414 351 1417 358
rect 1310 342 1313 348
rect 1422 342 1425 468
rect 1438 382 1441 1158
rect 1446 1002 1449 1278
rect 1478 1262 1481 1268
rect 1558 1262 1561 1268
rect 1598 1262 1601 1298
rect 1638 1262 1641 1278
rect 1654 1262 1657 1268
rect 1522 1258 1526 1261
rect 1642 1258 1649 1261
rect 1666 1258 1670 1261
rect 1462 1192 1465 1258
rect 1470 1252 1473 1258
rect 1490 1228 1494 1231
rect 1454 1162 1457 1168
rect 1454 1092 1457 1148
rect 1462 1142 1465 1188
rect 1486 1152 1489 1208
rect 1502 1192 1505 1258
rect 1494 1152 1497 1158
rect 1470 1132 1473 1148
rect 1502 1141 1505 1148
rect 1490 1138 1505 1141
rect 1470 1092 1473 1128
rect 1518 1102 1521 1258
rect 1530 1148 1534 1151
rect 1482 1088 1486 1091
rect 1454 1072 1457 1078
rect 1502 1062 1505 1068
rect 1526 1062 1529 1068
rect 1534 1012 1537 1128
rect 1494 962 1497 968
rect 1450 958 1454 961
rect 1450 948 1454 951
rect 1478 942 1481 948
rect 1502 942 1505 968
rect 1454 872 1457 898
rect 1454 862 1457 868
rect 1462 862 1465 868
rect 1454 742 1457 748
rect 1462 692 1465 838
rect 1470 722 1473 868
rect 1478 862 1481 908
rect 1486 872 1489 928
rect 1494 852 1497 918
rect 1542 912 1545 1258
rect 1566 1248 1574 1251
rect 1550 1142 1553 1198
rect 1558 1152 1561 1188
rect 1550 1072 1553 1118
rect 1566 1082 1569 1248
rect 1606 1242 1609 1258
rect 1614 1252 1617 1258
rect 1602 1188 1606 1191
rect 1586 1148 1590 1151
rect 1558 952 1561 958
rect 1566 942 1569 1038
rect 1598 952 1601 1178
rect 1630 1152 1633 1218
rect 1610 1148 1614 1151
rect 1630 1122 1633 1138
rect 1610 1068 1614 1071
rect 1630 1062 1633 1068
rect 1646 1062 1649 1258
rect 1678 1252 1681 1298
rect 1702 1262 1705 1328
rect 1718 1292 1721 1298
rect 1710 1272 1713 1278
rect 1726 1271 1729 1458
rect 1734 1452 1737 1458
rect 1758 1452 1761 1468
rect 1766 1461 1769 1508
rect 1790 1472 1793 1478
rect 1798 1472 1801 1488
rect 1778 1468 1782 1471
rect 1766 1458 1774 1461
rect 1734 1282 1737 1448
rect 1782 1442 1785 1458
rect 1814 1392 1817 1608
rect 1822 1462 1825 1468
rect 1778 1388 1782 1391
rect 1822 1361 1825 1388
rect 1814 1358 1825 1361
rect 1798 1352 1801 1358
rect 1786 1348 1790 1351
rect 1726 1268 1737 1271
rect 1690 1258 1694 1261
rect 1726 1242 1729 1248
rect 1726 1192 1729 1238
rect 1734 1192 1737 1268
rect 1758 1192 1761 1308
rect 1770 1258 1774 1261
rect 1694 1172 1697 1178
rect 1654 1152 1657 1158
rect 1770 1148 1774 1151
rect 1654 1092 1657 1128
rect 1678 1062 1681 1148
rect 1610 1058 1614 1061
rect 1614 992 1617 998
rect 1502 862 1505 908
rect 1542 872 1545 888
rect 1566 862 1569 868
rect 1486 672 1489 738
rect 1518 722 1521 818
rect 1590 792 1593 828
rect 1606 822 1609 838
rect 1614 811 1617 918
rect 1622 862 1625 888
rect 1630 862 1633 1058
rect 1654 992 1657 1008
rect 1686 992 1689 1078
rect 1734 1072 1737 1118
rect 1742 1102 1745 1128
rect 1782 1122 1785 1268
rect 1814 1262 1817 1358
rect 1822 1322 1825 1348
rect 1830 1292 1833 1718
rect 1838 1542 1841 1548
rect 1846 1542 1849 1638
rect 1838 1392 1841 1408
rect 1838 1302 1841 1318
rect 1846 1282 1849 1528
rect 1854 1482 1857 1588
rect 1862 1532 1865 1878
rect 2006 1862 2009 1928
rect 2022 1892 2025 1948
rect 2038 1892 2041 1898
rect 2046 1892 2049 1948
rect 2058 1938 2062 1941
rect 2086 1932 2089 1938
rect 2054 1888 2062 1891
rect 2014 1872 2017 1878
rect 2030 1872 2033 1878
rect 2054 1872 2057 1888
rect 2070 1862 2073 1868
rect 1962 1858 1966 1861
rect 1942 1852 1945 1858
rect 2034 1848 2038 1851
rect 1918 1752 1921 1758
rect 1934 1752 1937 1798
rect 1990 1792 1993 1848
rect 2002 1818 2006 1821
rect 2022 1792 2025 1848
rect 1974 1752 1977 1768
rect 2010 1758 2014 1761
rect 1906 1748 1910 1751
rect 1978 1748 1982 1751
rect 1934 1732 1937 1748
rect 1966 1742 1969 1748
rect 1978 1738 1982 1741
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1885 1703 1888 1707
rect 1922 1688 1926 1691
rect 1934 1662 1937 1688
rect 1942 1682 1945 1738
rect 1950 1722 1953 1728
rect 1958 1722 1961 1728
rect 1958 1692 1961 1698
rect 1966 1682 1969 1718
rect 1906 1658 1910 1661
rect 1934 1652 1937 1658
rect 1890 1648 1894 1651
rect 1894 1592 1897 1598
rect 1898 1588 1902 1591
rect 1942 1582 1945 1658
rect 1950 1612 1953 1658
rect 1918 1562 1921 1568
rect 1958 1562 1961 1628
rect 1966 1562 1969 1678
rect 1974 1672 1977 1688
rect 1966 1552 1969 1558
rect 1974 1542 1977 1658
rect 1990 1642 1993 1748
rect 2014 1732 2017 1738
rect 2022 1721 2025 1748
rect 2014 1718 2025 1721
rect 2014 1692 2017 1718
rect 2002 1648 2006 1651
rect 2006 1592 2009 1608
rect 2022 1592 2025 1668
rect 2030 1662 2033 1808
rect 2038 1732 2041 1758
rect 2046 1752 2049 1798
rect 2070 1772 2073 1818
rect 2054 1762 2057 1768
rect 2038 1682 2041 1708
rect 2046 1702 2049 1738
rect 2062 1732 2065 1758
rect 2046 1682 2049 1688
rect 2038 1672 2041 1678
rect 2062 1662 2065 1728
rect 2078 1692 2081 1758
rect 2086 1751 2089 1908
rect 2094 1802 2097 2158
rect 2102 2152 2105 2168
rect 2146 2148 2150 2151
rect 2150 2072 2153 2078
rect 2166 2072 2169 2268
rect 2190 2192 2193 2308
rect 2214 2262 2217 2408
rect 2222 2372 2225 2418
rect 2222 2352 2225 2358
rect 2222 2272 2225 2348
rect 2230 2332 2233 2508
rect 2254 2482 2257 2488
rect 2278 2462 2281 2518
rect 2286 2512 2289 2548
rect 2302 2542 2305 2658
rect 2314 2648 2318 2651
rect 2326 2642 2329 2688
rect 2342 2682 2345 2738
rect 2358 2702 2361 3138
rect 2390 3072 2393 3138
rect 2414 3062 2417 3238
rect 2446 3212 2449 3258
rect 2490 3248 2494 3251
rect 2426 3148 2430 3151
rect 2426 3068 2430 3071
rect 2454 3062 2457 3078
rect 2374 3052 2377 3059
rect 2406 3058 2414 3061
rect 2366 2992 2369 3048
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2397 3003 2400 3007
rect 2406 2952 2409 3058
rect 2438 3052 2441 3058
rect 2446 2952 2449 3048
rect 2454 2952 2457 2988
rect 2426 2948 2430 2951
rect 2446 2942 2449 2948
rect 2390 2922 2393 2928
rect 2390 2891 2393 2918
rect 2386 2888 2393 2891
rect 2366 2862 2369 2868
rect 2366 2852 2369 2858
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2397 2803 2400 2807
rect 2386 2768 2390 2771
rect 2406 2752 2409 2798
rect 2422 2672 2425 2858
rect 2422 2652 2425 2658
rect 2302 2492 2305 2498
rect 2238 2442 2241 2458
rect 2238 2362 2241 2438
rect 2246 2392 2249 2448
rect 2270 2442 2273 2458
rect 2286 2452 2289 2458
rect 2310 2392 2313 2618
rect 2334 2552 2337 2598
rect 2342 2492 2345 2628
rect 2358 2542 2361 2638
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2397 2603 2400 2607
rect 2430 2562 2433 2868
rect 2438 2862 2441 2918
rect 2454 2901 2457 2948
rect 2446 2898 2457 2901
rect 2446 2752 2449 2898
rect 2462 2822 2465 3248
rect 2470 3192 2473 3198
rect 2482 3158 2494 3161
rect 2490 3148 2494 3151
rect 2478 3142 2481 3148
rect 2502 3142 2505 3258
rect 2526 3212 2529 3248
rect 2510 3182 2513 3198
rect 2510 3162 2513 3178
rect 2518 3152 2521 3158
rect 2506 3138 2510 3141
rect 2486 3092 2489 3128
rect 2526 3092 2529 3208
rect 2534 3152 2537 3228
rect 2550 3162 2553 3338
rect 2558 3332 2561 3348
rect 2566 3272 2569 3298
rect 2582 3292 2585 3348
rect 2598 3322 2601 3518
rect 2622 3432 2625 3548
rect 2634 3478 2638 3481
rect 2638 3462 2641 3468
rect 2622 3382 2625 3428
rect 2618 3348 2622 3351
rect 2614 3312 2617 3318
rect 2622 3211 2625 3348
rect 2630 3342 2633 3358
rect 2634 3338 2638 3341
rect 2638 3322 2641 3328
rect 2638 3272 2641 3298
rect 2646 3282 2649 3488
rect 2662 3441 2665 3548
rect 2674 3538 2678 3541
rect 2686 3472 2689 3478
rect 2678 3462 2681 3468
rect 2698 3458 2702 3461
rect 2670 3442 2673 3458
rect 2710 3452 2713 3628
rect 2726 3612 2729 3678
rect 2734 3672 2737 3748
rect 2798 3742 2801 3748
rect 2742 3702 2745 3738
rect 2782 3732 2785 3738
rect 2790 3732 2793 3738
rect 2814 3722 2817 3758
rect 2838 3752 2841 3858
rect 2826 3748 2830 3751
rect 2838 3742 2841 3748
rect 2846 3742 2849 3858
rect 2854 3852 2857 3918
rect 2870 3862 2873 3918
rect 2888 3903 2890 3907
rect 2894 3903 2897 3907
rect 2901 3903 2904 3907
rect 2918 3882 2921 3938
rect 3054 3932 3057 3938
rect 3110 3932 3113 3938
rect 2926 3892 2929 3908
rect 2974 3892 2977 3898
rect 2878 3872 2881 3878
rect 2974 3872 2977 3888
rect 2906 3868 2910 3871
rect 2914 3858 2918 3861
rect 2970 3858 2974 3861
rect 2862 3852 2865 3858
rect 2902 3841 2905 3858
rect 2926 3842 2929 3848
rect 2902 3838 2913 3841
rect 2846 3702 2849 3738
rect 2866 3718 2870 3721
rect 2802 3688 2806 3691
rect 2834 3678 2838 3681
rect 2790 3672 2793 3678
rect 2742 3592 2745 3658
rect 2766 3652 2769 3658
rect 2774 3652 2777 3658
rect 2750 3642 2753 3648
rect 2782 3632 2785 3668
rect 2814 3662 2817 3678
rect 2878 3671 2881 3728
rect 2888 3703 2890 3707
rect 2894 3703 2897 3707
rect 2901 3703 2904 3707
rect 2874 3668 2881 3671
rect 2842 3658 2846 3661
rect 2766 3612 2769 3618
rect 2746 3548 2750 3551
rect 2790 3542 2793 3578
rect 2798 3552 2801 3648
rect 2814 3612 2817 3658
rect 2854 3652 2857 3658
rect 2842 3648 2846 3651
rect 2870 3602 2873 3658
rect 2878 3652 2881 3658
rect 2898 3648 2902 3651
rect 2830 3572 2833 3578
rect 2814 3562 2817 3568
rect 2846 3562 2849 3568
rect 2862 3562 2865 3598
rect 2878 3582 2881 3618
rect 2830 3552 2833 3558
rect 2818 3548 2822 3551
rect 2774 3532 2777 3538
rect 2790 3502 2793 3538
rect 2662 3438 2670 3441
rect 2662 3352 2665 3438
rect 2726 3422 2729 3468
rect 2750 3462 2753 3488
rect 2798 3472 2801 3548
rect 2818 3538 2822 3541
rect 2830 3512 2833 3548
rect 2898 3547 2902 3550
rect 2854 3532 2857 3538
rect 2838 3482 2841 3488
rect 2814 3472 2817 3478
rect 2862 3462 2865 3508
rect 2870 3472 2873 3518
rect 2878 3472 2881 3538
rect 2910 3512 2913 3838
rect 2982 3792 2985 3928
rect 3126 3912 3129 3928
rect 3114 3878 3118 3881
rect 3046 3862 3049 3868
rect 3094 3862 3097 3878
rect 3118 3868 3126 3871
rect 3118 3862 3121 3868
rect 3134 3862 3137 3938
rect 3150 3862 3153 3868
rect 3074 3858 3078 3861
rect 3130 3858 3134 3861
rect 3038 3832 3041 3838
rect 3086 3812 3089 3858
rect 2982 3752 2985 3788
rect 3050 3768 3054 3771
rect 3030 3762 3033 3768
rect 3022 3752 3025 3758
rect 2922 3748 2926 3751
rect 2950 3742 2953 3748
rect 2966 3712 2969 3728
rect 2974 3722 2977 3728
rect 2974 3701 2977 3708
rect 2966 3698 2977 3701
rect 2982 3702 2985 3738
rect 2998 3732 3001 3748
rect 2918 3672 2921 3698
rect 2966 3692 2969 3698
rect 2974 3682 2977 3688
rect 2986 3678 2990 3681
rect 2970 3668 2974 3671
rect 2918 3632 2921 3668
rect 2958 3662 2961 3668
rect 2982 3662 2985 3668
rect 3006 3662 3009 3748
rect 3046 3742 3049 3758
rect 3086 3752 3089 3788
rect 2930 3658 2934 3661
rect 2946 3658 2950 3661
rect 3014 3652 3017 3668
rect 2946 3648 2950 3651
rect 2926 3642 2929 3648
rect 2974 3592 2977 3648
rect 3022 3592 3025 3678
rect 3030 3672 3033 3718
rect 3102 3692 3105 3818
rect 3110 3712 3113 3748
rect 3090 3688 3094 3691
rect 3038 3672 3041 3688
rect 3118 3672 3121 3858
rect 3158 3792 3161 3938
rect 3198 3922 3201 3948
rect 3214 3922 3217 3928
rect 3182 3852 3185 3918
rect 3214 3882 3217 3918
rect 3226 3858 3230 3861
rect 3150 3742 3153 3758
rect 3158 3732 3161 3748
rect 3166 3672 3169 3818
rect 3174 3752 3177 3758
rect 3182 3752 3185 3828
rect 3206 3742 3209 3788
rect 3230 3752 3233 3758
rect 3238 3752 3241 4058
rect 3246 4052 3249 4138
rect 3278 4132 3281 4138
rect 3270 4082 3273 4088
rect 3278 4082 3281 4088
rect 3286 4072 3289 4198
rect 3262 4062 3265 4068
rect 3294 4062 3297 4218
rect 3302 4162 3305 4198
rect 3310 4102 3313 4138
rect 3302 4072 3305 4078
rect 3254 4052 3257 4058
rect 3246 4042 3249 4048
rect 3310 4042 3313 4048
rect 3286 3951 3289 3968
rect 3302 3942 3305 3998
rect 3318 3952 3321 4178
rect 3374 4152 3377 4338
rect 3390 4322 3393 4338
rect 3422 4332 3425 4468
rect 3430 4352 3433 4778
rect 3446 4752 3449 4968
rect 3462 4952 3465 4978
rect 3470 4901 3473 5008
rect 3550 5002 3553 5058
rect 3558 4982 3561 5058
rect 3630 4992 3633 5058
rect 3654 5012 3657 5058
rect 3542 4972 3545 4978
rect 3530 4968 3534 4971
rect 3558 4962 3561 4968
rect 3490 4947 3494 4950
rect 3462 4898 3473 4901
rect 3462 4862 3465 4898
rect 3502 4872 3505 4878
rect 3510 4862 3513 4958
rect 3542 4952 3545 4958
rect 3630 4952 3633 4978
rect 3662 4962 3665 4968
rect 3650 4958 3654 4961
rect 3554 4948 3558 4951
rect 3658 4948 3662 4951
rect 3574 4942 3577 4948
rect 3590 4942 3593 4948
rect 3614 4942 3617 4948
rect 3658 4938 3665 4941
rect 3550 4882 3553 4938
rect 3582 4922 3585 4938
rect 3566 4872 3569 4918
rect 3614 4892 3617 4938
rect 3622 4922 3625 4938
rect 3626 4918 3633 4921
rect 3594 4888 3598 4891
rect 3550 4862 3553 4868
rect 3498 4838 3502 4841
rect 3478 4792 3481 4838
rect 3526 4802 3529 4838
rect 3542 4752 3545 4858
rect 3446 4742 3449 4748
rect 3494 4742 3497 4748
rect 3462 4672 3465 4678
rect 3438 4662 3441 4668
rect 3470 4662 3473 4738
rect 3486 4652 3489 4698
rect 3502 4662 3505 4708
rect 3518 4692 3521 4748
rect 3494 4652 3497 4658
rect 3458 4648 3462 4651
rect 3438 4481 3441 4618
rect 3450 4548 3454 4551
rect 3446 4532 3449 4538
rect 3462 4532 3465 4548
rect 3470 4542 3473 4618
rect 3494 4582 3497 4648
rect 3478 4552 3481 4558
rect 3494 4522 3497 4578
rect 3502 4542 3505 4618
rect 3542 4571 3545 4738
rect 3566 4732 3569 4868
rect 3614 4862 3617 4888
rect 3622 4872 3625 4878
rect 3630 4872 3633 4918
rect 3654 4892 3657 4918
rect 3662 4872 3665 4938
rect 3670 4882 3673 5058
rect 3702 5042 3705 5058
rect 3710 5052 3713 5058
rect 3726 5052 3729 5058
rect 3678 4942 3681 4958
rect 3686 4942 3689 5018
rect 3694 4952 3697 5038
rect 3702 4992 3705 4998
rect 3718 4952 3721 5038
rect 3734 5022 3737 5058
rect 3694 4872 3697 4938
rect 3718 4931 3721 4948
rect 3726 4942 3729 4948
rect 3718 4928 3729 4931
rect 3574 4852 3577 4858
rect 3594 4848 3598 4851
rect 3614 4842 3617 4848
rect 3602 4838 3606 4841
rect 3582 4792 3585 4798
rect 3606 4791 3609 4838
rect 3622 4812 3625 4868
rect 3606 4788 3617 4791
rect 3574 4712 3577 4718
rect 3550 4682 3553 4708
rect 3566 4662 3569 4678
rect 3590 4652 3593 4678
rect 3598 4671 3601 4728
rect 3614 4672 3617 4788
rect 3598 4668 3606 4671
rect 3630 4662 3633 4858
rect 3654 4842 3657 4848
rect 3662 4812 3665 4868
rect 3674 4858 3678 4861
rect 3702 4861 3705 4928
rect 3694 4858 3705 4861
rect 3670 4842 3673 4848
rect 3638 4752 3641 4758
rect 3662 4742 3665 4748
rect 3678 4742 3681 4808
rect 3686 4752 3689 4858
rect 3694 4852 3697 4858
rect 3714 4848 3718 4851
rect 3702 4762 3705 4768
rect 3726 4752 3729 4928
rect 3758 4922 3761 4947
rect 3766 4942 3769 5008
rect 3798 4992 3801 5058
rect 3838 5052 3841 5058
rect 3838 5002 3841 5048
rect 3846 4972 3849 4988
rect 3790 4952 3793 4958
rect 3734 4862 3737 4878
rect 3742 4852 3745 4868
rect 3750 4832 3753 4868
rect 3758 4862 3761 4888
rect 3734 4792 3737 4818
rect 3662 4701 3665 4738
rect 3678 4712 3681 4738
rect 3662 4698 3673 4701
rect 3638 4682 3641 4688
rect 3670 4682 3673 4698
rect 3678 4662 3681 4668
rect 3542 4568 3553 4571
rect 3510 4542 3513 4558
rect 3530 4548 3534 4551
rect 3550 4542 3553 4568
rect 3530 4538 3534 4541
rect 3438 4478 3449 4481
rect 3438 4362 3441 4468
rect 3446 4382 3449 4478
rect 3430 4331 3433 4348
rect 3438 4342 3441 4358
rect 3446 4342 3449 4348
rect 3430 4328 3441 4331
rect 3390 4262 3393 4268
rect 3438 4262 3441 4328
rect 3454 4261 3457 4518
rect 3450 4258 3457 4261
rect 3462 4262 3465 4448
rect 3334 4142 3337 4148
rect 3358 4132 3361 4138
rect 3326 4092 3329 4128
rect 3350 4072 3353 4078
rect 3326 3972 3329 3978
rect 3318 3942 3321 3948
rect 3262 3902 3265 3938
rect 3262 3872 3265 3898
rect 3286 3892 3289 3928
rect 3318 3902 3321 3918
rect 3318 3892 3321 3898
rect 3278 3872 3281 3878
rect 3306 3858 3310 3861
rect 3294 3842 3297 3848
rect 3266 3778 3270 3781
rect 3218 3748 3222 3751
rect 3182 3732 3185 3738
rect 3266 3728 3270 3731
rect 3198 3722 3201 3728
rect 3254 3702 3257 3718
rect 3242 3668 3246 3671
rect 3046 3662 3049 3668
rect 3086 3662 3089 3668
rect 3034 3658 3038 3661
rect 3162 3658 3166 3661
rect 3054 3642 3057 3658
rect 3058 3588 3062 3591
rect 2962 3568 2966 3571
rect 2994 3558 2998 3561
rect 2974 3552 2977 3558
rect 3030 3552 3033 3568
rect 3054 3562 3057 3568
rect 3050 3548 3054 3551
rect 2888 3503 2890 3507
rect 2894 3503 2897 3507
rect 2901 3503 2904 3507
rect 2822 3452 2825 3458
rect 2750 3442 2753 3448
rect 2846 3442 2849 3448
rect 2810 3438 2814 3441
rect 2678 3362 2681 3398
rect 2694 3382 2697 3418
rect 2674 3358 2678 3361
rect 2694 3352 2697 3368
rect 2710 3352 2713 3408
rect 2738 3358 2742 3361
rect 2750 3352 2753 3438
rect 2722 3348 2726 3351
rect 2762 3348 2766 3351
rect 2654 3342 2657 3348
rect 2702 3342 2705 3348
rect 2782 3342 2785 3418
rect 2798 3351 2801 3358
rect 2654 3292 2657 3338
rect 2670 3321 2673 3328
rect 2662 3318 2673 3321
rect 2662 3312 2665 3318
rect 2662 3272 2665 3308
rect 2670 3262 2673 3288
rect 2678 3272 2681 3288
rect 2686 3281 2689 3338
rect 2766 3332 2769 3338
rect 2710 3292 2713 3318
rect 2686 3278 2694 3281
rect 2726 3272 2729 3278
rect 2742 3272 2745 3298
rect 2690 3268 2694 3271
rect 2622 3208 2633 3211
rect 2606 3192 2609 3198
rect 2546 3158 2550 3161
rect 2574 3152 2577 3178
rect 2618 3158 2622 3161
rect 2566 3142 2569 3148
rect 2630 3142 2633 3208
rect 2638 3152 2641 3168
rect 2646 3151 2649 3228
rect 2654 3162 2657 3168
rect 2646 3148 2654 3151
rect 2662 3142 2665 3258
rect 2670 3222 2673 3258
rect 2670 3162 2673 3168
rect 2534 3132 2537 3138
rect 2546 3118 2550 3121
rect 2478 3082 2481 3088
rect 2494 3072 2497 3088
rect 2558 3082 2561 3138
rect 2598 3102 2601 3138
rect 2566 3092 2569 3098
rect 2630 3092 2633 3138
rect 2654 3132 2657 3138
rect 2662 3122 2665 3138
rect 2678 3082 2681 3268
rect 2790 3262 2793 3308
rect 2806 3272 2809 3378
rect 2862 3342 2865 3368
rect 2886 3352 2889 3438
rect 2902 3352 2905 3448
rect 2926 3412 2929 3548
rect 2962 3538 2966 3541
rect 2998 3522 3001 3548
rect 3006 3492 3009 3538
rect 3022 3532 3025 3548
rect 3122 3547 3126 3550
rect 3142 3542 3145 3658
rect 3190 3642 3193 3668
rect 3206 3652 3209 3668
rect 3270 3662 3273 3668
rect 3234 3658 3238 3661
rect 3214 3652 3217 3658
rect 3214 3611 3217 3618
rect 3214 3608 3222 3611
rect 3246 3592 3249 3598
rect 3158 3562 3161 3588
rect 3174 3572 3177 3578
rect 3190 3562 3193 3568
rect 3186 3548 3190 3551
rect 3242 3548 3246 3551
rect 3034 3538 3038 3541
rect 2950 3472 2953 3488
rect 2978 3478 2982 3481
rect 3006 3472 3009 3488
rect 2966 3462 2969 3468
rect 2990 3462 2993 3468
rect 3078 3462 3081 3478
rect 3102 3472 3105 3538
rect 3174 3531 3177 3548
rect 3186 3538 3190 3541
rect 3174 3528 3185 3531
rect 3158 3492 3161 3518
rect 3182 3492 3185 3528
rect 3206 3522 3209 3548
rect 3214 3502 3217 3538
rect 3254 3532 3257 3618
rect 3222 3522 3225 3528
rect 3206 3472 3209 3488
rect 3170 3468 3174 3471
rect 3002 3458 3006 3461
rect 2950 3452 2953 3458
rect 2950 3422 2953 3448
rect 2942 3351 2945 3418
rect 2898 3338 2902 3341
rect 2966 3322 2969 3458
rect 2974 3352 2977 3408
rect 2870 3302 2873 3318
rect 2888 3303 2890 3307
rect 2894 3303 2897 3307
rect 2901 3303 2904 3307
rect 2814 3262 2817 3298
rect 2838 3272 2841 3288
rect 2870 3272 2873 3288
rect 2926 3262 2929 3298
rect 2946 3288 2950 3291
rect 2958 3262 2961 3288
rect 2966 3272 2969 3298
rect 2990 3282 2993 3328
rect 2990 3272 2993 3278
rect 2834 3258 2846 3261
rect 2890 3258 2894 3261
rect 2702 3252 2705 3258
rect 2718 3242 2721 3248
rect 2750 3232 2753 3258
rect 2758 3252 2761 3258
rect 2726 3182 2729 3218
rect 2766 3202 2769 3258
rect 2834 3248 2838 3251
rect 2782 3182 2785 3218
rect 2794 3168 2801 3171
rect 2686 3162 2689 3168
rect 2790 3162 2793 3168
rect 2798 3152 2801 3168
rect 2726 3132 2729 3148
rect 2790 3142 2793 3148
rect 2558 3072 2561 3078
rect 2594 3068 2598 3071
rect 2470 3062 2473 3068
rect 2558 3062 2561 3068
rect 2606 3062 2609 3068
rect 2630 3062 2633 3068
rect 2638 3062 2641 3068
rect 2514 3058 2518 3061
rect 2594 3058 2598 3061
rect 2610 3058 2614 3061
rect 2470 3022 2473 3058
rect 2470 2992 2473 2998
rect 2502 2972 2505 3058
rect 2582 3052 2585 3058
rect 2538 3048 2542 3051
rect 2626 3048 2630 3051
rect 2478 2892 2481 2968
rect 2506 2948 2510 2951
rect 2490 2938 2494 2941
rect 2526 2941 2529 3018
rect 2550 2982 2553 3018
rect 2566 3012 2569 3048
rect 2566 2952 2569 2988
rect 2682 2968 2686 2971
rect 2574 2952 2577 2958
rect 2646 2952 2649 2958
rect 2518 2938 2529 2941
rect 2618 2948 2622 2951
rect 2510 2922 2513 2938
rect 2442 2738 2446 2741
rect 2446 2642 2449 2668
rect 2462 2662 2465 2808
rect 2486 2802 2489 2918
rect 2510 2862 2513 2868
rect 2518 2852 2521 2938
rect 2526 2882 2529 2928
rect 2534 2912 2537 2948
rect 2562 2938 2566 2941
rect 2554 2928 2558 2931
rect 2582 2922 2585 2948
rect 2654 2942 2657 2948
rect 2598 2902 2601 2918
rect 2602 2888 2606 2891
rect 2574 2882 2577 2888
rect 2486 2752 2489 2768
rect 2502 2762 2505 2768
rect 2518 2762 2521 2848
rect 2526 2822 2529 2878
rect 2558 2872 2561 2878
rect 2614 2872 2617 2938
rect 2622 2892 2625 2928
rect 2630 2902 2633 2918
rect 2638 2912 2641 2938
rect 2670 2932 2673 2958
rect 2702 2952 2705 3088
rect 2718 3072 2721 3128
rect 2782 3092 2785 3118
rect 2790 3112 2793 3138
rect 2758 3072 2761 3078
rect 2718 3052 2721 3058
rect 2726 2972 2729 3068
rect 2778 3058 2782 3061
rect 2778 3048 2782 3051
rect 2806 3051 2809 3238
rect 2858 3218 2862 3221
rect 2818 3158 2822 3161
rect 2814 3062 2817 3118
rect 2830 3062 2833 3208
rect 2870 3192 2873 3258
rect 2902 3242 2905 3258
rect 2838 3162 2841 3168
rect 2846 3142 2849 3148
rect 2854 3142 2857 3158
rect 2838 3132 2841 3138
rect 2878 3102 2881 3158
rect 2894 3152 2897 3188
rect 2902 3132 2905 3138
rect 2888 3103 2890 3107
rect 2894 3103 2897 3107
rect 2901 3103 2904 3107
rect 2838 3062 2841 3068
rect 2846 3062 2849 3078
rect 2878 3062 2881 3088
rect 2858 3058 2862 3061
rect 2890 3058 2894 3061
rect 2830 3052 2833 3058
rect 2806 3048 2814 3051
rect 2778 3038 2782 3041
rect 2814 2972 2817 3048
rect 2866 3038 2870 3041
rect 2710 2962 2713 2968
rect 2766 2952 2769 2968
rect 2638 2872 2641 2878
rect 2542 2863 2545 2868
rect 2590 2862 2593 2868
rect 2614 2862 2617 2868
rect 2622 2862 2625 2868
rect 2658 2859 2662 2862
rect 2558 2762 2561 2768
rect 2494 2752 2497 2758
rect 2534 2752 2537 2758
rect 2546 2748 2550 2751
rect 2478 2722 2481 2748
rect 2510 2732 2513 2748
rect 2558 2741 2561 2758
rect 2606 2752 2609 2758
rect 2550 2738 2561 2741
rect 2634 2748 2638 2751
rect 2510 2722 2513 2728
rect 2462 2612 2465 2658
rect 2470 2652 2473 2718
rect 2478 2692 2481 2698
rect 2502 2642 2505 2668
rect 2518 2652 2521 2659
rect 2402 2558 2406 2561
rect 2446 2542 2449 2558
rect 2374 2462 2377 2478
rect 2382 2472 2385 2518
rect 2254 2352 2257 2368
rect 2262 2352 2265 2358
rect 2294 2352 2297 2358
rect 2242 2348 2246 2351
rect 2242 2338 2246 2341
rect 2230 2292 2233 2308
rect 2246 2262 2249 2268
rect 2254 2262 2257 2348
rect 2290 2338 2294 2341
rect 2270 2302 2273 2338
rect 2278 2282 2281 2338
rect 2286 2322 2289 2328
rect 2318 2322 2321 2458
rect 2326 2442 2329 2458
rect 2326 2352 2329 2438
rect 2342 2352 2345 2398
rect 2326 2291 2329 2348
rect 2334 2332 2337 2348
rect 2334 2302 2337 2328
rect 2326 2288 2334 2291
rect 2334 2272 2337 2288
rect 2282 2268 2286 2271
rect 2198 2162 2201 2218
rect 2214 2192 2217 2218
rect 2238 2152 2241 2198
rect 2246 2192 2249 2238
rect 2254 2162 2257 2258
rect 2262 2172 2265 2268
rect 2350 2262 2353 2458
rect 2358 2382 2361 2448
rect 2382 2442 2385 2468
rect 2406 2452 2409 2518
rect 2422 2462 2425 2498
rect 2430 2472 2433 2538
rect 2414 2452 2417 2458
rect 2374 2432 2377 2438
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2397 2403 2400 2407
rect 2430 2401 2433 2438
rect 2438 2412 2441 2518
rect 2478 2492 2481 2528
rect 2478 2472 2481 2488
rect 2458 2458 2462 2461
rect 2430 2398 2441 2401
rect 2358 2302 2361 2318
rect 2298 2258 2302 2261
rect 2278 2202 2281 2218
rect 2178 2148 2182 2151
rect 2294 2151 2297 2218
rect 2302 2212 2305 2258
rect 2310 2252 2313 2258
rect 2302 2162 2305 2168
rect 2286 2148 2297 2151
rect 2310 2151 2313 2188
rect 2318 2172 2321 2258
rect 2358 2202 2361 2268
rect 2318 2152 2321 2158
rect 2310 2148 2318 2151
rect 2102 2062 2105 2068
rect 2110 2052 2113 2068
rect 2102 1972 2105 2048
rect 2110 1992 2113 2028
rect 2118 1992 2121 2058
rect 2126 2052 2129 2058
rect 2134 2052 2137 2058
rect 2134 1992 2137 1998
rect 2126 1952 2129 1968
rect 2114 1948 2118 1951
rect 2114 1938 2118 1941
rect 2126 1932 2129 1938
rect 2142 1932 2145 2038
rect 2150 1962 2153 2058
rect 2166 2052 2169 2059
rect 2158 1872 2161 1918
rect 2166 1902 2169 1918
rect 2214 1892 2217 2098
rect 2230 2052 2233 2148
rect 2254 2142 2257 2148
rect 2278 2142 2281 2148
rect 2266 2138 2270 2141
rect 2286 2132 2289 2148
rect 2302 2142 2305 2148
rect 2254 2112 2257 2128
rect 2238 2082 2241 2088
rect 2246 2082 2249 2088
rect 2246 2068 2254 2071
rect 2230 1972 2233 2018
rect 2246 1972 2249 2068
rect 2270 2062 2273 2128
rect 2294 2122 2297 2138
rect 2310 2092 2313 2108
rect 2326 2072 2329 2148
rect 2350 2142 2353 2148
rect 2358 2072 2361 2148
rect 2366 2082 2369 2348
rect 2374 2342 2377 2388
rect 2418 2368 2422 2371
rect 2402 2348 2406 2351
rect 2374 2312 2377 2338
rect 2374 2272 2377 2308
rect 2374 2252 2377 2258
rect 2382 2242 2385 2258
rect 2410 2248 2414 2251
rect 2374 2192 2377 2208
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2397 2203 2400 2207
rect 2414 2192 2417 2228
rect 2414 2102 2417 2118
rect 2422 2092 2425 2358
rect 2430 2352 2433 2358
rect 2438 2352 2441 2398
rect 2446 2392 2449 2418
rect 2462 2392 2465 2448
rect 2438 2272 2441 2348
rect 2446 2272 2449 2348
rect 2430 2262 2433 2268
rect 2438 2152 2441 2168
rect 2446 2152 2449 2218
rect 2430 2112 2433 2148
rect 2438 2122 2441 2148
rect 2418 2078 2422 2081
rect 2298 2068 2302 2071
rect 2262 2022 2265 2058
rect 2226 1938 2230 1941
rect 2262 1922 2265 1938
rect 2174 1872 2177 1878
rect 2222 1872 2225 1898
rect 2230 1882 2233 1918
rect 2270 1892 2273 2058
rect 2294 2052 2297 2068
rect 2326 2062 2329 2068
rect 2358 2062 2361 2068
rect 2438 2062 2441 2108
rect 2386 2028 2390 2031
rect 2314 2018 2318 2021
rect 2342 1992 2345 2018
rect 2374 1992 2377 2008
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2397 2003 2400 2007
rect 2430 1992 2433 2058
rect 2286 1892 2289 1948
rect 2294 1942 2297 1958
rect 2362 1948 2366 1951
rect 2410 1948 2414 1951
rect 2334 1922 2337 1928
rect 2330 1888 2334 1891
rect 2270 1872 2273 1878
rect 2342 1872 2345 1888
rect 2086 1748 2094 1751
rect 2102 1742 2105 1778
rect 2118 1752 2121 1868
rect 2238 1862 2241 1868
rect 2186 1858 2190 1861
rect 2134 1792 2137 1858
rect 2162 1778 2166 1781
rect 2086 1692 2089 1738
rect 2102 1702 2105 1738
rect 2034 1658 2041 1661
rect 1930 1538 1934 1541
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1885 1503 1888 1507
rect 1926 1501 1929 1518
rect 1922 1498 1929 1501
rect 1854 1462 1857 1478
rect 1862 1472 1865 1498
rect 1934 1481 1937 1538
rect 1966 1532 1969 1538
rect 1958 1512 1961 1518
rect 1926 1478 1937 1481
rect 1942 1482 1945 1508
rect 1918 1462 1921 1468
rect 1890 1458 1894 1461
rect 1906 1458 1910 1461
rect 1838 1272 1841 1278
rect 1822 1262 1825 1268
rect 1842 1258 1846 1261
rect 1854 1192 1857 1438
rect 1862 1332 1865 1358
rect 1894 1351 1897 1398
rect 1878 1342 1881 1348
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1885 1303 1888 1307
rect 1862 1282 1865 1288
rect 1822 1162 1825 1168
rect 1842 1148 1846 1151
rect 1758 1112 1761 1118
rect 1758 1092 1761 1098
rect 1798 1092 1801 1118
rect 1822 1082 1825 1118
rect 1718 1062 1721 1068
rect 1750 1062 1753 1068
rect 1738 1058 1742 1061
rect 1810 1058 1814 1061
rect 1710 1042 1713 1058
rect 1670 952 1673 958
rect 1658 948 1662 951
rect 1638 922 1641 948
rect 1678 942 1681 948
rect 1686 902 1689 958
rect 1694 882 1697 1018
rect 1706 948 1710 951
rect 1742 942 1745 948
rect 1730 938 1734 941
rect 1646 862 1649 878
rect 1686 872 1689 878
rect 1654 862 1657 868
rect 1630 852 1633 858
rect 1670 852 1673 868
rect 1702 862 1705 928
rect 1718 922 1721 928
rect 1726 892 1729 908
rect 1714 868 1718 871
rect 1690 858 1694 861
rect 1730 858 1734 861
rect 1614 808 1622 811
rect 1614 752 1617 798
rect 1678 792 1681 858
rect 1742 852 1745 858
rect 1714 848 1718 851
rect 1750 842 1753 948
rect 1762 918 1766 921
rect 1758 862 1761 888
rect 1758 852 1761 858
rect 1694 772 1697 818
rect 1750 762 1753 838
rect 1766 812 1769 918
rect 1530 748 1534 751
rect 1658 748 1662 751
rect 1542 732 1545 738
rect 1502 692 1505 708
rect 1542 692 1545 728
rect 1542 682 1545 688
rect 1574 682 1577 748
rect 1606 732 1609 748
rect 1630 742 1633 748
rect 1710 722 1713 738
rect 1718 722 1721 738
rect 1610 688 1614 691
rect 1450 658 1454 661
rect 1490 658 1494 661
rect 1470 602 1473 648
rect 1510 642 1513 678
rect 1638 672 1641 708
rect 1670 672 1673 718
rect 1678 682 1681 688
rect 1686 682 1689 688
rect 1650 668 1654 671
rect 1562 658 1566 661
rect 1490 588 1494 591
rect 1510 552 1513 628
rect 1574 621 1577 658
rect 1614 652 1617 668
rect 1678 662 1681 678
rect 1718 662 1721 668
rect 1622 652 1625 658
rect 1574 618 1585 621
rect 1574 562 1577 608
rect 1502 532 1505 538
rect 1466 488 1470 491
rect 1486 472 1489 478
rect 1526 462 1529 518
rect 1534 482 1537 558
rect 1574 552 1577 558
rect 1550 542 1553 548
rect 1558 542 1561 548
rect 1566 532 1569 538
rect 1570 488 1574 491
rect 1582 472 1585 618
rect 1590 562 1593 568
rect 1598 552 1601 638
rect 1630 632 1633 658
rect 1646 652 1649 658
rect 1662 652 1665 658
rect 1726 652 1729 748
rect 1742 742 1745 758
rect 1766 752 1769 788
rect 1750 742 1753 748
rect 1758 682 1761 738
rect 1774 691 1777 978
rect 1806 942 1809 948
rect 1806 871 1809 918
rect 1822 872 1825 888
rect 1798 870 1809 871
rect 1798 868 1806 870
rect 1782 862 1785 868
rect 1782 752 1785 808
rect 1790 742 1793 778
rect 1782 732 1785 738
rect 1774 688 1785 691
rect 1774 672 1777 678
rect 1782 662 1785 688
rect 1790 682 1793 738
rect 1798 702 1801 868
rect 1818 868 1822 871
rect 1806 792 1809 848
rect 1822 752 1825 768
rect 1830 741 1833 858
rect 1838 792 1841 1098
rect 1854 1062 1857 1068
rect 1862 1062 1865 1278
rect 1926 1272 1929 1478
rect 1946 1468 1950 1471
rect 1934 1462 1937 1468
rect 1958 1412 1961 1468
rect 1966 1462 1969 1488
rect 1974 1462 1977 1468
rect 1982 1422 1985 1578
rect 1994 1558 1998 1561
rect 2026 1558 2030 1561
rect 2038 1552 2041 1658
rect 2030 1542 2033 1548
rect 2046 1542 2049 1548
rect 2002 1538 2006 1541
rect 2034 1528 2038 1531
rect 1998 1492 2001 1528
rect 2026 1468 2033 1471
rect 2014 1462 2017 1468
rect 1974 1392 1977 1408
rect 1958 1362 1961 1368
rect 1982 1351 1985 1418
rect 1978 1348 1985 1351
rect 1942 1272 1945 1278
rect 1938 1248 1942 1251
rect 1894 1202 1897 1218
rect 1950 1202 1953 1258
rect 1958 1242 1961 1348
rect 1966 1332 1969 1338
rect 1970 1288 1974 1291
rect 1982 1282 1985 1298
rect 1982 1272 1985 1278
rect 1990 1262 1993 1458
rect 2006 1441 2009 1458
rect 2022 1452 2025 1458
rect 2006 1438 2014 1441
rect 2030 1392 2033 1468
rect 2038 1451 2041 1528
rect 2046 1492 2049 1518
rect 2054 1472 2057 1498
rect 2062 1472 2065 1658
rect 2070 1652 2073 1668
rect 2086 1652 2089 1678
rect 2094 1652 2097 1688
rect 2110 1662 2113 1748
rect 2142 1742 2145 1748
rect 2158 1732 2161 1748
rect 2166 1682 2169 1768
rect 2174 1722 2177 1728
rect 2182 1692 2185 1858
rect 2202 1848 2206 1851
rect 2118 1662 2121 1668
rect 2126 1662 2129 1668
rect 2114 1638 2118 1641
rect 2110 1552 2113 1588
rect 2134 1552 2137 1618
rect 2166 1592 2169 1678
rect 2174 1592 2177 1658
rect 2190 1552 2193 1838
rect 2178 1548 2182 1551
rect 2078 1492 2081 1547
rect 2142 1522 2145 1528
rect 2138 1518 2142 1521
rect 2058 1458 2062 1461
rect 2086 1452 2089 1518
rect 2150 1512 2153 1548
rect 2122 1488 2126 1491
rect 2114 1468 2118 1471
rect 2038 1448 2046 1451
rect 2078 1442 2081 1448
rect 2102 1442 2105 1448
rect 2014 1362 2017 1368
rect 2046 1352 2049 1358
rect 2094 1352 2097 1368
rect 2034 1348 2038 1351
rect 2014 1342 2017 1348
rect 1998 1322 2001 1338
rect 2014 1292 2017 1308
rect 2014 1272 2017 1288
rect 2022 1262 2025 1338
rect 2010 1258 2014 1261
rect 1982 1192 1985 1208
rect 1874 1148 1878 1151
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1885 1103 1888 1107
rect 1894 1092 1897 1108
rect 1918 1092 1921 1147
rect 1934 1122 1937 1138
rect 1950 1082 1953 1128
rect 1990 1072 1993 1258
rect 2022 1252 2025 1258
rect 2006 1242 2009 1248
rect 2022 1232 2025 1238
rect 2030 1192 2033 1328
rect 2078 1272 2081 1328
rect 2110 1312 2113 1458
rect 2038 1252 2041 1258
rect 2070 1252 2073 1259
rect 2030 1182 2033 1188
rect 2070 1152 2073 1188
rect 2058 1148 2062 1151
rect 2014 1142 2017 1148
rect 1998 1072 2001 1118
rect 2006 1082 2009 1088
rect 2038 1082 2041 1118
rect 2046 1102 2049 1148
rect 1910 1062 1913 1068
rect 1958 1062 1961 1068
rect 1966 1062 1969 1068
rect 1938 1058 1942 1061
rect 1862 892 1865 1058
rect 1882 1048 1886 1051
rect 1902 982 1905 1058
rect 1982 1042 1985 1048
rect 1962 968 1966 971
rect 1966 952 1969 958
rect 1990 952 1993 1058
rect 2038 1052 2041 1059
rect 1998 972 2001 988
rect 2030 972 2033 1008
rect 2054 992 2057 1128
rect 2070 1012 2073 1128
rect 2078 1122 2081 1268
rect 2102 1252 2105 1258
rect 2090 1168 2094 1171
rect 2094 1152 2097 1158
rect 2102 1142 2105 1218
rect 2126 1192 2129 1448
rect 2142 1362 2145 1368
rect 2150 1352 2153 1458
rect 2158 1422 2161 1548
rect 2182 1482 2185 1518
rect 2174 1462 2177 1478
rect 2198 1382 2201 1848
rect 2230 1822 2233 1858
rect 2222 1792 2225 1798
rect 2206 1752 2209 1768
rect 2214 1732 2217 1738
rect 2214 1632 2217 1728
rect 2230 1672 2233 1688
rect 2254 1662 2257 1748
rect 2262 1712 2265 1868
rect 2270 1792 2273 1828
rect 2318 1822 2321 1868
rect 2334 1862 2337 1868
rect 2246 1602 2249 1618
rect 2230 1562 2233 1588
rect 2214 1472 2217 1518
rect 2222 1472 2225 1478
rect 2230 1462 2233 1558
rect 2254 1552 2257 1658
rect 2262 1642 2265 1708
rect 2286 1692 2289 1808
rect 2310 1752 2313 1818
rect 2326 1792 2329 1828
rect 2294 1662 2297 1718
rect 2342 1662 2345 1748
rect 2358 1732 2361 1928
rect 2422 1912 2425 1918
rect 2406 1862 2409 1888
rect 2414 1872 2417 1898
rect 2430 1892 2433 1988
rect 2438 1952 2441 2058
rect 2446 1962 2449 2078
rect 2454 2062 2457 2328
rect 2462 2262 2465 2268
rect 2470 2262 2473 2468
rect 2486 2392 2489 2608
rect 2502 2552 2505 2638
rect 2494 2542 2497 2548
rect 2502 2352 2505 2358
rect 2510 2352 2513 2508
rect 2518 2332 2521 2338
rect 2486 2292 2489 2328
rect 2494 2282 2497 2308
rect 2526 2301 2529 2738
rect 2542 2722 2545 2738
rect 2550 2702 2553 2738
rect 2558 2702 2561 2728
rect 2582 2722 2585 2748
rect 2570 2718 2574 2721
rect 2590 2712 2593 2738
rect 2598 2732 2601 2748
rect 2606 2742 2609 2748
rect 2634 2738 2638 2741
rect 2614 2728 2622 2731
rect 2582 2692 2585 2698
rect 2598 2692 2601 2718
rect 2566 2552 2569 2608
rect 2574 2552 2577 2558
rect 2554 2548 2558 2551
rect 2594 2548 2598 2551
rect 2614 2551 2617 2728
rect 2638 2692 2641 2698
rect 2622 2642 2625 2658
rect 2646 2642 2649 2658
rect 2654 2631 2657 2778
rect 2670 2692 2673 2828
rect 2678 2772 2681 2908
rect 2678 2742 2681 2748
rect 2686 2742 2689 2858
rect 2670 2682 2673 2688
rect 2686 2682 2689 2738
rect 2682 2668 2686 2671
rect 2702 2662 2705 2938
rect 2726 2872 2729 2918
rect 2742 2761 2745 2898
rect 2750 2782 2753 2858
rect 2758 2771 2761 2938
rect 2770 2858 2774 2861
rect 2786 2858 2790 2861
rect 2766 2842 2769 2848
rect 2774 2792 2777 2848
rect 2790 2782 2793 2818
rect 2806 2772 2809 2878
rect 2830 2862 2833 3018
rect 2838 2952 2841 3008
rect 2862 2952 2865 2958
rect 2888 2903 2890 2907
rect 2894 2903 2897 2907
rect 2901 2903 2904 2907
rect 2858 2868 2862 2871
rect 2870 2862 2873 2868
rect 2818 2858 2822 2861
rect 2842 2858 2846 2861
rect 2854 2792 2857 2848
rect 2758 2768 2769 2771
rect 2742 2758 2758 2761
rect 2754 2748 2758 2751
rect 2766 2731 2769 2768
rect 2774 2742 2777 2748
rect 2782 2742 2785 2768
rect 2822 2762 2825 2778
rect 2794 2748 2798 2751
rect 2846 2742 2849 2768
rect 2862 2762 2865 2858
rect 2874 2748 2878 2751
rect 2790 2731 2793 2738
rect 2766 2728 2793 2731
rect 2814 2722 2817 2728
rect 2806 2712 2809 2718
rect 2742 2692 2745 2708
rect 2750 2682 2753 2688
rect 2766 2672 2769 2678
rect 2722 2658 2726 2661
rect 2702 2652 2705 2658
rect 2782 2652 2785 2659
rect 2730 2648 2734 2651
rect 2646 2628 2657 2631
rect 2646 2561 2649 2628
rect 2642 2558 2649 2561
rect 2614 2548 2622 2551
rect 2582 2532 2585 2538
rect 2622 2502 2625 2548
rect 2558 2482 2561 2488
rect 2534 2472 2537 2478
rect 2534 2452 2537 2468
rect 2574 2462 2577 2468
rect 2598 2462 2601 2488
rect 2542 2452 2545 2458
rect 2554 2428 2558 2431
rect 2554 2408 2561 2411
rect 2534 2392 2537 2398
rect 2558 2392 2561 2408
rect 2622 2392 2625 2448
rect 2638 2392 2641 2548
rect 2646 2392 2649 2558
rect 2666 2548 2670 2551
rect 2654 2492 2657 2548
rect 2678 2541 2681 2598
rect 2726 2552 2729 2558
rect 2734 2552 2737 2618
rect 2758 2552 2761 2558
rect 2698 2548 2702 2551
rect 2718 2542 2721 2548
rect 2766 2542 2769 2628
rect 2794 2558 2798 2561
rect 2794 2548 2798 2551
rect 2674 2538 2681 2541
rect 2670 2492 2673 2508
rect 2678 2472 2681 2528
rect 2694 2492 2697 2538
rect 2782 2532 2785 2538
rect 2746 2528 2750 2531
rect 2702 2472 2705 2488
rect 2662 2412 2665 2448
rect 2686 2432 2689 2468
rect 2694 2462 2697 2468
rect 2710 2462 2713 2468
rect 2718 2462 2721 2468
rect 2726 2462 2729 2478
rect 2734 2472 2737 2508
rect 2742 2482 2745 2518
rect 2782 2512 2785 2528
rect 2790 2492 2793 2538
rect 2806 2532 2809 2628
rect 2822 2592 2825 2618
rect 2798 2481 2801 2528
rect 2806 2522 2809 2528
rect 2790 2478 2801 2481
rect 2754 2468 2758 2471
rect 2754 2458 2758 2461
rect 2738 2428 2742 2431
rect 2766 2412 2769 2468
rect 2774 2462 2777 2478
rect 2662 2392 2665 2398
rect 2566 2352 2569 2388
rect 2606 2352 2609 2358
rect 2614 2352 2617 2368
rect 2554 2348 2558 2351
rect 2534 2312 2537 2338
rect 2542 2332 2545 2348
rect 2594 2328 2598 2331
rect 2566 2322 2569 2328
rect 2526 2298 2537 2301
rect 2482 2268 2486 2271
rect 2474 2258 2478 2261
rect 2494 2212 2497 2268
rect 2526 2262 2529 2288
rect 2534 2272 2537 2298
rect 2566 2262 2569 2268
rect 2510 2242 2513 2258
rect 2530 2238 2537 2241
rect 2502 2192 2505 2228
rect 2526 2212 2529 2218
rect 2462 2142 2465 2148
rect 2462 2112 2465 2138
rect 2470 2132 2473 2158
rect 2514 2148 2518 2151
rect 2466 2078 2470 2081
rect 2478 2061 2481 2118
rect 2486 2102 2489 2138
rect 2478 2058 2486 2061
rect 2494 2042 2497 2138
rect 2534 2122 2537 2238
rect 2550 2222 2553 2248
rect 2542 2192 2545 2198
rect 2506 2048 2510 2051
rect 2542 2042 2545 2118
rect 2454 1972 2457 2018
rect 2486 1972 2489 2018
rect 2474 1968 2478 1971
rect 2446 1902 2449 1958
rect 2502 1952 2505 1988
rect 2518 1952 2521 2008
rect 2550 1982 2553 2218
rect 2566 2192 2569 2258
rect 2574 2172 2577 2328
rect 2606 2272 2609 2308
rect 2614 2282 2617 2318
rect 2622 2312 2625 2378
rect 2630 2362 2633 2368
rect 2706 2358 2710 2361
rect 2646 2352 2649 2358
rect 2654 2352 2657 2358
rect 2638 2342 2641 2348
rect 2686 2342 2689 2348
rect 2726 2342 2729 2398
rect 2750 2392 2753 2408
rect 2782 2392 2785 2468
rect 2790 2462 2793 2478
rect 2830 2472 2833 2718
rect 2854 2702 2857 2718
rect 2862 2692 2865 2728
rect 2842 2688 2846 2691
rect 2878 2662 2881 2748
rect 2886 2732 2889 2738
rect 2888 2703 2890 2707
rect 2894 2703 2897 2707
rect 2901 2703 2904 2707
rect 2898 2658 2902 2661
rect 2902 2642 2905 2658
rect 2902 2552 2905 2638
rect 2910 2562 2913 3218
rect 2918 3142 2921 3218
rect 2926 3082 2929 3148
rect 2926 2992 2929 3058
rect 2934 2942 2937 3258
rect 2942 3252 2945 3258
rect 2990 3252 2993 3258
rect 2974 3242 2977 3248
rect 2950 3132 2953 3138
rect 2958 3132 2961 3158
rect 2970 3148 2974 3151
rect 2942 3052 2945 3118
rect 2982 3072 2985 3198
rect 2990 3152 2993 3158
rect 2998 3152 3001 3458
rect 3038 3412 3041 3438
rect 3102 3372 3105 3468
rect 3230 3462 3233 3518
rect 3238 3472 3241 3478
rect 3138 3458 3142 3461
rect 3210 3458 3214 3461
rect 3146 3448 3150 3451
rect 3182 3422 3185 3428
rect 3198 3422 3201 3458
rect 3246 3442 3249 3458
rect 3006 3352 3009 3368
rect 3070 3362 3073 3368
rect 3046 3352 3049 3358
rect 3126 3352 3129 3418
rect 3142 3352 3145 3368
rect 3166 3352 3169 3358
rect 3034 3348 3038 3351
rect 3082 3348 3086 3351
rect 3054 3342 3057 3348
rect 3042 3338 3046 3341
rect 3090 3338 3094 3341
rect 3206 3332 3209 3338
rect 3014 3292 3017 3318
rect 3086 3292 3089 3308
rect 3102 3292 3105 3298
rect 3062 3272 3065 3288
rect 3126 3272 3129 3278
rect 3006 3202 3009 3218
rect 3010 3168 3014 3171
rect 3046 3152 3049 3198
rect 3054 3152 3057 3158
rect 2998 3142 3001 3148
rect 3006 3102 3009 3148
rect 3070 3112 3073 3258
rect 3102 3222 3105 3248
rect 3118 3232 3121 3258
rect 3118 3202 3121 3228
rect 3126 3162 3129 3168
rect 3134 3142 3137 3228
rect 3142 3212 3145 3268
rect 3166 3262 3169 3298
rect 3142 3152 3145 3158
rect 3198 3152 3201 3158
rect 3178 3148 3182 3151
rect 3110 3132 3113 3138
rect 3166 3122 3169 3148
rect 3118 3092 3121 3118
rect 3022 3062 3025 3068
rect 2982 3042 2985 3058
rect 2942 2952 2945 3038
rect 3030 3032 3033 3058
rect 3054 3051 3057 3088
rect 3130 3068 3134 3071
rect 3062 3062 3065 3068
rect 3094 3062 3097 3068
rect 3082 3058 3086 3061
rect 3142 3052 3145 3058
rect 3050 3048 3057 3051
rect 3014 2992 3017 2998
rect 3030 2962 3033 3018
rect 3046 2992 3049 3018
rect 3070 3012 3073 3018
rect 2934 2901 2937 2938
rect 2926 2898 2937 2901
rect 2926 2772 2929 2898
rect 2942 2862 2945 2948
rect 2950 2942 2953 2958
rect 2990 2952 2993 2958
rect 2970 2948 2974 2951
rect 2998 2942 3001 2948
rect 3030 2932 3033 2948
rect 3070 2932 3073 2948
rect 2926 2752 2929 2758
rect 2918 2712 2921 2748
rect 2934 2742 2937 2758
rect 2918 2602 2921 2618
rect 2842 2548 2846 2551
rect 2882 2548 2886 2551
rect 2934 2541 2937 2718
rect 2942 2692 2945 2818
rect 2950 2762 2953 2918
rect 2966 2862 2969 2868
rect 2958 2752 2961 2758
rect 2950 2742 2953 2748
rect 2966 2712 2969 2748
rect 2990 2742 2993 2928
rect 3014 2881 3017 2918
rect 3014 2878 3025 2881
rect 3006 2802 3009 2868
rect 3014 2792 3017 2868
rect 2990 2692 2993 2738
rect 2998 2712 3001 2748
rect 2990 2662 2993 2668
rect 2998 2662 3001 2708
rect 3014 2692 3017 2778
rect 3022 2772 3025 2878
rect 3054 2862 3057 2868
rect 3030 2812 3033 2818
rect 3030 2692 3033 2808
rect 3038 2782 3041 2788
rect 3026 2668 3030 2671
rect 3002 2658 3006 2661
rect 2966 2652 2969 2658
rect 2946 2638 2950 2641
rect 2974 2572 2977 2618
rect 2954 2548 2958 2551
rect 2974 2542 2977 2558
rect 2982 2542 2985 2548
rect 2990 2542 2993 2618
rect 2998 2552 3001 2568
rect 3018 2558 3022 2561
rect 3034 2558 3038 2561
rect 3046 2552 3049 2828
rect 3078 2792 3081 3038
rect 3066 2748 3070 2751
rect 3078 2662 3081 2668
rect 3062 2642 3065 2658
rect 3086 2562 3089 3048
rect 3094 2942 3097 3048
rect 3158 3032 3161 3118
rect 3174 3072 3177 3138
rect 3182 3072 3185 3118
rect 3206 3102 3209 3148
rect 3214 3101 3217 3418
rect 3230 3392 3233 3418
rect 3230 3322 3233 3368
rect 3246 3342 3249 3398
rect 3254 3372 3257 3458
rect 3254 3342 3257 3348
rect 3222 3272 3225 3278
rect 3230 3262 3233 3318
rect 3238 3262 3241 3268
rect 3222 3172 3225 3218
rect 3222 3142 3225 3148
rect 3230 3141 3233 3258
rect 3238 3162 3241 3168
rect 3226 3138 3233 3141
rect 3214 3098 3225 3101
rect 3210 3088 3214 3091
rect 3202 3078 3206 3081
rect 3174 3032 3177 3058
rect 3106 3018 3110 3021
rect 3158 2962 3161 3018
rect 3174 3002 3177 3028
rect 3198 2982 3201 3018
rect 3146 2948 3150 2951
rect 3094 2862 3097 2868
rect 3126 2862 3129 2928
rect 3146 2888 3150 2891
rect 3098 2748 3102 2751
rect 3110 2692 3113 2808
rect 3126 2742 3129 2848
rect 3134 2792 3137 2878
rect 3158 2862 3161 2958
rect 3170 2868 3174 2871
rect 3182 2762 3185 2978
rect 3194 2968 3198 2971
rect 3222 2961 3225 3098
rect 3246 3062 3249 3338
rect 3254 3272 3257 3338
rect 3262 3262 3265 3508
rect 3278 3502 3281 3808
rect 3286 3742 3289 3758
rect 3326 3742 3329 3948
rect 3334 3862 3337 4028
rect 3342 3961 3345 3988
rect 3350 3971 3353 4058
rect 3358 4012 3361 4058
rect 3374 4002 3377 4148
rect 3350 3968 3361 3971
rect 3342 3958 3350 3961
rect 3346 3868 3350 3871
rect 3358 3862 3361 3968
rect 3366 3902 3369 3948
rect 3374 3942 3377 3988
rect 3382 3952 3385 4218
rect 3400 4203 3402 4207
rect 3406 4203 3409 4207
rect 3413 4203 3416 4207
rect 3406 4142 3409 4147
rect 3438 4092 3441 4258
rect 3446 4222 3449 4258
rect 3470 4172 3473 4218
rect 3478 4162 3481 4518
rect 3502 4462 3505 4478
rect 3542 4472 3545 4498
rect 3550 4492 3553 4538
rect 3566 4512 3569 4618
rect 3622 4592 3625 4658
rect 3638 4642 3641 4648
rect 3686 4642 3689 4748
rect 3710 4712 3713 4718
rect 3726 4622 3729 4748
rect 3734 4732 3737 4738
rect 3738 4688 3742 4691
rect 3750 4662 3753 4778
rect 3766 4742 3769 4938
rect 3774 4852 3777 4918
rect 3782 4892 3785 4948
rect 3822 4932 3825 4968
rect 3862 4962 3865 5018
rect 3982 4952 3985 5018
rect 3882 4948 3886 4951
rect 3826 4918 3830 4921
rect 3774 4762 3777 4848
rect 3798 4822 3801 4858
rect 3806 4802 3809 4868
rect 3870 4862 3873 4938
rect 3974 4912 3977 4948
rect 3982 4942 3985 4948
rect 3920 4903 3922 4907
rect 3926 4903 3929 4907
rect 3933 4903 3936 4907
rect 3850 4858 3854 4861
rect 3774 4712 3777 4748
rect 3758 4672 3761 4678
rect 3742 4652 3745 4658
rect 3750 4652 3753 4658
rect 3614 4562 3617 4568
rect 3682 4548 3686 4551
rect 3574 4542 3577 4548
rect 3654 4542 3657 4548
rect 3582 4482 3585 4488
rect 3598 4472 3601 4538
rect 3662 4532 3665 4548
rect 3670 4532 3673 4538
rect 3694 4502 3697 4548
rect 3702 4522 3705 4548
rect 3710 4542 3713 4548
rect 3726 4532 3729 4578
rect 3774 4552 3777 4658
rect 3790 4652 3793 4798
rect 3838 4772 3841 4848
rect 3906 4838 3910 4841
rect 3926 4832 3929 4868
rect 3934 4862 3937 4888
rect 3998 4872 4001 5018
rect 4006 4892 4009 4908
rect 3958 4862 3961 4868
rect 3950 4842 3953 4848
rect 3954 4838 3961 4841
rect 3814 4762 3817 4768
rect 3838 4742 3841 4768
rect 3866 4758 3870 4761
rect 3906 4758 3910 4761
rect 3846 4752 3849 4758
rect 3830 4712 3833 4718
rect 3798 4682 3801 4688
rect 3854 4682 3857 4738
rect 3862 4682 3865 4718
rect 3862 4662 3865 4668
rect 3870 4662 3873 4748
rect 3878 4742 3881 4748
rect 3886 4692 3889 4718
rect 3902 4702 3905 4758
rect 3920 4703 3922 4707
rect 3926 4703 3929 4707
rect 3933 4703 3936 4707
rect 3818 4658 3822 4661
rect 3790 4552 3793 4648
rect 3814 4602 3817 4638
rect 3822 4612 3825 4618
rect 3806 4552 3809 4558
rect 3814 4551 3817 4598
rect 3838 4562 3841 4588
rect 3826 4558 3830 4561
rect 3874 4558 3878 4561
rect 3814 4548 3822 4551
rect 3734 4542 3737 4548
rect 3674 4488 3678 4491
rect 3562 4468 3566 4471
rect 3486 4392 3489 4418
rect 3494 4322 3497 4418
rect 3494 4262 3497 4318
rect 3502 4272 3505 4428
rect 3518 4342 3521 4358
rect 3526 4352 3529 4458
rect 3534 4442 3537 4468
rect 3542 4462 3545 4468
rect 3614 4463 3617 4468
rect 3566 4452 3569 4458
rect 3534 4352 3537 4438
rect 3558 4362 3561 4368
rect 3546 4358 3550 4361
rect 3614 4352 3617 4388
rect 3554 4348 3558 4351
rect 3510 4332 3513 4338
rect 3486 4242 3489 4258
rect 3502 4152 3505 4178
rect 3510 4162 3513 4218
rect 3518 4162 3521 4338
rect 3526 4312 3529 4348
rect 3534 4282 3537 4348
rect 3542 4342 3545 4348
rect 3542 4292 3545 4328
rect 3550 4302 3553 4338
rect 3582 4272 3585 4318
rect 3622 4272 3625 4378
rect 3638 4342 3641 4348
rect 3630 4262 3633 4288
rect 3594 4258 3598 4261
rect 3610 4258 3614 4261
rect 3526 4252 3529 4258
rect 3550 4232 3553 4258
rect 3558 4252 3561 4258
rect 3558 4232 3561 4248
rect 3614 4222 3617 4248
rect 3630 4242 3633 4248
rect 3450 4138 3454 4141
rect 3450 4128 3454 4131
rect 3470 4112 3473 4148
rect 3478 4142 3481 4148
rect 3494 4112 3497 4138
rect 3390 4062 3393 4068
rect 3426 4059 3430 4062
rect 3454 4062 3457 4078
rect 3494 4062 3497 4098
rect 3502 4072 3505 4138
rect 3510 4092 3513 4148
rect 3526 4132 3529 4168
rect 3558 4142 3561 4147
rect 3542 4132 3545 4138
rect 3518 4082 3521 4118
rect 3502 4062 3505 4068
rect 3390 3992 3393 4048
rect 3400 4003 3402 4007
rect 3406 4003 3409 4007
rect 3413 4003 3416 4007
rect 3422 3962 3425 4008
rect 3434 3978 3438 3981
rect 3430 3952 3433 3958
rect 3386 3938 3390 3941
rect 3366 3832 3369 3848
rect 3358 3771 3361 3818
rect 3350 3768 3361 3771
rect 3286 3692 3289 3738
rect 3278 3462 3281 3468
rect 3286 3462 3289 3478
rect 3302 3452 3305 3658
rect 3318 3652 3321 3738
rect 3334 3732 3337 3747
rect 3342 3682 3345 3688
rect 3338 3668 3342 3671
rect 3350 3662 3353 3768
rect 3366 3742 3369 3748
rect 3374 3742 3377 3898
rect 3382 3892 3385 3938
rect 3402 3888 3406 3891
rect 3438 3872 3441 3918
rect 3382 3852 3385 3858
rect 3400 3803 3402 3807
rect 3406 3803 3409 3807
rect 3413 3803 3416 3807
rect 3446 3782 3449 3928
rect 3454 3922 3457 4058
rect 3470 3992 3473 4058
rect 3526 4032 3529 4128
rect 3542 4032 3545 4048
rect 3486 4012 3489 4018
rect 3462 3948 3470 3951
rect 3482 3948 3486 3951
rect 3462 3912 3465 3948
rect 3494 3941 3497 4018
rect 3506 3958 3510 3961
rect 3526 3952 3529 4018
rect 3514 3948 3518 3951
rect 3490 3938 3497 3941
rect 3530 3938 3534 3941
rect 3470 3932 3473 3938
rect 3542 3922 3545 3938
rect 3494 3882 3497 3918
rect 3526 3862 3529 3868
rect 3534 3862 3537 3888
rect 3542 3882 3545 3918
rect 3494 3852 3497 3859
rect 3542 3842 3545 3848
rect 3382 3742 3385 3748
rect 3390 3732 3393 3748
rect 3398 3732 3401 3778
rect 3474 3758 3478 3761
rect 3494 3752 3497 3838
rect 3502 3752 3505 3798
rect 3526 3752 3529 3778
rect 3482 3748 3486 3751
rect 3518 3748 3526 3751
rect 3414 3742 3417 3748
rect 3458 3738 3462 3741
rect 3450 3728 3454 3731
rect 3330 3658 3334 3661
rect 3310 3512 3313 3648
rect 3318 3642 3321 3648
rect 3318 3542 3321 3638
rect 3326 3592 3329 3618
rect 3326 3551 3329 3558
rect 3366 3552 3369 3658
rect 3358 3542 3361 3548
rect 3326 3472 3329 3528
rect 3322 3459 3326 3462
rect 3350 3432 3353 3458
rect 3366 3422 3369 3548
rect 3294 3392 3297 3408
rect 3318 3392 3321 3418
rect 3358 3362 3361 3368
rect 3274 3358 3278 3361
rect 3282 3348 3286 3351
rect 3334 3332 3337 3348
rect 3270 3302 3273 3318
rect 3294 3292 3297 3318
rect 3286 3272 3289 3288
rect 3318 3272 3321 3318
rect 3266 3258 3270 3261
rect 3254 3242 3257 3248
rect 3318 3182 3321 3268
rect 3326 3252 3329 3258
rect 3334 3252 3337 3328
rect 3342 3282 3345 3358
rect 3350 3282 3353 3348
rect 3358 3312 3361 3348
rect 3374 3342 3377 3688
rect 3458 3668 3462 3671
rect 3422 3663 3425 3668
rect 3470 3662 3473 3748
rect 3494 3712 3497 3738
rect 3502 3692 3505 3748
rect 3518 3732 3521 3748
rect 3550 3742 3553 4018
rect 3566 3992 3569 4128
rect 3574 3992 3577 4218
rect 3646 4191 3649 4328
rect 3662 4272 3665 4388
rect 3686 4362 3689 4478
rect 3702 4462 3705 4518
rect 3718 4492 3721 4518
rect 3734 4482 3737 4528
rect 3750 4491 3753 4528
rect 3774 4522 3777 4548
rect 3766 4512 3769 4518
rect 3746 4488 3753 4491
rect 3722 4468 3726 4471
rect 3694 4392 3697 4418
rect 3710 4412 3713 4458
rect 3734 4442 3737 4448
rect 3782 4382 3785 4538
rect 3790 4462 3793 4548
rect 3806 4532 3809 4538
rect 3814 4501 3817 4538
rect 3806 4498 3817 4501
rect 3798 4452 3801 4458
rect 3654 4262 3657 4268
rect 3638 4188 3649 4191
rect 3670 4242 3673 4248
rect 3618 4168 3622 4171
rect 3622 4112 3625 4158
rect 3638 4142 3641 4188
rect 3662 4152 3665 4158
rect 3606 4072 3609 4078
rect 3622 4072 3625 4108
rect 3638 4102 3641 4138
rect 3638 4082 3641 4098
rect 3590 4052 3593 4059
rect 3558 3862 3561 3968
rect 3598 3942 3601 4018
rect 3622 3992 3625 4068
rect 3670 4062 3673 4238
rect 3678 4072 3681 4298
rect 3686 4262 3689 4358
rect 3714 4348 3718 4351
rect 3766 4342 3769 4378
rect 3774 4358 3782 4361
rect 3774 4352 3777 4358
rect 3786 4348 3790 4351
rect 3770 4338 3774 4341
rect 3758 4272 3761 4338
rect 3798 4332 3801 4358
rect 3806 4342 3809 4498
rect 3822 4492 3825 4548
rect 3838 4482 3841 4558
rect 3874 4548 3878 4551
rect 3846 4542 3849 4548
rect 3854 4502 3857 4548
rect 3878 4512 3881 4538
rect 3846 4472 3849 4498
rect 3822 4462 3825 4468
rect 3838 4452 3841 4458
rect 3854 4392 3857 4488
rect 3862 4482 3865 4488
rect 3870 4472 3873 4478
rect 3878 4462 3881 4498
rect 3886 4472 3889 4548
rect 3902 4542 3905 4548
rect 3910 4542 3913 4678
rect 3922 4538 3926 4541
rect 3934 4532 3937 4618
rect 3942 4582 3945 4748
rect 3950 4742 3953 4768
rect 3958 4752 3961 4838
rect 3974 4822 3977 4858
rect 3982 4802 3985 4868
rect 3990 4842 3993 4858
rect 3990 4782 3993 4838
rect 3998 4782 4001 4868
rect 4014 4862 4017 5028
rect 4070 4962 4073 5068
rect 4082 5058 4086 5061
rect 4222 5062 4225 5068
rect 4206 5032 4209 5059
rect 4286 5042 4289 5058
rect 4310 5052 4313 5058
rect 4138 5018 4142 5021
rect 4246 4972 4249 5018
rect 4070 4952 4073 4958
rect 4138 4948 4142 4951
rect 4042 4918 4046 4921
rect 4030 4911 4033 4918
rect 4030 4908 4041 4911
rect 4038 4882 4041 4908
rect 4022 4862 4025 4868
rect 3978 4758 3982 4761
rect 3998 4742 4001 4768
rect 4006 4742 4009 4748
rect 3954 4738 3958 4741
rect 3990 4722 3993 4728
rect 3962 4668 3966 4671
rect 3990 4662 3993 4668
rect 3998 4662 4001 4728
rect 4014 4672 4017 4858
rect 4022 4792 4025 4848
rect 4038 4812 4041 4878
rect 4054 4872 4057 4918
rect 4094 4892 4097 4948
rect 4134 4932 4137 4938
rect 4158 4922 4161 4958
rect 4230 4952 4233 4958
rect 4170 4948 4174 4951
rect 4250 4948 4254 4951
rect 4102 4882 4105 4888
rect 4142 4882 4145 4918
rect 4122 4878 4126 4881
rect 4110 4872 4113 4878
rect 4046 4852 4049 4868
rect 4054 4862 4057 4868
rect 4086 4862 4089 4868
rect 4122 4858 4126 4861
rect 4146 4858 4150 4861
rect 4078 4852 4081 4858
rect 4046 4752 4049 4778
rect 4034 4748 4038 4751
rect 4046 4742 4049 4748
rect 4054 4691 4057 4818
rect 4070 4762 4073 4848
rect 4086 4782 4089 4858
rect 4062 4712 4065 4728
rect 4054 4688 4065 4691
rect 4014 4662 4017 4668
rect 4034 4658 4038 4661
rect 3990 4652 3993 4658
rect 3998 4632 4001 4658
rect 3950 4542 3953 4548
rect 3966 4542 3969 4568
rect 3982 4532 3985 4547
rect 3862 4362 3865 4418
rect 3878 4382 3881 4458
rect 3894 4442 3897 4448
rect 3902 4362 3905 4518
rect 3920 4503 3922 4507
rect 3926 4503 3929 4507
rect 3933 4503 3936 4507
rect 4006 4492 4009 4658
rect 3910 4472 3913 4478
rect 3942 4372 3945 4488
rect 3950 4392 3953 4458
rect 3890 4358 3894 4361
rect 3814 4342 3817 4348
rect 3766 4312 3769 4318
rect 3806 4302 3809 4338
rect 3822 4332 3825 4338
rect 3830 4332 3833 4358
rect 3838 4352 3841 4358
rect 3790 4272 3793 4298
rect 3730 4268 3734 4271
rect 3694 4262 3697 4268
rect 3714 4258 3718 4261
rect 3686 4132 3689 4258
rect 3702 4252 3705 4258
rect 3718 4092 3721 4248
rect 3726 4182 3729 4258
rect 3750 4252 3753 4258
rect 3734 4162 3737 4218
rect 3742 4142 3745 4148
rect 3710 4072 3713 4078
rect 3726 4072 3729 4138
rect 3758 4112 3761 4268
rect 3782 4262 3785 4268
rect 3766 4192 3769 4258
rect 3790 4252 3793 4258
rect 3822 4252 3825 4278
rect 3838 4262 3841 4308
rect 3846 4272 3849 4358
rect 3942 4352 3945 4368
rect 3890 4348 3894 4351
rect 3930 4348 3934 4351
rect 3858 4338 3862 4341
rect 3874 4338 3878 4341
rect 3870 4312 3873 4338
rect 3878 4282 3881 4318
rect 3902 4292 3905 4318
rect 3910 4292 3913 4328
rect 3920 4303 3922 4307
rect 3926 4303 3929 4307
rect 3933 4303 3936 4307
rect 3958 4282 3961 4468
rect 4014 4442 4017 4658
rect 4030 4642 4033 4648
rect 4042 4588 4046 4591
rect 4054 4552 4057 4678
rect 4062 4622 4065 4688
rect 4062 4562 4065 4568
rect 4070 4562 4073 4758
rect 4094 4752 4097 4848
rect 4102 4752 4105 4848
rect 4182 4822 4185 4948
rect 4190 4932 4193 4938
rect 4194 4918 4198 4921
rect 4206 4892 4209 4938
rect 4230 4882 4233 4948
rect 4190 4852 4193 4858
rect 4122 4788 4126 4791
rect 4134 4752 4137 4818
rect 4166 4792 4169 4818
rect 4082 4738 4086 4741
rect 4078 4652 4081 4718
rect 4094 4672 4097 4748
rect 4074 4558 4078 4561
rect 4086 4552 4089 4618
rect 4102 4592 4105 4748
rect 4134 4722 4137 4748
rect 4126 4682 4129 4688
rect 4142 4662 4145 4748
rect 4150 4732 4153 4748
rect 4158 4742 4161 4748
rect 4110 4642 4113 4658
rect 4118 4552 4121 4598
rect 4134 4562 4137 4578
rect 4142 4542 4145 4608
rect 4158 4582 4161 4618
rect 4166 4572 4169 4788
rect 4174 4611 4177 4808
rect 4182 4752 4185 4768
rect 4190 4742 4193 4748
rect 4206 4682 4209 4878
rect 4214 4862 4217 4868
rect 4230 4862 4233 4868
rect 4238 4862 4241 4898
rect 4246 4882 4249 4918
rect 4294 4902 4297 4948
rect 4302 4942 4305 4998
rect 4342 4992 4345 5028
rect 4358 4982 4361 5018
rect 4358 4952 4361 4968
rect 4318 4932 4321 4948
rect 4310 4912 4313 4918
rect 4282 4888 4286 4891
rect 4294 4882 4297 4888
rect 4326 4882 4329 4888
rect 4266 4878 4270 4881
rect 4286 4872 4289 4878
rect 4306 4868 4310 4871
rect 4270 4862 4273 4868
rect 4306 4858 4310 4861
rect 4214 4752 4217 4858
rect 4222 4852 4225 4858
rect 4238 4731 4241 4858
rect 4270 4852 4273 4858
rect 4318 4842 4321 4858
rect 4234 4728 4241 4731
rect 4214 4722 4217 4728
rect 4234 4718 4238 4721
rect 4222 4682 4225 4718
rect 4206 4672 4209 4678
rect 4174 4608 4185 4611
rect 4150 4552 4153 4558
rect 4054 4522 4057 4538
rect 4102 4532 4105 4538
rect 4110 4532 4113 4538
rect 4166 4532 4169 4548
rect 4174 4542 4177 4558
rect 4182 4532 4185 4608
rect 4222 4592 4225 4659
rect 4198 4542 4201 4548
rect 4194 4528 4198 4531
rect 4134 4522 4137 4528
rect 4206 4522 4209 4558
rect 4222 4552 4225 4558
rect 4230 4542 4233 4578
rect 4054 4472 4057 4518
rect 4094 4512 4097 4518
rect 4166 4482 4169 4518
rect 4102 4462 4105 4468
rect 4190 4462 4193 4468
rect 4026 4458 4030 4461
rect 4066 4458 4070 4461
rect 4094 4452 4097 4458
rect 3982 4362 3985 4418
rect 3970 4348 3974 4351
rect 3998 4332 4001 4348
rect 4006 4342 4009 4358
rect 4022 4352 4025 4418
rect 4046 4361 4049 4418
rect 4086 4372 4089 4418
rect 4094 4392 4097 4438
rect 4042 4358 4049 4361
rect 4030 4352 4033 4358
rect 4062 4352 4065 4358
rect 4082 4348 4086 4351
rect 4070 4342 4073 4348
rect 3970 4288 3974 4291
rect 3878 4263 3881 4268
rect 3910 4262 3913 4278
rect 3782 4242 3785 4248
rect 3774 4152 3777 4178
rect 3790 4162 3793 4248
rect 3798 4242 3801 4248
rect 3814 4222 3817 4248
rect 3798 4192 3801 4208
rect 3782 4122 3785 4148
rect 3790 4142 3793 4148
rect 3806 4132 3809 4158
rect 3766 4062 3769 4088
rect 3790 4072 3793 4098
rect 3814 4092 3817 4118
rect 3774 4062 3777 4068
rect 3634 4058 3638 4061
rect 3706 4058 3710 4061
rect 3722 4058 3729 4061
rect 3738 4058 3742 4061
rect 3630 4042 3633 4048
rect 3646 3992 3649 4038
rect 3654 4032 3657 4048
rect 3622 3962 3625 3968
rect 3606 3952 3609 3958
rect 3638 3952 3641 3958
rect 3670 3952 3673 4058
rect 3678 4022 3681 4058
rect 3710 4048 3718 4051
rect 3618 3948 3622 3951
rect 3662 3948 3670 3951
rect 3610 3938 3614 3941
rect 3582 3922 3585 3928
rect 3566 3882 3569 3908
rect 3574 3872 3577 3918
rect 3590 3902 3593 3918
rect 3614 3892 3617 3898
rect 3638 3892 3641 3938
rect 3586 3888 3590 3891
rect 3646 3882 3649 3948
rect 3662 3932 3665 3948
rect 3670 3902 3673 3938
rect 3558 3762 3561 3858
rect 3526 3732 3529 3738
rect 3510 3722 3513 3728
rect 3502 3662 3505 3678
rect 3510 3662 3513 3718
rect 3542 3712 3545 3728
rect 3526 3692 3529 3698
rect 3518 3672 3521 3688
rect 3550 3672 3553 3738
rect 3574 3692 3577 3868
rect 3650 3858 3654 3861
rect 3586 3848 3590 3851
rect 3598 3822 3601 3858
rect 3662 3792 3665 3878
rect 3678 3872 3681 3928
rect 3686 3892 3689 4048
rect 3694 3942 3697 3958
rect 3698 3868 3702 3871
rect 3678 3862 3681 3868
rect 3710 3862 3713 4048
rect 3726 4032 3729 4058
rect 3722 3958 3726 3961
rect 3722 3948 3726 3951
rect 3726 3932 3729 3938
rect 3726 3882 3729 3928
rect 3734 3922 3737 3938
rect 3750 3922 3753 4048
rect 3782 3952 3785 3958
rect 3790 3942 3793 4068
rect 3818 4058 3822 4061
rect 3626 3788 3630 3791
rect 3610 3748 3614 3751
rect 3658 3748 3662 3751
rect 3686 3751 3689 3818
rect 3702 3742 3705 3828
rect 3710 3812 3713 3858
rect 3718 3852 3721 3858
rect 3734 3842 3737 3918
rect 3742 3862 3745 3868
rect 3750 3822 3753 3838
rect 3782 3832 3785 3858
rect 3742 3818 3750 3821
rect 3718 3752 3721 3758
rect 3726 3742 3729 3778
rect 3570 3668 3574 3671
rect 3474 3658 3478 3661
rect 3390 3652 3393 3658
rect 3518 3651 3521 3668
rect 3558 3652 3561 3658
rect 3510 3648 3521 3651
rect 3400 3603 3402 3607
rect 3406 3603 3409 3607
rect 3413 3603 3416 3607
rect 3422 3602 3425 3618
rect 3390 3552 3393 3598
rect 3422 3552 3425 3598
rect 3478 3592 3481 3618
rect 3402 3548 3406 3551
rect 3430 3542 3433 3568
rect 3454 3552 3457 3588
rect 3466 3558 3470 3561
rect 3494 3552 3497 3558
rect 3502 3552 3505 3558
rect 3478 3542 3481 3548
rect 3502 3542 3505 3548
rect 3490 3538 3494 3541
rect 3446 3532 3449 3538
rect 3434 3518 3438 3521
rect 3402 3478 3406 3481
rect 3430 3462 3433 3488
rect 3446 3452 3449 3518
rect 3510 3462 3513 3648
rect 3534 3641 3537 3648
rect 3530 3638 3537 3641
rect 3518 3541 3521 3638
rect 3542 3592 3545 3618
rect 3574 3592 3577 3658
rect 3590 3642 3593 3648
rect 3590 3602 3593 3638
rect 3598 3622 3601 3668
rect 3610 3658 3614 3661
rect 3546 3558 3550 3561
rect 3530 3548 3534 3551
rect 3518 3538 3529 3541
rect 3538 3538 3542 3541
rect 3526 3492 3529 3538
rect 3590 3492 3593 3588
rect 3606 3542 3609 3548
rect 3542 3472 3545 3488
rect 3562 3478 3566 3481
rect 3550 3472 3553 3478
rect 3574 3472 3577 3488
rect 3606 3472 3609 3498
rect 3454 3432 3457 3458
rect 3518 3422 3521 3468
rect 3542 3462 3545 3468
rect 3566 3462 3569 3468
rect 3586 3458 3590 3461
rect 3400 3403 3402 3407
rect 3406 3403 3409 3407
rect 3413 3403 3416 3407
rect 3286 3151 3289 3158
rect 3358 3152 3361 3158
rect 3254 3142 3257 3148
rect 3270 3063 3273 3078
rect 3286 3072 3289 3128
rect 3302 3082 3305 3088
rect 3326 3072 3329 3078
rect 3214 2958 3225 2961
rect 3198 2952 3201 2958
rect 3202 2938 3206 2941
rect 3190 2862 3193 2888
rect 3198 2862 3201 2868
rect 3206 2862 3209 2928
rect 3206 2752 3209 2858
rect 3214 2761 3217 2958
rect 3230 2952 3233 2968
rect 3246 2952 3249 3018
rect 3254 2952 3257 2958
rect 3222 2942 3225 2948
rect 3230 2932 3233 2948
rect 3246 2942 3249 2948
rect 3270 2942 3273 2998
rect 3286 2942 3289 3068
rect 3318 3062 3321 3068
rect 3350 3062 3353 3068
rect 3330 3058 3334 3061
rect 3366 3061 3369 3288
rect 3382 3262 3385 3278
rect 3398 3242 3401 3278
rect 3414 3262 3417 3378
rect 3430 3362 3433 3418
rect 3526 3392 3529 3448
rect 3542 3432 3545 3438
rect 3482 3368 3486 3371
rect 3442 3348 3446 3351
rect 3422 3322 3425 3348
rect 3438 3282 3441 3308
rect 3446 3272 3449 3338
rect 3462 3291 3465 3358
rect 3542 3352 3545 3428
rect 3550 3352 3553 3358
rect 3458 3288 3465 3291
rect 3454 3272 3457 3288
rect 3470 3282 3473 3288
rect 3486 3272 3489 3348
rect 3534 3342 3537 3348
rect 3558 3342 3561 3458
rect 3590 3412 3593 3448
rect 3570 3358 3574 3361
rect 3586 3358 3590 3361
rect 3598 3352 3601 3368
rect 3590 3342 3593 3348
rect 3566 3332 3569 3338
rect 3598 3332 3601 3338
rect 3522 3318 3526 3321
rect 3558 3282 3561 3318
rect 3566 3292 3569 3328
rect 3582 3272 3585 3278
rect 3446 3262 3449 3268
rect 3470 3262 3473 3268
rect 3502 3263 3505 3268
rect 3534 3262 3537 3268
rect 3414 3232 3417 3258
rect 3430 3222 3433 3258
rect 3362 3058 3369 3061
rect 3302 2932 3305 2947
rect 3242 2928 3246 2931
rect 3222 2922 3225 2928
rect 3238 2872 3241 2888
rect 3246 2862 3249 2908
rect 3254 2851 3257 2918
rect 3286 2892 3289 2928
rect 3266 2888 3270 2891
rect 3278 2862 3281 2868
rect 3266 2858 3270 2861
rect 3254 2848 3262 2851
rect 3222 2842 3225 2848
rect 3214 2758 3222 2761
rect 3162 2748 3166 2751
rect 3234 2748 3238 2751
rect 3126 2622 3129 2738
rect 3150 2671 3153 2748
rect 3174 2722 3177 2728
rect 3150 2668 3158 2671
rect 3134 2662 3137 2668
rect 3158 2662 3161 2668
rect 3150 2642 3153 2658
rect 3166 2552 3169 2718
rect 3174 2602 3177 2618
rect 3174 2552 3177 2568
rect 3010 2548 3014 2551
rect 3130 2548 3134 2551
rect 2934 2538 2942 2541
rect 2838 2472 2841 2538
rect 2846 2502 2849 2538
rect 2890 2518 2894 2521
rect 2878 2492 2881 2508
rect 2888 2503 2890 2507
rect 2894 2503 2897 2507
rect 2901 2503 2904 2507
rect 2874 2478 2878 2481
rect 2850 2468 2854 2471
rect 2798 2462 2801 2468
rect 2862 2462 2865 2468
rect 2846 2452 2849 2458
rect 2834 2428 2838 2431
rect 2870 2421 2873 2478
rect 2878 2452 2881 2468
rect 2878 2432 2881 2448
rect 2894 2432 2897 2458
rect 2862 2418 2873 2421
rect 2790 2402 2793 2418
rect 2734 2352 2737 2368
rect 2750 2352 2753 2378
rect 2770 2358 2774 2361
rect 2670 2332 2673 2338
rect 2638 2302 2641 2318
rect 2662 2312 2665 2328
rect 2646 2292 2649 2298
rect 2678 2292 2681 2338
rect 2702 2292 2705 2328
rect 2626 2288 2630 2291
rect 2586 2258 2590 2261
rect 2630 2252 2633 2258
rect 2602 2168 2606 2171
rect 2654 2152 2657 2278
rect 2718 2272 2721 2318
rect 2726 2292 2729 2298
rect 2742 2282 2745 2338
rect 2774 2302 2777 2348
rect 2790 2332 2793 2368
rect 2798 2352 2801 2408
rect 2830 2352 2833 2358
rect 2846 2352 2849 2368
rect 2862 2362 2865 2418
rect 2834 2348 2838 2351
rect 2858 2348 2862 2351
rect 2870 2342 2873 2408
rect 2910 2352 2913 2538
rect 2926 2532 2929 2538
rect 2918 2472 2921 2508
rect 2926 2502 2929 2528
rect 2890 2348 2894 2351
rect 2846 2338 2854 2341
rect 2890 2338 2894 2341
rect 2806 2292 2809 2338
rect 2814 2332 2817 2338
rect 2822 2312 2825 2338
rect 2838 2302 2841 2338
rect 2846 2292 2849 2338
rect 2862 2292 2865 2318
rect 2888 2303 2890 2307
rect 2894 2303 2897 2307
rect 2901 2303 2904 2307
rect 2918 2292 2921 2368
rect 2926 2361 2929 2478
rect 2950 2472 2953 2538
rect 2958 2472 2961 2528
rect 2990 2492 2993 2528
rect 2974 2462 2977 2468
rect 2942 2452 2945 2458
rect 2950 2441 2953 2458
rect 2958 2452 2961 2458
rect 2982 2452 2985 2458
rect 2990 2452 2993 2468
rect 2942 2438 2953 2441
rect 2934 2412 2937 2418
rect 2926 2358 2934 2361
rect 2934 2352 2937 2358
rect 2926 2312 2929 2338
rect 2898 2288 2902 2291
rect 2854 2272 2857 2278
rect 2686 2262 2689 2268
rect 2694 2262 2697 2268
rect 2710 2262 2713 2268
rect 2666 2258 2670 2261
rect 2686 2248 2694 2251
rect 2718 2251 2721 2258
rect 2710 2248 2721 2251
rect 2726 2252 2729 2258
rect 2686 2192 2689 2248
rect 2710 2182 2713 2248
rect 2718 2192 2721 2228
rect 2734 2212 2737 2258
rect 2742 2232 2745 2258
rect 2742 2192 2745 2198
rect 2570 2148 2574 2151
rect 2626 2148 2630 2151
rect 2670 2142 2673 2148
rect 2702 2142 2705 2148
rect 2558 2132 2561 2138
rect 2558 2072 2561 2118
rect 2558 1972 2561 2068
rect 2574 2062 2577 2138
rect 2614 2132 2617 2138
rect 2622 2082 2625 2118
rect 2646 2102 2649 2118
rect 2574 2022 2577 2058
rect 2598 2052 2601 2058
rect 2630 2052 2633 2059
rect 2598 2032 2601 2048
rect 2566 2012 2569 2018
rect 2662 2012 2665 2068
rect 2678 2052 2681 2058
rect 2490 1948 2494 1951
rect 2470 1902 2473 1938
rect 2502 1932 2505 1938
rect 2446 1892 2449 1898
rect 2422 1862 2425 1878
rect 2438 1862 2441 1888
rect 2462 1882 2465 1888
rect 2366 1852 2369 1858
rect 2454 1842 2457 1868
rect 2470 1852 2473 1898
rect 2510 1892 2513 1928
rect 2478 1882 2481 1888
rect 2518 1882 2521 1948
rect 2530 1928 2534 1931
rect 2546 1928 2550 1931
rect 2486 1862 2489 1878
rect 2534 1862 2537 1928
rect 2558 1922 2561 1928
rect 2550 1918 2558 1921
rect 2550 1882 2553 1918
rect 2558 1882 2561 1888
rect 2434 1838 2438 1841
rect 2366 1792 2369 1808
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2397 1803 2400 1807
rect 2406 1762 2409 1818
rect 2486 1792 2489 1858
rect 2550 1852 2553 1878
rect 2566 1862 2569 1948
rect 2582 1932 2585 2008
rect 2694 1992 2697 2058
rect 2710 1992 2713 2068
rect 2718 2062 2721 2148
rect 2726 2031 2729 2138
rect 2734 2062 2737 2078
rect 2742 2072 2745 2118
rect 2750 2082 2753 2268
rect 2822 2262 2825 2268
rect 2786 2258 2790 2261
rect 2758 2212 2761 2258
rect 2766 2252 2769 2258
rect 2814 2192 2817 2248
rect 2830 2232 2833 2258
rect 2838 2192 2841 2268
rect 2862 2162 2865 2268
rect 2874 2258 2878 2261
rect 2870 2212 2873 2258
rect 2886 2252 2889 2268
rect 2934 2262 2937 2348
rect 2942 2292 2945 2438
rect 2982 2392 2985 2408
rect 2950 2312 2953 2358
rect 2990 2352 2993 2428
rect 2998 2362 3001 2548
rect 3018 2538 3022 2541
rect 3030 2532 3033 2548
rect 3078 2542 3081 2548
rect 3050 2538 3054 2541
rect 3006 2492 3009 2528
rect 3030 2492 3033 2518
rect 3038 2502 3041 2518
rect 3062 2492 3065 2528
rect 3070 2502 3073 2518
rect 3014 2472 3017 2488
rect 3086 2482 3089 2548
rect 3118 2542 3121 2548
rect 3106 2538 3110 2541
rect 3150 2532 3153 2548
rect 3174 2542 3177 2548
rect 3162 2538 3166 2541
rect 3102 2492 3105 2528
rect 3118 2522 3121 2528
rect 3006 2362 3009 2458
rect 3030 2352 3033 2378
rect 2966 2342 2969 2348
rect 2998 2342 3001 2348
rect 2986 2338 2990 2341
rect 3018 2338 3022 2341
rect 2974 2292 2977 2338
rect 3006 2322 3009 2338
rect 3022 2322 3025 2328
rect 3014 2312 3017 2318
rect 2962 2268 2966 2271
rect 2946 2258 2950 2261
rect 2886 2212 2889 2248
rect 2934 2192 2937 2258
rect 2990 2252 2993 2258
rect 3022 2252 3025 2258
rect 2942 2182 2945 2248
rect 3030 2222 3033 2348
rect 3038 2322 3041 2468
rect 3058 2458 3062 2461
rect 3054 2422 3057 2438
rect 3062 2352 3065 2418
rect 3070 2392 3073 2418
rect 3078 2371 3081 2458
rect 3070 2368 3081 2371
rect 3054 2332 3057 2348
rect 3046 2292 3049 2318
rect 3062 2312 3065 2338
rect 3070 2292 3073 2368
rect 3110 2362 3113 2518
rect 3118 2462 3121 2468
rect 3126 2452 3129 2458
rect 3134 2402 3137 2518
rect 3170 2468 3174 2471
rect 3150 2452 3153 2458
rect 3166 2442 3169 2448
rect 3142 2422 3145 2428
rect 3086 2342 3089 2358
rect 3126 2352 3129 2358
rect 3098 2348 3102 2351
rect 3114 2348 3118 2351
rect 3134 2342 3137 2368
rect 3094 2331 3097 2338
rect 3090 2328 3097 2331
rect 3126 2302 3129 2318
rect 3150 2272 3153 2428
rect 3162 2348 3166 2351
rect 3182 2351 3185 2718
rect 3198 2612 3201 2618
rect 3206 2601 3209 2738
rect 3214 2662 3217 2678
rect 3198 2598 3209 2601
rect 3190 2552 3193 2558
rect 3198 2551 3201 2598
rect 3210 2558 3214 2561
rect 3194 2548 3201 2551
rect 3222 2551 3225 2718
rect 3246 2702 3249 2718
rect 3238 2692 3241 2698
rect 3246 2562 3249 2698
rect 3254 2662 3257 2678
rect 3262 2662 3265 2748
rect 3270 2692 3273 2828
rect 3278 2792 3281 2798
rect 3302 2792 3305 2858
rect 3310 2761 3313 2938
rect 3334 2892 3337 3038
rect 3350 2942 3353 3058
rect 3358 3012 3361 3058
rect 3374 3052 3377 3148
rect 3390 3131 3393 3218
rect 3400 3203 3402 3207
rect 3406 3203 3409 3207
rect 3413 3203 3416 3207
rect 3422 3142 3425 3218
rect 3430 3182 3433 3218
rect 3426 3138 3430 3141
rect 3390 3128 3398 3131
rect 3390 3072 3393 3098
rect 3438 3082 3441 3198
rect 3450 3158 3454 3161
rect 3446 3132 3449 3148
rect 3462 3131 3465 3238
rect 3470 3152 3473 3208
rect 3510 3152 3513 3178
rect 3478 3142 3481 3148
rect 3474 3138 3478 3141
rect 3502 3141 3505 3148
rect 3550 3142 3553 3178
rect 3558 3152 3561 3258
rect 3590 3142 3593 3147
rect 3502 3138 3513 3141
rect 3458 3128 3465 3131
rect 3418 3068 3422 3071
rect 3382 3052 3385 3068
rect 3366 3042 3369 3048
rect 3390 2992 3393 3058
rect 3414 3052 3417 3058
rect 3400 3003 3402 3007
rect 3406 3003 3409 3007
rect 3413 3003 3416 3007
rect 3438 2972 3441 2988
rect 3378 2948 3382 2951
rect 3390 2942 3393 2948
rect 3370 2938 3374 2941
rect 3318 2872 3321 2878
rect 3338 2868 3342 2871
rect 3350 2862 3353 2888
rect 3366 2872 3369 2918
rect 3382 2862 3385 2928
rect 3414 2862 3417 2968
rect 3426 2938 3430 2941
rect 3446 2862 3449 3118
rect 3454 3062 3457 3088
rect 3454 3052 3457 3058
rect 3454 2992 3457 3038
rect 3426 2858 3430 2861
rect 3366 2852 3369 2858
rect 3322 2848 3326 2851
rect 3306 2758 3313 2761
rect 3302 2752 3305 2758
rect 3294 2662 3297 2668
rect 3310 2662 3313 2678
rect 3318 2662 3321 2668
rect 3310 2642 3313 2658
rect 3326 2592 3329 2838
rect 3334 2692 3337 2778
rect 3342 2672 3345 2728
rect 3294 2572 3297 2578
rect 3310 2552 3313 2558
rect 3342 2552 3345 2558
rect 3222 2548 3233 2551
rect 3242 2548 3246 2551
rect 3198 2542 3201 2548
rect 3218 2538 3222 2541
rect 3194 2528 3198 2531
rect 3190 2482 3193 2508
rect 3198 2482 3201 2508
rect 3190 2472 3193 2478
rect 3198 2461 3201 2468
rect 3194 2458 3201 2461
rect 3198 2402 3201 2418
rect 3214 2362 3217 2518
rect 3230 2511 3233 2548
rect 3254 2542 3257 2548
rect 3310 2542 3313 2548
rect 3254 2522 3257 2538
rect 3222 2508 3233 2511
rect 3222 2462 3225 2508
rect 3230 2472 3233 2498
rect 3230 2432 3233 2458
rect 3238 2431 3241 2508
rect 3262 2492 3265 2528
rect 3270 2502 3273 2518
rect 3326 2512 3329 2518
rect 3350 2482 3353 2828
rect 3390 2812 3393 2858
rect 3414 2851 3417 2858
rect 3414 2848 3425 2851
rect 3422 2812 3425 2848
rect 3462 2842 3465 3128
rect 3470 3062 3473 3068
rect 3478 3051 3481 3088
rect 3490 3068 3494 3071
rect 3474 3048 3481 3051
rect 3470 2892 3473 3008
rect 3478 2992 3481 3018
rect 3494 2992 3497 3018
rect 3510 2962 3513 3138
rect 3538 3138 3542 3141
rect 3526 3132 3529 3138
rect 3518 3122 3521 3128
rect 3534 3122 3537 3128
rect 3542 3063 3545 3078
rect 3558 3072 3561 3138
rect 3574 3072 3577 3078
rect 3558 3002 3561 3068
rect 3518 2972 3521 2978
rect 3562 2948 3566 2951
rect 3582 2951 3585 3108
rect 3598 3072 3601 3078
rect 3606 3072 3609 3468
rect 3614 3332 3617 3648
rect 3622 3632 3625 3668
rect 3630 3662 3633 3738
rect 3702 3672 3705 3738
rect 3726 3732 3729 3738
rect 3734 3712 3737 3718
rect 3658 3668 3662 3671
rect 3638 3662 3641 3668
rect 3650 3658 3654 3661
rect 3638 3612 3641 3648
rect 3670 3572 3673 3628
rect 3694 3552 3697 3668
rect 3710 3662 3713 3708
rect 3742 3632 3745 3818
rect 3750 3752 3753 3778
rect 3798 3771 3801 3988
rect 3830 3972 3833 4258
rect 3946 4218 3950 4221
rect 3982 4172 3985 4318
rect 4014 4212 4017 4338
rect 4058 4328 4062 4331
rect 4046 4312 4049 4328
rect 4062 4282 4065 4288
rect 4046 4272 4049 4278
rect 4030 4263 4033 4268
rect 4078 4262 4081 4268
rect 4094 4242 4097 4378
rect 4102 4352 4105 4448
rect 4150 4442 4153 4458
rect 4102 4292 4105 4348
rect 4110 4332 4113 4418
rect 4158 4392 4161 4428
rect 4134 4352 4137 4358
rect 4122 4348 4126 4351
rect 4146 4348 4150 4351
rect 4126 4332 4129 4338
rect 4134 4292 4137 4338
rect 4154 4268 4158 4271
rect 4110 4262 4113 4268
rect 4118 4262 4121 4268
rect 4166 4262 4169 4398
rect 4198 4372 4201 4438
rect 4230 4422 4233 4538
rect 4238 4532 4241 4708
rect 4254 4691 4257 4818
rect 4334 4802 4337 4948
rect 4366 4872 4369 4948
rect 4374 4922 4377 4928
rect 4378 4858 4382 4861
rect 4290 4748 4294 4751
rect 4318 4742 4321 4748
rect 4334 4742 4337 4748
rect 4390 4741 4393 5068
rect 4406 5062 4409 5068
rect 4590 5062 4593 5068
rect 4398 5032 4401 5058
rect 4406 4942 4409 5058
rect 4574 5052 4577 5059
rect 4474 5028 4481 5031
rect 4424 5003 4426 5007
rect 4430 5003 4433 5007
rect 4437 5003 4440 5007
rect 4406 4872 4409 4938
rect 4422 4862 4425 4968
rect 4430 4942 4433 4948
rect 4454 4932 4457 4938
rect 4446 4882 4449 4898
rect 4390 4738 4398 4741
rect 4342 4692 4345 4708
rect 4250 4688 4257 4691
rect 4278 4652 4281 4659
rect 4266 4558 4270 4561
rect 4286 4552 4289 4688
rect 4250 4528 4254 4531
rect 4206 4362 4209 4418
rect 4174 4352 4177 4358
rect 4238 4352 4241 4518
rect 4254 4472 4257 4478
rect 4262 4422 4265 4548
rect 4206 4342 4209 4348
rect 4230 4342 4233 4348
rect 4238 4342 4241 4348
rect 4178 4338 4182 4341
rect 4218 4338 4222 4341
rect 4046 4152 4049 4178
rect 4070 4172 4073 4178
rect 3866 4148 3870 4151
rect 3846 4102 3849 4148
rect 4034 4148 4038 4151
rect 3950 4111 3953 4147
rect 3942 4108 3953 4111
rect 3920 4103 3922 4107
rect 3926 4103 3929 4107
rect 3933 4103 3936 4107
rect 3886 4082 3889 4088
rect 3894 4078 3902 4081
rect 3894 4072 3897 4078
rect 3942 4072 3945 4108
rect 3958 4072 3961 4148
rect 3982 4092 3985 4138
rect 4038 4132 4041 4138
rect 4062 4132 4065 4158
rect 4094 4152 4097 4238
rect 4102 4152 4105 4168
rect 4086 4142 4089 4148
rect 4110 4141 4113 4248
rect 4150 4232 4153 4258
rect 4190 4252 4193 4318
rect 4210 4268 4214 4271
rect 4206 4252 4209 4258
rect 4230 4252 4233 4258
rect 4126 4152 4129 4158
rect 4106 4138 4113 4141
rect 4134 4132 4137 4218
rect 4166 4182 4169 4218
rect 4182 4202 4185 4248
rect 4150 4152 4153 4158
rect 4182 4152 4185 4158
rect 4158 4142 4161 4148
rect 4178 4138 4182 4141
rect 4062 4122 4065 4128
rect 3990 4062 3993 4068
rect 4006 4062 4009 4078
rect 4030 4062 4033 4088
rect 3910 4042 3913 4048
rect 3950 4042 3953 4058
rect 3862 3932 3865 3948
rect 3870 3872 3873 3878
rect 3910 3872 3913 3948
rect 3918 3942 3921 3968
rect 3950 3952 3953 4038
rect 3966 3962 3969 4058
rect 4006 3992 4009 4038
rect 4038 3992 4041 4108
rect 4046 4072 4049 4088
rect 4054 4062 4057 4068
rect 4046 3982 4049 4058
rect 3938 3948 3942 3951
rect 3970 3948 3974 3951
rect 3950 3942 3953 3948
rect 3990 3932 3993 3938
rect 3958 3922 3961 3928
rect 3920 3903 3922 3907
rect 3926 3903 3929 3907
rect 3933 3903 3936 3907
rect 3942 3892 3945 3898
rect 3974 3892 3977 3908
rect 3866 3868 3870 3871
rect 3914 3868 3918 3871
rect 3814 3852 3817 3859
rect 3858 3858 3862 3861
rect 3882 3858 3886 3861
rect 3846 3842 3849 3848
rect 3790 3768 3801 3771
rect 3774 3742 3777 3768
rect 3790 3762 3793 3768
rect 3806 3742 3809 3828
rect 3854 3802 3857 3858
rect 3874 3848 3878 3851
rect 3862 3842 3865 3848
rect 3830 3752 3833 3758
rect 3766 3691 3769 3728
rect 3762 3688 3769 3691
rect 3766 3662 3769 3688
rect 3774 3681 3777 3738
rect 3782 3702 3785 3718
rect 3786 3688 3790 3691
rect 3774 3678 3785 3681
rect 3794 3678 3830 3681
rect 3774 3652 3777 3668
rect 3782 3642 3785 3678
rect 3838 3671 3841 3688
rect 3826 3668 3841 3671
rect 3854 3672 3857 3788
rect 3890 3778 3894 3781
rect 3902 3752 3905 3858
rect 3910 3752 3913 3758
rect 3894 3742 3897 3748
rect 3902 3712 3905 3748
rect 3918 3732 3921 3858
rect 3950 3782 3953 3868
rect 3926 3772 3929 3778
rect 3958 3752 3961 3798
rect 3966 3742 3969 3878
rect 3974 3842 3977 3848
rect 3982 3792 3985 3818
rect 3998 3812 4001 3938
rect 4014 3932 4017 3958
rect 4054 3952 4057 4008
rect 4062 3992 4065 4098
rect 4070 4082 4073 4088
rect 4126 4072 4129 4118
rect 4142 4072 4145 4118
rect 4086 4062 4089 4068
rect 4110 4062 4113 4068
rect 4190 4062 4193 4168
rect 4198 4132 4201 4178
rect 4206 4172 4209 4218
rect 4222 4212 4225 4248
rect 4214 4142 4217 4158
rect 4226 4148 4230 4151
rect 4206 4112 4209 4118
rect 4198 4072 4201 4078
rect 4222 4062 4225 4088
rect 4230 4072 4233 4078
rect 4170 4058 4174 4061
rect 4210 4058 4214 4061
rect 4074 4048 4078 4051
rect 4086 3952 4089 4008
rect 4094 3992 4097 4018
rect 4118 3972 4121 4058
rect 4146 4048 4150 4051
rect 4110 3952 4113 3958
rect 4022 3942 4025 3948
rect 4078 3942 4081 3948
rect 4066 3928 4070 3931
rect 4086 3891 4089 3948
rect 4118 3942 4121 3948
rect 4078 3888 4089 3891
rect 3982 3782 3985 3788
rect 3990 3752 3993 3758
rect 3842 3658 3846 3661
rect 3798 3642 3801 3648
rect 3814 3582 3817 3618
rect 3822 3612 3825 3658
rect 3834 3648 3838 3651
rect 3706 3558 3710 3561
rect 3754 3558 3758 3561
rect 3726 3552 3729 3558
rect 3638 3542 3641 3548
rect 3622 3462 3625 3468
rect 3630 3462 3633 3498
rect 3626 3348 3630 3351
rect 3618 3328 3622 3331
rect 3638 3331 3641 3538
rect 3654 3521 3657 3538
rect 3678 3532 3681 3538
rect 3686 3522 3689 3548
rect 3630 3328 3641 3331
rect 3646 3518 3657 3521
rect 3666 3518 3670 3521
rect 3614 3262 3617 3268
rect 3630 3262 3633 3328
rect 3638 3312 3641 3318
rect 3646 3302 3649 3518
rect 3654 3341 3657 3418
rect 3662 3352 3665 3488
rect 3694 3462 3697 3548
rect 3734 3541 3737 3548
rect 3714 3538 3737 3541
rect 3774 3542 3777 3548
rect 3714 3528 3718 3531
rect 3758 3482 3761 3518
rect 3766 3492 3769 3518
rect 3806 3492 3809 3548
rect 3778 3468 3782 3471
rect 3706 3458 3710 3461
rect 3754 3458 3758 3461
rect 3798 3452 3801 3458
rect 3770 3438 3774 3441
rect 3710 3392 3713 3408
rect 3730 3358 3734 3361
rect 3694 3352 3697 3358
rect 3758 3352 3761 3398
rect 3814 3392 3817 3548
rect 3822 3462 3825 3598
rect 3886 3551 3889 3558
rect 3894 3542 3897 3668
rect 3902 3642 3905 3708
rect 3920 3703 3922 3707
rect 3926 3703 3929 3707
rect 3933 3703 3936 3707
rect 3950 3692 3953 3698
rect 3966 3692 3969 3738
rect 3994 3728 3998 3731
rect 4006 3731 4009 3798
rect 4014 3742 4017 3828
rect 4022 3752 4025 3758
rect 4030 3752 4033 3878
rect 4054 3792 4057 3858
rect 4062 3822 4065 3868
rect 4038 3752 4041 3778
rect 4078 3771 4081 3888
rect 4094 3832 4097 3868
rect 4106 3858 4110 3861
rect 4118 3852 4121 3868
rect 4126 3852 4129 3858
rect 4070 3768 4081 3771
rect 4070 3752 4073 3768
rect 4030 3742 4033 3748
rect 4110 3742 4113 3818
rect 4006 3728 4017 3731
rect 3974 3722 3977 3728
rect 3982 3722 3985 3728
rect 3974 3712 3977 3718
rect 4006 3712 4009 3718
rect 4006 3672 4009 3688
rect 3910 3632 3913 3658
rect 3966 3642 3969 3658
rect 3974 3642 3977 3668
rect 4014 3662 4017 3728
rect 4038 3672 4041 3698
rect 4038 3652 4041 3668
rect 4086 3662 4089 3668
rect 4102 3662 4105 3738
rect 4118 3692 4121 3748
rect 4054 3652 4057 3658
rect 4002 3648 4014 3651
rect 3950 3552 3953 3568
rect 3846 3518 3854 3521
rect 3846 3482 3849 3518
rect 3862 3482 3865 3488
rect 3894 3482 3897 3538
rect 3920 3503 3922 3507
rect 3926 3503 3929 3507
rect 3933 3503 3936 3507
rect 3950 3482 3953 3548
rect 3958 3492 3961 3558
rect 3766 3352 3769 3378
rect 3706 3348 3710 3351
rect 3678 3342 3681 3348
rect 3654 3338 3665 3341
rect 3662 3332 3665 3338
rect 3750 3332 3753 3338
rect 3782 3332 3785 3358
rect 3718 3292 3721 3308
rect 3670 3272 3673 3288
rect 3690 3268 3694 3271
rect 3718 3262 3721 3288
rect 3742 3272 3745 3328
rect 3782 3282 3785 3318
rect 3762 3278 3766 3281
rect 3730 3268 3734 3271
rect 3682 3258 3686 3261
rect 3738 3258 3745 3261
rect 3742 3242 3745 3258
rect 3774 3242 3777 3258
rect 3790 3242 3793 3348
rect 3798 3332 3801 3348
rect 3666 3238 3670 3241
rect 3706 3238 3710 3241
rect 3714 3238 3721 3241
rect 3686 3162 3689 3178
rect 3662 3142 3665 3148
rect 3654 3122 3657 3128
rect 3662 3092 3665 3098
rect 3630 3082 3633 3088
rect 3674 3078 3678 3081
rect 3710 3072 3713 3148
rect 3718 3132 3721 3238
rect 3742 3192 3745 3238
rect 3758 3202 3761 3218
rect 3790 3152 3793 3218
rect 3730 3148 3734 3151
rect 3798 3122 3801 3258
rect 3806 3242 3809 3258
rect 3814 3252 3817 3258
rect 3822 3242 3825 3458
rect 3846 3382 3849 3478
rect 3894 3421 3897 3459
rect 3922 3458 3926 3461
rect 3886 3418 3897 3421
rect 3854 3362 3857 3418
rect 3886 3392 3889 3418
rect 3902 3362 3905 3398
rect 3958 3362 3961 3418
rect 3866 3358 3870 3361
rect 3830 3352 3833 3358
rect 3950 3352 3953 3358
rect 3966 3352 3969 3638
rect 3986 3628 3990 3631
rect 4046 3622 4049 3628
rect 3990 3572 3993 3578
rect 3974 3532 3977 3558
rect 3990 3552 3993 3558
rect 3998 3542 4001 3568
rect 4022 3562 4025 3568
rect 4010 3558 4014 3561
rect 4034 3558 4038 3561
rect 4054 3552 4057 3578
rect 4062 3572 4065 3658
rect 4094 3622 4097 3658
rect 4102 3642 4105 3658
rect 4078 3612 4081 3618
rect 4126 3602 4129 3848
rect 4134 3792 4137 4018
rect 4150 3942 4153 3947
rect 4142 3872 4145 3908
rect 4158 3862 4161 4058
rect 4174 4042 4177 4048
rect 4182 4032 4185 4058
rect 4238 4042 4241 4338
rect 4250 4328 4254 4331
rect 4246 4272 4249 4318
rect 4270 4272 4273 4538
rect 4286 4492 4289 4538
rect 4350 4522 4353 4658
rect 4358 4542 4361 4738
rect 4366 4682 4369 4688
rect 4382 4672 4385 4678
rect 4390 4662 4393 4668
rect 4398 4632 4401 4738
rect 4406 4712 4409 4838
rect 4426 4818 4430 4821
rect 4424 4803 4426 4807
rect 4430 4803 4433 4807
rect 4437 4803 4440 4807
rect 4414 4762 4417 4768
rect 4446 4762 4449 4878
rect 4454 4752 4457 4788
rect 4406 4662 4409 4708
rect 4430 4702 4433 4748
rect 4418 4688 4422 4691
rect 4454 4662 4457 4738
rect 4462 4662 4465 4738
rect 4470 4732 4473 5018
rect 4478 5002 4481 5028
rect 4514 5018 4518 5021
rect 4478 4952 4481 4998
rect 4494 4952 4497 4958
rect 4478 4902 4481 4938
rect 4486 4882 4489 4928
rect 4494 4862 4497 4868
rect 4494 4752 4497 4758
rect 4486 4732 4489 4738
rect 4478 4722 4481 4728
rect 4294 4512 4297 4518
rect 4318 4472 4321 4508
rect 4278 4432 4281 4458
rect 4286 4351 4289 4358
rect 4302 4342 4305 4468
rect 4350 4462 4353 4498
rect 4358 4462 4361 4508
rect 4374 4492 4377 4547
rect 4390 4462 4393 4568
rect 4398 4472 4401 4488
rect 4406 4481 4409 4658
rect 4470 4652 4473 4718
rect 4478 4662 4481 4668
rect 4424 4603 4426 4607
rect 4430 4603 4433 4607
rect 4437 4603 4440 4607
rect 4502 4602 4505 5018
rect 4566 4992 4569 5038
rect 4514 4958 4518 4961
rect 4526 4951 4529 4978
rect 4522 4948 4529 4951
rect 4526 4902 4529 4938
rect 4542 4932 4545 4958
rect 4558 4952 4561 4978
rect 4606 4972 4609 5018
rect 4606 4952 4609 4958
rect 4534 4762 4537 4918
rect 4542 4902 4545 4928
rect 4570 4868 4574 4871
rect 4582 4862 4585 4948
rect 4590 4942 4593 4948
rect 4606 4862 4609 4948
rect 4638 4942 4641 4948
rect 4646 4892 4649 4908
rect 4550 4802 4553 4818
rect 4514 4758 4518 4761
rect 4550 4752 4553 4758
rect 4566 4752 4569 4858
rect 4606 4852 4609 4858
rect 4518 4732 4521 4738
rect 4510 4702 4513 4718
rect 4526 4692 4529 4718
rect 4534 4682 4537 4688
rect 4566 4682 4569 4748
rect 4574 4742 4577 4748
rect 4582 4732 4585 4768
rect 4614 4752 4617 4858
rect 4630 4852 4633 4858
rect 4630 4792 4633 4848
rect 4654 4792 4657 4938
rect 4670 4772 4673 5059
rect 4686 5042 4689 5068
rect 4782 5062 4785 5068
rect 4694 4932 4697 4938
rect 4678 4882 4681 4918
rect 4686 4842 4689 4858
rect 4694 4852 4697 4858
rect 4638 4752 4641 4758
rect 4630 4722 4633 4738
rect 4518 4672 4521 4678
rect 4550 4672 4553 4678
rect 4574 4672 4577 4718
rect 4626 4688 4630 4691
rect 4646 4672 4649 4748
rect 4678 4742 4681 4748
rect 4686 4742 4689 4788
rect 4702 4752 4705 5018
rect 4714 4948 4718 4951
rect 4742 4942 4745 4948
rect 4758 4932 4761 4998
rect 4722 4868 4726 4871
rect 4710 4752 4713 4778
rect 4734 4772 4737 4818
rect 4742 4752 4745 4758
rect 4698 4728 4702 4731
rect 4642 4668 4646 4671
rect 4522 4658 4526 4661
rect 4526 4612 4529 4658
rect 4566 4652 4569 4659
rect 4430 4552 4433 4558
rect 4486 4552 4489 4558
rect 4450 4548 4454 4551
rect 4506 4548 4510 4551
rect 4494 4542 4497 4548
rect 4414 4492 4417 4518
rect 4462 4492 4465 4538
rect 4470 4522 4473 4528
rect 4406 4478 4417 4481
rect 4442 4478 4446 4481
rect 4322 4458 4326 4461
rect 4330 4448 4334 4451
rect 4342 4402 4345 4448
rect 4382 4392 4385 4458
rect 4398 4361 4401 4468
rect 4406 4372 4409 4418
rect 4398 4358 4409 4361
rect 4394 4348 4398 4351
rect 4374 4342 4377 4348
rect 4394 4338 4398 4341
rect 4302 4282 4305 4338
rect 4350 4322 4353 4328
rect 4358 4322 4361 4328
rect 4334 4282 4337 4288
rect 4314 4278 4318 4281
rect 4258 4268 4262 4271
rect 4282 4268 4286 4271
rect 4290 4258 4294 4261
rect 4246 4152 4249 4258
rect 4262 4252 4265 4258
rect 4278 4252 4281 4258
rect 4262 4192 4265 4218
rect 4262 4062 4265 4068
rect 4278 4062 4281 4108
rect 4286 4102 4289 4258
rect 4294 4242 4297 4248
rect 4302 4182 4305 4278
rect 4350 4272 4353 4318
rect 4374 4302 4377 4338
rect 4406 4312 4409 4358
rect 4414 4352 4417 4478
rect 4462 4472 4465 4488
rect 4424 4403 4426 4407
rect 4430 4403 4433 4407
rect 4437 4403 4440 4407
rect 4322 4258 4326 4261
rect 4354 4258 4361 4261
rect 4302 4142 4305 4148
rect 4326 4142 4329 4178
rect 4350 4172 4353 4218
rect 4358 4192 4361 4258
rect 4366 4252 4369 4258
rect 4374 4192 4377 4278
rect 4406 4272 4409 4308
rect 4414 4302 4417 4348
rect 4426 4318 4430 4321
rect 4414 4272 4417 4278
rect 4398 4262 4401 4268
rect 4406 4262 4409 4268
rect 4446 4262 4449 4318
rect 4470 4292 4473 4518
rect 4494 4492 4497 4538
rect 4506 4518 4510 4521
rect 4478 4462 4481 4478
rect 4506 4468 4510 4471
rect 4518 4462 4521 4468
rect 4526 4462 4529 4588
rect 4550 4552 4553 4558
rect 4574 4542 4577 4668
rect 4642 4658 4646 4661
rect 4666 4658 4670 4661
rect 4666 4648 4670 4651
rect 4614 4552 4617 4648
rect 4646 4601 4649 4618
rect 4646 4598 4654 4601
rect 4638 4562 4641 4588
rect 4626 4558 4630 4561
rect 4534 4482 4537 4488
rect 4574 4462 4577 4468
rect 4482 4348 4486 4351
rect 4494 4272 4497 4458
rect 4526 4401 4529 4458
rect 4526 4398 4537 4401
rect 4510 4332 4513 4338
rect 4522 4318 4526 4321
rect 4526 4282 4529 4288
rect 4518 4272 4521 4278
rect 4522 4268 4529 4271
rect 4422 4252 4425 4258
rect 4346 4158 4350 4161
rect 4366 4152 4369 4168
rect 4362 4138 4366 4141
rect 4382 4122 4385 4248
rect 4424 4203 4426 4207
rect 4430 4203 4433 4207
rect 4437 4203 4440 4207
rect 4390 4172 4393 4178
rect 4430 4142 4433 4148
rect 4454 4142 4457 4258
rect 4310 4092 4313 4118
rect 4374 4112 4377 4118
rect 4342 4082 4345 4108
rect 4390 4092 4393 4138
rect 4494 4112 4497 4268
rect 4518 4152 4521 4158
rect 4330 4078 4334 4081
rect 4290 4068 4294 4071
rect 4326 4062 4329 4068
rect 4254 4052 4257 4058
rect 4266 4048 4270 4051
rect 4294 4022 4297 4058
rect 4222 3952 4225 3958
rect 4166 3912 4169 3938
rect 4238 3922 4241 4018
rect 4246 3952 4249 3998
rect 4258 3958 4262 3961
rect 4290 3948 4294 3951
rect 4230 3882 4233 3908
rect 4154 3828 4158 3831
rect 4198 3792 4201 3868
rect 4222 3852 4225 3858
rect 4230 3822 4233 3878
rect 4174 3782 4177 3788
rect 4134 3692 4137 3778
rect 4166 3722 4169 3728
rect 4134 3662 4137 3688
rect 4166 3672 4169 3688
rect 4158 3662 4161 3668
rect 4174 3652 4177 3768
rect 4182 3722 4185 3728
rect 4198 3672 4201 3778
rect 4210 3748 4214 3751
rect 4230 3742 4233 3818
rect 4246 3712 4249 3948
rect 4270 3942 4273 3948
rect 4302 3932 4305 3948
rect 4310 3942 4313 3948
rect 4326 3922 4329 4058
rect 4334 3952 4337 4028
rect 4350 4002 4353 4068
rect 4358 4062 4361 4088
rect 4378 4078 4382 4081
rect 4398 4072 4401 4108
rect 4518 4092 4521 4118
rect 4526 4072 4529 4268
rect 4534 4092 4537 4398
rect 4558 4332 4561 4338
rect 4542 4262 4545 4308
rect 4582 4272 4585 4478
rect 4590 4472 4593 4538
rect 4606 4532 4609 4538
rect 4630 4482 4633 4518
rect 4630 4452 4633 4458
rect 4630 4352 4633 4378
rect 4638 4362 4641 4518
rect 4646 4492 4649 4588
rect 4654 4542 4657 4548
rect 4646 4372 4649 4418
rect 4654 4382 4657 4458
rect 4662 4452 4665 4558
rect 4670 4522 4673 4528
rect 4666 4448 4670 4451
rect 4650 4358 4654 4361
rect 4590 4342 4593 4347
rect 4670 4342 4673 4348
rect 4590 4282 4593 4328
rect 4606 4292 4609 4338
rect 4622 4332 4625 4338
rect 4594 4268 4598 4271
rect 4578 4258 4582 4261
rect 4594 4258 4598 4261
rect 4550 4241 4553 4258
rect 4562 4248 4566 4251
rect 4550 4238 4561 4241
rect 4558 4182 4561 4238
rect 4570 4168 4574 4171
rect 4598 4142 4601 4148
rect 4606 4142 4609 4148
rect 4614 4142 4617 4308
rect 4622 4282 4625 4318
rect 4646 4302 4649 4318
rect 4642 4288 4646 4291
rect 4654 4291 4657 4328
rect 4650 4288 4657 4291
rect 4638 4262 4641 4268
rect 4662 4242 4665 4278
rect 4646 4192 4649 4228
rect 4634 4148 4638 4151
rect 4618 4138 4622 4141
rect 4634 4138 4638 4141
rect 4630 4092 4633 4098
rect 4394 4068 4398 4071
rect 4618 4068 4622 4071
rect 4382 4052 4385 4068
rect 4410 4058 4414 4061
rect 4454 4052 4457 4059
rect 4370 4048 4374 4051
rect 4358 3992 4361 4048
rect 4424 4003 4426 4007
rect 4430 4003 4433 4007
rect 4437 4003 4440 4007
rect 4270 3862 4273 3868
rect 4206 3691 4209 3698
rect 4206 3688 4214 3691
rect 4190 3662 4193 3668
rect 4206 3662 4209 3678
rect 4222 3672 4225 3678
rect 4186 3658 4190 3661
rect 4142 3632 4145 3648
rect 4162 3638 4166 3641
rect 4102 3552 4105 3578
rect 4026 3548 4030 3551
rect 4090 3548 4094 3551
rect 4114 3548 4118 3551
rect 4062 3542 4065 3548
rect 4030 3531 4033 3538
rect 4026 3528 4033 3531
rect 4046 3532 4049 3538
rect 4070 3532 4073 3548
rect 3990 3492 3993 3518
rect 4022 3482 4025 3488
rect 3998 3472 4001 3478
rect 4042 3468 4046 3471
rect 4062 3462 4065 3468
rect 4070 3462 4073 3468
rect 3982 3412 3985 3458
rect 3998 3452 4001 3458
rect 3982 3392 3985 3398
rect 3850 3348 3854 3351
rect 3906 3348 3910 3351
rect 3886 3342 3889 3348
rect 3834 3338 3838 3341
rect 3918 3341 3921 3348
rect 4014 3342 4017 3458
rect 3910 3338 3921 3341
rect 3970 3338 3974 3341
rect 3886 3332 3889 3338
rect 3830 3292 3833 3328
rect 3846 3262 3849 3318
rect 3874 3268 3878 3271
rect 3886 3262 3889 3288
rect 3854 3162 3857 3218
rect 3862 3161 3865 3218
rect 3894 3162 3897 3338
rect 3910 3292 3913 3338
rect 3942 3312 3945 3338
rect 3954 3328 3958 3331
rect 3920 3303 3922 3307
rect 3926 3303 3929 3307
rect 3933 3303 3936 3307
rect 4014 3292 4017 3338
rect 3990 3282 3993 3288
rect 4022 3282 4025 3418
rect 4030 3342 4033 3458
rect 4086 3442 4089 3528
rect 4094 3522 4097 3538
rect 4118 3502 4121 3518
rect 4126 3492 4129 3538
rect 3942 3262 3945 3278
rect 3990 3263 3993 3268
rect 4022 3262 4025 3268
rect 3918 3252 3921 3258
rect 3862 3158 3873 3161
rect 3810 3148 3814 3151
rect 3858 3148 3862 3151
rect 3838 3142 3841 3148
rect 3758 3082 3761 3088
rect 3766 3082 3769 3088
rect 3610 3068 3614 3071
rect 3658 3068 3662 3071
rect 3674 3068 3678 3071
rect 3590 3062 3593 3068
rect 3718 3062 3721 3078
rect 3750 3062 3753 3068
rect 3626 3058 3630 3061
rect 3642 3058 3646 3061
rect 3690 3058 3694 3061
rect 3590 3032 3593 3058
rect 3626 3048 3630 3051
rect 3706 3048 3710 3051
rect 3718 3042 3721 3048
rect 3578 2948 3585 2951
rect 3478 2942 3481 2948
rect 3534 2942 3537 2948
rect 3494 2872 3497 2918
rect 3510 2892 3513 2918
rect 3522 2888 3526 2891
rect 3462 2822 3465 2838
rect 3494 2822 3497 2858
rect 3526 2852 3529 2868
rect 3534 2822 3537 2938
rect 3574 2932 3577 2948
rect 3598 2942 3601 2998
rect 3678 2972 3681 3028
rect 3642 2948 3646 2951
rect 3550 2902 3553 2918
rect 3566 2892 3569 2918
rect 3542 2872 3545 2888
rect 3550 2872 3553 2888
rect 3558 2872 3561 2878
rect 3590 2872 3593 2918
rect 3542 2852 3545 2858
rect 3574 2852 3577 2868
rect 3590 2862 3593 2868
rect 3630 2862 3633 2938
rect 3642 2888 3646 2891
rect 3582 2852 3585 2858
rect 3400 2803 3402 2807
rect 3406 2803 3409 2807
rect 3413 2803 3416 2807
rect 3418 2748 3422 2751
rect 3390 2742 3393 2748
rect 3358 2732 3361 2738
rect 3390 2732 3393 2738
rect 3382 2642 3385 2658
rect 3430 2642 3433 2658
rect 3398 2622 3401 2628
rect 3400 2603 3402 2607
rect 3406 2603 3409 2607
rect 3413 2603 3416 2607
rect 3374 2552 3377 2558
rect 3382 2552 3385 2568
rect 3406 2552 3409 2558
rect 3390 2542 3393 2548
rect 3358 2502 3361 2518
rect 3250 2478 3254 2481
rect 3274 2478 3278 2481
rect 3294 2472 3297 2478
rect 3326 2472 3329 2478
rect 3358 2472 3361 2478
rect 3374 2472 3377 2478
rect 3406 2472 3409 2528
rect 3338 2468 3342 2471
rect 3254 2452 3257 2458
rect 3238 2428 3246 2431
rect 3234 2418 3238 2421
rect 3246 2361 3249 2428
rect 3254 2372 3257 2408
rect 3238 2358 3249 2361
rect 3238 2352 3241 2358
rect 3178 2348 3185 2351
rect 3250 2348 3254 2351
rect 3198 2342 3201 2348
rect 3158 2332 3161 2338
rect 3166 2332 3169 2338
rect 3182 2292 3185 2338
rect 3194 2328 3198 2331
rect 3114 2268 3118 2271
rect 3098 2258 3126 2261
rect 3134 2261 3137 2268
rect 3130 2258 3137 2261
rect 3158 2262 3161 2268
rect 3198 2262 3201 2318
rect 3206 2292 3209 2348
rect 3214 2272 3217 2348
rect 3222 2332 3225 2338
rect 3238 2332 3241 2348
rect 3270 2342 3273 2468
rect 3286 2352 3289 2418
rect 3294 2362 3297 2468
rect 3302 2462 3305 2468
rect 3338 2458 3342 2461
rect 3354 2458 3358 2461
rect 3266 2328 3270 2331
rect 3226 2298 3233 2301
rect 3230 2262 3233 2298
rect 3278 2292 3281 2348
rect 3286 2312 3289 2348
rect 3294 2332 3297 2348
rect 3302 2321 3305 2448
rect 3318 2442 3321 2458
rect 3318 2352 3321 2378
rect 3358 2362 3361 2388
rect 3366 2382 3369 2468
rect 3354 2358 3358 2361
rect 3334 2352 3337 2358
rect 3366 2352 3369 2358
rect 3374 2352 3377 2398
rect 3382 2352 3385 2458
rect 3398 2452 3401 2458
rect 3438 2412 3441 2818
rect 3470 2762 3473 2768
rect 3478 2752 3481 2788
rect 3446 2692 3449 2708
rect 3454 2662 3457 2678
rect 3454 2542 3457 2628
rect 3470 2592 3473 2738
rect 3478 2712 3481 2748
rect 3494 2732 3497 2758
rect 3506 2748 3510 2751
rect 3522 2748 3526 2751
rect 3502 2738 3518 2741
rect 3454 2522 3457 2538
rect 3478 2532 3481 2708
rect 3494 2672 3497 2728
rect 3502 2712 3505 2738
rect 3542 2732 3545 2738
rect 3514 2678 3518 2681
rect 3522 2668 3526 2671
rect 3542 2662 3545 2668
rect 3558 2662 3561 2818
rect 3606 2762 3609 2818
rect 3622 2802 3625 2858
rect 3654 2842 3657 2948
rect 3638 2792 3641 2798
rect 3650 2778 3654 2781
rect 3566 2752 3569 2758
rect 3678 2752 3681 2858
rect 3678 2732 3681 2748
rect 3602 2668 3609 2671
rect 3590 2662 3593 2668
rect 3606 2662 3609 2668
rect 3614 2662 3617 2668
rect 3554 2658 3558 2661
rect 3486 2642 3489 2658
rect 3542 2642 3545 2648
rect 3486 2552 3489 2638
rect 3622 2622 3625 2698
rect 3662 2692 3665 2728
rect 3686 2712 3689 3018
rect 3734 3002 3737 3048
rect 3742 2992 3745 3058
rect 3782 3032 3785 3068
rect 3806 3062 3809 3078
rect 3846 3062 3849 3068
rect 3814 2992 3817 3028
rect 3714 2988 3718 2991
rect 3694 2852 3697 2858
rect 3686 2682 3689 2688
rect 3654 2662 3657 2668
rect 3666 2658 3670 2661
rect 3646 2652 3649 2658
rect 3502 2592 3505 2618
rect 3566 2602 3569 2618
rect 3554 2598 3561 2601
rect 3558 2562 3561 2598
rect 3582 2552 3585 2568
rect 3486 2542 3489 2548
rect 3518 2542 3521 2548
rect 3570 2538 3574 2541
rect 3598 2532 3601 2538
rect 3542 2522 3545 2528
rect 3630 2522 3633 2618
rect 3638 2542 3641 2548
rect 3678 2542 3681 2548
rect 3618 2518 3622 2521
rect 3446 2492 3449 2498
rect 3486 2472 3489 2478
rect 3542 2472 3545 2518
rect 3550 2472 3553 2478
rect 3514 2468 3518 2471
rect 3494 2462 3497 2468
rect 3526 2462 3529 2468
rect 3446 2422 3449 2458
rect 3400 2403 3402 2407
rect 3406 2403 3409 2407
rect 3413 2403 3416 2407
rect 3394 2358 3398 2361
rect 3350 2342 3353 2348
rect 3338 2338 3342 2341
rect 3326 2332 3329 2338
rect 3294 2318 3305 2321
rect 3286 2292 3289 2298
rect 3266 2288 3270 2291
rect 3242 2268 3246 2271
rect 3086 2222 3089 2258
rect 3010 2218 3014 2221
rect 3178 2218 3182 2221
rect 3046 2212 3049 2218
rect 2758 2142 2761 2148
rect 2766 2142 2769 2148
rect 2782 2142 2785 2148
rect 2834 2138 2841 2141
rect 2758 2082 2761 2118
rect 2766 2112 2769 2138
rect 2782 2132 2785 2138
rect 2814 2102 2817 2118
rect 2838 2082 2841 2138
rect 2738 2058 2742 2061
rect 2774 2032 2777 2068
rect 2814 2062 2817 2078
rect 2822 2072 2825 2078
rect 2726 2028 2737 2031
rect 2626 1988 2630 1991
rect 2598 1962 2601 1968
rect 2674 1958 2678 1961
rect 2590 1952 2593 1958
rect 2614 1952 2617 1958
rect 2686 1952 2689 1988
rect 2662 1942 2665 1948
rect 2674 1938 2678 1941
rect 2606 1922 2609 1928
rect 2574 1902 2577 1918
rect 2606 1892 2609 1918
rect 2574 1872 2577 1888
rect 2502 1848 2510 1851
rect 2562 1848 2566 1851
rect 2422 1751 2425 1758
rect 2494 1742 2497 1798
rect 2502 1792 2505 1848
rect 2542 1842 2545 1848
rect 2574 1822 2577 1868
rect 2594 1858 2598 1861
rect 2606 1852 2609 1888
rect 2614 1872 2617 1928
rect 2630 1892 2633 1938
rect 2642 1928 2646 1931
rect 2654 1922 2657 1928
rect 2646 1918 2654 1921
rect 2646 1892 2649 1918
rect 2614 1852 2617 1868
rect 2638 1862 2641 1878
rect 2678 1862 2681 1888
rect 2670 1852 2673 1858
rect 2678 1852 2681 1858
rect 2630 1842 2633 1848
rect 2694 1842 2697 1958
rect 2710 1902 2713 1928
rect 2702 1862 2705 1898
rect 2710 1852 2713 1858
rect 2586 1838 2590 1841
rect 2658 1838 2662 1841
rect 2690 1838 2694 1841
rect 2702 1822 2705 1828
rect 2542 1812 2545 1818
rect 2550 1782 2553 1788
rect 2598 1782 2601 1818
rect 2622 1802 2625 1818
rect 2670 1812 2673 1818
rect 2502 1752 2505 1778
rect 2534 1752 2537 1768
rect 2390 1692 2393 1738
rect 2390 1672 2393 1688
rect 2446 1672 2449 1728
rect 2518 1722 2521 1748
rect 2550 1742 2553 1778
rect 2646 1762 2649 1768
rect 2610 1758 2614 1761
rect 2526 1712 2529 1738
rect 2574 1732 2577 1738
rect 2590 1722 2593 1748
rect 2598 1742 2601 1748
rect 2598 1712 2601 1738
rect 2274 1658 2278 1661
rect 2330 1658 2334 1661
rect 2278 1592 2281 1598
rect 2286 1562 2289 1618
rect 2318 1542 2321 1618
rect 2350 1582 2353 1618
rect 2338 1548 2342 1551
rect 2238 1502 2241 1518
rect 2238 1472 2241 1488
rect 2246 1482 2249 1498
rect 2214 1432 2217 1448
rect 2238 1432 2241 1458
rect 2246 1452 2249 1478
rect 2246 1422 2249 1428
rect 2254 1422 2257 1538
rect 2286 1522 2289 1538
rect 2262 1462 2265 1508
rect 2270 1472 2273 1478
rect 2278 1472 2281 1488
rect 2310 1472 2313 1478
rect 2302 1462 2305 1468
rect 2286 1432 2289 1458
rect 2298 1448 2302 1451
rect 2162 1368 2166 1371
rect 2194 1368 2198 1371
rect 2174 1362 2177 1368
rect 2214 1362 2217 1368
rect 2202 1358 2206 1361
rect 2190 1342 2193 1348
rect 2150 1302 2153 1338
rect 2182 1312 2185 1338
rect 2134 1262 2137 1288
rect 2150 1252 2153 1268
rect 2174 1252 2177 1258
rect 2158 1158 2174 1161
rect 2110 1152 2113 1158
rect 2158 1152 2161 1158
rect 2182 1151 2185 1168
rect 2178 1148 2185 1151
rect 2170 1138 2174 1141
rect 2134 1112 2137 1138
rect 2146 1128 2150 1131
rect 2158 1092 2161 1108
rect 2098 1088 2102 1091
rect 2114 1048 2118 1051
rect 2126 1042 2129 1048
rect 2126 1022 2129 1038
rect 2134 992 2137 1068
rect 2142 1062 2145 1078
rect 2166 1062 2169 1098
rect 2154 1048 2158 1051
rect 2026 968 2030 971
rect 2042 968 2046 971
rect 1910 942 1913 948
rect 1974 942 1977 948
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1885 903 1888 907
rect 1902 872 1905 938
rect 1982 932 1985 938
rect 1998 932 2001 968
rect 2006 902 2009 968
rect 2054 962 2057 968
rect 2070 962 2073 988
rect 2106 978 2110 981
rect 2134 972 2137 988
rect 2070 952 2073 958
rect 2094 952 2097 968
rect 2118 952 2121 958
rect 2018 948 2022 951
rect 2038 942 2041 948
rect 1990 892 1993 898
rect 1918 872 1921 878
rect 1978 868 1982 871
rect 1882 859 1886 862
rect 1854 822 1857 858
rect 1926 822 1929 868
rect 1950 862 1953 868
rect 1958 862 1961 868
rect 1886 762 1889 768
rect 1886 752 1889 758
rect 1926 752 1929 818
rect 1842 748 1846 751
rect 1854 742 1857 748
rect 1830 738 1841 741
rect 1806 692 1809 728
rect 1806 652 1809 658
rect 1702 642 1705 648
rect 1798 642 1801 648
rect 1678 582 1681 588
rect 1610 568 1614 571
rect 1654 562 1657 568
rect 1626 558 1633 561
rect 1606 552 1609 558
rect 1618 548 1622 551
rect 1598 542 1601 548
rect 1606 542 1609 548
rect 1590 501 1593 518
rect 1590 498 1601 501
rect 1598 463 1601 498
rect 1566 392 1569 438
rect 1474 368 1478 371
rect 1510 362 1513 378
rect 1606 362 1609 408
rect 1582 358 1590 361
rect 1534 352 1537 358
rect 1582 352 1585 358
rect 1522 348 1526 351
rect 1546 348 1550 351
rect 1594 348 1598 351
rect 1614 342 1617 428
rect 1622 372 1625 508
rect 1630 492 1633 558
rect 1638 552 1641 558
rect 1682 548 1686 551
rect 1682 538 1686 541
rect 1662 492 1665 518
rect 1658 488 1662 491
rect 1670 482 1673 488
rect 1694 472 1697 478
rect 1630 462 1633 468
rect 1702 452 1705 558
rect 1718 551 1721 578
rect 1718 472 1721 528
rect 1742 512 1745 618
rect 1766 592 1769 618
rect 1782 582 1785 618
rect 1786 568 1790 571
rect 1790 522 1793 528
rect 1726 472 1729 498
rect 1734 482 1737 488
rect 1746 478 1750 481
rect 1770 478 1774 481
rect 1666 448 1670 451
rect 1662 422 1665 428
rect 1622 352 1625 368
rect 1638 362 1641 398
rect 1662 352 1665 418
rect 1650 348 1654 351
rect 1670 342 1673 388
rect 1702 382 1705 448
rect 1702 351 1705 358
rect 1718 342 1721 468
rect 1790 462 1793 468
rect 1734 402 1737 458
rect 1766 392 1769 398
rect 1790 382 1793 458
rect 1790 362 1793 368
rect 1346 338 1350 341
rect 1278 292 1281 318
rect 1294 282 1297 288
rect 1278 262 1281 268
rect 1302 262 1305 338
rect 1314 268 1318 271
rect 1138 258 1142 261
rect 1110 242 1113 258
rect 1166 252 1169 258
rect 1310 252 1313 258
rect 1102 192 1105 218
rect 1102 152 1105 168
rect 1150 152 1153 218
rect 1214 192 1217 248
rect 1318 192 1321 268
rect 1326 262 1329 338
rect 1342 332 1345 338
rect 1398 282 1401 338
rect 1438 292 1441 298
rect 1434 288 1438 291
rect 1378 278 1382 281
rect 1222 152 1225 168
rect 1034 148 1038 151
rect 1066 148 1070 151
rect 1250 148 1254 151
rect 1038 132 1041 138
rect 1030 82 1033 88
rect 1046 72 1049 148
rect 1078 142 1081 148
rect 1082 128 1086 131
rect 1062 102 1065 128
rect 1062 82 1065 98
rect 1078 72 1081 118
rect 1102 72 1105 148
rect 1118 122 1121 138
rect 1022 62 1025 68
rect 1110 62 1113 78
rect 1182 62 1185 138
rect 1222 112 1225 148
rect 1278 142 1281 158
rect 1234 138 1238 141
rect 1202 78 1206 81
rect 1214 62 1217 98
rect 1238 62 1241 118
rect 1254 82 1257 118
rect 1270 92 1273 128
rect 1318 92 1321 178
rect 1326 172 1329 258
rect 1334 192 1337 268
rect 1454 262 1457 268
rect 1374 252 1377 259
rect 1352 203 1354 207
rect 1358 203 1361 207
rect 1365 203 1368 207
rect 1458 168 1462 171
rect 1470 161 1473 308
rect 1478 262 1481 278
rect 1486 272 1489 338
rect 1542 332 1545 338
rect 1574 332 1577 338
rect 1582 332 1585 338
rect 1510 322 1513 328
rect 1518 302 1521 328
rect 1670 312 1673 338
rect 1534 292 1537 298
rect 1462 158 1473 161
rect 1494 242 1497 288
rect 1582 272 1585 288
rect 1590 282 1593 288
rect 1622 282 1625 298
rect 1518 242 1521 248
rect 1342 92 1345 158
rect 1462 152 1465 158
rect 1494 152 1497 238
rect 1534 192 1537 238
rect 1514 158 1518 161
rect 1534 152 1537 168
rect 1314 88 1318 91
rect 1350 82 1353 88
rect 1042 58 1046 61
rect 1170 58 1174 61
rect 1258 59 1262 62
rect 1326 62 1329 68
rect 1190 52 1193 58
rect 1334 52 1337 68
rect 890 48 894 51
rect 1350 42 1353 78
rect 1358 62 1361 138
rect 1374 122 1377 138
rect 1398 132 1401 148
rect 1462 102 1465 148
rect 1470 142 1473 148
rect 1534 132 1537 148
rect 1542 142 1545 268
rect 1582 262 1585 268
rect 1602 258 1606 261
rect 1566 232 1569 258
rect 1574 222 1577 258
rect 1638 252 1641 268
rect 1662 262 1665 278
rect 1686 272 1689 338
rect 1722 288 1726 291
rect 1738 278 1742 281
rect 1726 272 1729 278
rect 1742 262 1745 268
rect 1750 262 1753 308
rect 1774 302 1777 358
rect 1798 352 1801 598
rect 1814 592 1817 738
rect 1822 662 1825 668
rect 1838 592 1841 738
rect 1846 692 1849 738
rect 1958 732 1961 747
rect 1858 728 1862 731
rect 1846 672 1849 678
rect 1854 662 1857 708
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1885 703 1888 707
rect 1902 672 1905 708
rect 1958 672 1961 698
rect 1966 672 1969 688
rect 1910 622 1913 658
rect 1926 652 1929 668
rect 1942 658 1950 661
rect 1866 558 1870 561
rect 1806 542 1809 548
rect 1786 338 1790 341
rect 1798 332 1801 338
rect 1798 292 1801 318
rect 1770 278 1774 281
rect 1770 268 1774 271
rect 1782 262 1785 288
rect 1806 282 1809 528
rect 1822 502 1825 548
rect 1830 542 1833 548
rect 1838 542 1841 548
rect 1878 532 1881 578
rect 1902 552 1905 618
rect 1942 612 1945 658
rect 1954 648 1958 651
rect 1894 532 1897 538
rect 1910 532 1913 568
rect 1926 532 1929 548
rect 1934 542 1937 588
rect 1954 568 1958 571
rect 1962 558 1966 561
rect 1890 518 1897 521
rect 1822 492 1825 498
rect 1862 472 1865 518
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1885 503 1888 507
rect 1870 472 1873 478
rect 1822 463 1825 468
rect 1854 392 1857 458
rect 1862 452 1865 468
rect 1894 452 1897 518
rect 1902 472 1905 478
rect 1918 472 1921 518
rect 1926 492 1929 528
rect 1942 462 1945 468
rect 1930 458 1934 461
rect 1918 442 1921 458
rect 1950 452 1953 528
rect 1950 442 1953 448
rect 1818 358 1822 361
rect 1830 352 1833 368
rect 1818 348 1822 351
rect 1826 338 1830 341
rect 1854 322 1857 358
rect 1838 272 1841 288
rect 1482 128 1486 131
rect 1514 128 1518 131
rect 1422 82 1425 88
rect 1382 62 1385 78
rect 1486 72 1489 118
rect 1542 72 1545 138
rect 1582 132 1585 148
rect 1566 62 1569 98
rect 1574 72 1577 128
rect 1622 82 1625 88
rect 1630 62 1633 218
rect 1670 152 1673 218
rect 1658 148 1662 151
rect 1662 132 1665 138
rect 1646 92 1649 98
rect 1666 78 1670 81
rect 1678 72 1681 198
rect 1694 152 1697 208
rect 1702 152 1705 178
rect 1742 172 1745 258
rect 1790 212 1793 268
rect 1854 262 1857 318
rect 1862 292 1865 398
rect 1878 392 1881 408
rect 1878 342 1881 358
rect 1918 352 1921 428
rect 1958 412 1961 468
rect 1966 462 1969 508
rect 1974 472 1977 858
rect 1982 842 1985 858
rect 1982 782 1985 838
rect 1990 752 1993 788
rect 2038 772 2041 938
rect 2046 932 2049 938
rect 2054 911 2057 918
rect 2046 908 2057 911
rect 2046 862 2049 908
rect 2054 882 2057 898
rect 1990 702 1993 748
rect 1998 742 2001 748
rect 1986 558 1990 561
rect 1986 548 1990 551
rect 1998 522 2001 738
rect 2022 732 2025 758
rect 2034 748 2038 751
rect 2046 742 2049 748
rect 2006 722 2009 728
rect 2062 692 2065 798
rect 2070 752 2073 948
rect 2086 942 2089 948
rect 2078 932 2081 938
rect 2078 892 2081 928
rect 2086 862 2089 878
rect 2110 872 2113 938
rect 2182 922 2185 1018
rect 2174 908 2182 911
rect 2090 748 2094 751
rect 2074 738 2078 741
rect 2090 738 2094 741
rect 2006 592 2009 688
rect 2046 662 2049 668
rect 2022 652 2025 658
rect 2062 612 2065 648
rect 2038 592 2041 608
rect 2070 582 2073 678
rect 2086 672 2089 678
rect 2078 642 2081 658
rect 2102 652 2105 818
rect 2110 752 2113 868
rect 2118 862 2121 908
rect 2174 892 2177 908
rect 2190 871 2193 1278
rect 2198 1222 2201 1258
rect 2214 1151 2217 1318
rect 2210 1148 2217 1151
rect 2198 1142 2201 1148
rect 2214 1102 2217 1118
rect 2198 1062 2201 1098
rect 2222 1072 2225 1398
rect 2238 1352 2241 1358
rect 2230 1342 2233 1348
rect 2238 1331 2241 1338
rect 2230 1328 2241 1331
rect 2230 1242 2233 1328
rect 2238 1272 2241 1278
rect 2246 1262 2249 1418
rect 2258 1358 2262 1361
rect 2286 1342 2289 1348
rect 2262 1332 2265 1338
rect 2270 1261 2273 1328
rect 2262 1258 2273 1261
rect 2286 1262 2289 1308
rect 2294 1272 2297 1398
rect 2302 1392 2305 1418
rect 2310 1402 2313 1468
rect 2318 1462 2321 1508
rect 2350 1472 2353 1548
rect 2366 1472 2369 1668
rect 2494 1662 2497 1688
rect 2510 1672 2513 1678
rect 2482 1658 2486 1661
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2397 1603 2400 1607
rect 2394 1578 2398 1581
rect 2422 1562 2425 1608
rect 2454 1592 2457 1658
rect 2470 1652 2473 1658
rect 2526 1652 2529 1659
rect 2462 1582 2465 1628
rect 2462 1562 2465 1578
rect 2502 1572 2505 1578
rect 2446 1552 2449 1558
rect 2434 1548 2438 1551
rect 2406 1532 2409 1538
rect 2430 1522 2433 1538
rect 2386 1459 2390 1461
rect 2382 1458 2390 1459
rect 2322 1448 2326 1451
rect 2338 1448 2342 1451
rect 2350 1392 2353 1408
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2397 1403 2400 1407
rect 2310 1368 2329 1371
rect 2310 1351 2313 1368
rect 2326 1362 2329 1368
rect 2306 1348 2313 1351
rect 2398 1358 2406 1361
rect 2414 1361 2417 1518
rect 2430 1492 2433 1518
rect 2430 1452 2433 1458
rect 2438 1442 2441 1548
rect 2462 1492 2465 1528
rect 2486 1512 2489 1548
rect 2534 1542 2537 1708
rect 2598 1662 2601 1668
rect 2566 1562 2569 1568
rect 2486 1492 2489 1508
rect 2458 1478 2462 1481
rect 2414 1358 2422 1361
rect 2318 1352 2321 1358
rect 2398 1352 2401 1358
rect 2430 1352 2433 1418
rect 2446 1392 2449 1428
rect 2454 1392 2457 1478
rect 2494 1472 2497 1538
rect 2542 1532 2545 1538
rect 2522 1518 2526 1521
rect 2550 1512 2553 1548
rect 2574 1542 2577 1638
rect 2606 1592 2609 1718
rect 2614 1712 2617 1758
rect 2638 1752 2641 1758
rect 2678 1751 2681 1758
rect 2710 1752 2713 1788
rect 2726 1762 2729 2018
rect 2734 1942 2737 2028
rect 2734 1912 2737 1918
rect 2742 1882 2745 2028
rect 2750 1972 2753 2018
rect 2806 1992 2809 2008
rect 2822 1982 2825 2058
rect 2846 2052 2849 2118
rect 2774 1978 2801 1981
rect 2774 1972 2777 1978
rect 2790 1962 2793 1968
rect 2798 1962 2801 1978
rect 2786 1958 2790 1961
rect 2810 1958 2814 1961
rect 2774 1948 2782 1951
rect 2742 1792 2745 1878
rect 2750 1862 2753 1928
rect 2766 1922 2769 1948
rect 2774 1942 2777 1948
rect 2814 1942 2817 1948
rect 2786 1918 2790 1921
rect 2790 1882 2793 1888
rect 2766 1842 2769 1858
rect 2766 1772 2769 1778
rect 2630 1742 2633 1748
rect 2766 1742 2769 1748
rect 2774 1742 2777 1848
rect 2798 1762 2801 1928
rect 2806 1872 2809 1918
rect 2814 1872 2817 1928
rect 2822 1872 2825 1978
rect 2838 1962 2841 1968
rect 2846 1952 2849 2028
rect 2854 2002 2857 2158
rect 2974 2152 2977 2158
rect 3054 2151 3057 2158
rect 3126 2152 3129 2218
rect 3214 2212 3217 2218
rect 3222 2182 3225 2258
rect 3142 2172 3145 2178
rect 2878 2121 2881 2138
rect 2870 2118 2881 2121
rect 2870 2072 2873 2118
rect 2918 2112 2921 2148
rect 2966 2122 2969 2148
rect 3006 2142 3009 2148
rect 3126 2142 3129 2148
rect 2888 2103 2890 2107
rect 2894 2103 2897 2107
rect 2901 2103 2904 2107
rect 2958 2102 2961 2118
rect 3022 2112 3025 2128
rect 2966 2082 2969 2088
rect 2906 2078 2910 2081
rect 2922 2068 2926 2071
rect 2878 2062 2881 2068
rect 3046 2063 3049 2088
rect 3062 2072 3065 2138
rect 3078 2082 3081 2118
rect 3118 2112 3121 2118
rect 3106 2088 3110 2091
rect 2922 2058 2926 2061
rect 3102 2062 3105 2078
rect 3150 2062 3153 2178
rect 3238 2162 3241 2258
rect 3246 2162 3249 2188
rect 3234 2148 3238 2151
rect 3182 2132 3185 2148
rect 3218 2138 3222 2141
rect 3170 2118 3174 2121
rect 3166 2092 3169 2098
rect 3182 2062 3185 2108
rect 3206 2092 3209 2118
rect 3190 2072 3193 2078
rect 3214 2062 3217 2128
rect 3046 2058 3049 2059
rect 3122 2058 3126 2061
rect 2950 2052 2953 2058
rect 2930 2048 2934 2051
rect 2954 2038 2958 2041
rect 3014 1972 3017 2058
rect 3134 2052 3137 2058
rect 3082 2038 3086 2041
rect 3150 2012 3153 2058
rect 2934 1962 2937 1968
rect 2862 1942 2865 1958
rect 2918 1952 2921 1958
rect 3030 1952 3033 1968
rect 3070 1962 3073 1968
rect 3050 1958 3054 1961
rect 3090 1958 3094 1961
rect 3062 1952 3065 1958
rect 2890 1938 2894 1941
rect 2814 1862 2817 1868
rect 2822 1862 2825 1868
rect 2830 1842 2833 1858
rect 2846 1852 2849 1878
rect 2854 1842 2857 1918
rect 2862 1912 2865 1938
rect 2902 1932 2905 1938
rect 2870 1912 2873 1918
rect 2888 1903 2890 1907
rect 2894 1903 2897 1907
rect 2901 1903 2904 1907
rect 2918 1902 2921 1948
rect 2934 1942 2937 1948
rect 3078 1951 3081 1958
rect 3078 1948 3086 1951
rect 2966 1942 2969 1947
rect 2870 1872 2873 1878
rect 2950 1872 2953 1938
rect 2870 1852 2873 1868
rect 2878 1852 2881 1858
rect 2782 1742 2785 1758
rect 2814 1752 2817 1808
rect 2846 1792 2849 1828
rect 2902 1792 2905 1868
rect 2942 1842 2945 1858
rect 2966 1782 2969 1788
rect 2974 1772 2977 1898
rect 3038 1882 3041 1938
rect 3046 1931 3049 1948
rect 3102 1942 3105 1998
rect 3126 1982 3129 1988
rect 3122 1948 3126 1951
rect 3046 1928 3057 1931
rect 3046 1872 3049 1878
rect 2986 1868 2990 1871
rect 2986 1858 2990 1861
rect 2830 1762 2833 1768
rect 2858 1758 2862 1761
rect 2742 1732 2745 1738
rect 2654 1672 2657 1688
rect 2694 1682 2697 1688
rect 2754 1678 2758 1681
rect 2666 1668 2670 1671
rect 2614 1632 2617 1668
rect 2622 1662 2625 1668
rect 2654 1662 2657 1668
rect 2682 1658 2686 1661
rect 2638 1652 2641 1658
rect 2646 1652 2649 1658
rect 2626 1628 2630 1631
rect 2582 1552 2585 1578
rect 2590 1552 2593 1558
rect 2630 1551 2633 1578
rect 2558 1472 2561 1478
rect 2522 1468 2526 1471
rect 2466 1458 2470 1461
rect 2462 1352 2465 1398
rect 2494 1372 2497 1468
rect 2542 1462 2545 1468
rect 2502 1412 2505 1458
rect 2510 1452 2513 1458
rect 2550 1451 2553 1458
rect 2538 1448 2553 1451
rect 2518 1362 2521 1378
rect 2490 1358 2502 1361
rect 2478 1352 2481 1358
rect 2526 1352 2529 1358
rect 2542 1352 2545 1378
rect 2550 1352 2553 1398
rect 2574 1382 2577 1518
rect 2590 1492 2593 1548
rect 2598 1522 2601 1538
rect 2614 1532 2617 1538
rect 2594 1459 2598 1462
rect 2566 1372 2569 1378
rect 2426 1348 2430 1351
rect 2514 1348 2518 1351
rect 2334 1342 2337 1348
rect 2326 1332 2329 1338
rect 2310 1292 2313 1298
rect 2334 1292 2337 1338
rect 2342 1332 2345 1348
rect 2406 1342 2409 1348
rect 2398 1302 2401 1338
rect 2462 1332 2465 1338
rect 2406 1282 2409 1298
rect 2442 1288 2446 1291
rect 2414 1278 2422 1281
rect 2302 1262 2305 1278
rect 2382 1262 2385 1268
rect 2250 1248 2254 1251
rect 2234 1238 2238 1241
rect 2262 1212 2265 1258
rect 2270 1242 2273 1248
rect 2326 1242 2329 1248
rect 2302 1192 2305 1238
rect 2326 1192 2329 1228
rect 2342 1222 2345 1238
rect 2278 1152 2281 1168
rect 2298 1158 2302 1161
rect 2326 1152 2329 1188
rect 2234 1148 2238 1151
rect 2266 1148 2270 1151
rect 2342 1142 2345 1218
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2397 1203 2400 1207
rect 2366 1152 2369 1158
rect 2274 1138 2281 1141
rect 2246 1122 2249 1128
rect 2270 1072 2273 1098
rect 2266 1058 2270 1061
rect 2198 952 2201 978
rect 2186 868 2193 871
rect 2214 872 2217 1048
rect 2266 948 2270 951
rect 2246 942 2249 948
rect 2266 938 2270 941
rect 2230 912 2233 938
rect 2250 928 2254 931
rect 2270 882 2273 928
rect 2134 802 2137 818
rect 2110 742 2113 748
rect 2022 562 2025 568
rect 2050 558 2054 561
rect 2070 552 2073 578
rect 2094 572 2097 618
rect 2014 532 2017 538
rect 2014 522 2017 528
rect 2022 502 2025 548
rect 2030 482 2033 488
rect 1990 472 1993 478
rect 2014 472 2017 478
rect 2002 468 2006 471
rect 1982 452 1985 458
rect 1930 358 1934 361
rect 1906 348 1910 351
rect 1894 342 1897 348
rect 1934 342 1937 348
rect 1950 342 1953 378
rect 1966 342 1969 347
rect 1874 328 1878 331
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1885 303 1888 307
rect 1810 248 1814 251
rect 1830 162 1833 238
rect 1910 222 1913 338
rect 1918 262 1921 308
rect 1974 292 1977 368
rect 1998 332 2001 458
rect 2022 452 2025 458
rect 2038 402 2041 548
rect 2078 542 2081 568
rect 2046 522 2049 538
rect 2086 522 2089 548
rect 2094 542 2097 558
rect 2102 541 2105 618
rect 2110 592 2113 638
rect 2118 552 2121 768
rect 2126 732 2129 768
rect 2142 742 2145 818
rect 2158 772 2161 858
rect 2174 832 2177 848
rect 2158 751 2161 758
rect 2182 702 2185 868
rect 2222 862 2225 878
rect 2270 863 2273 868
rect 2210 858 2214 861
rect 2190 852 2193 858
rect 2210 848 2214 851
rect 2142 672 2145 678
rect 2166 662 2169 688
rect 2126 642 2129 648
rect 2138 558 2142 561
rect 2174 552 2177 698
rect 2190 682 2193 848
rect 2222 842 2225 848
rect 2238 842 2241 848
rect 2278 792 2281 1138
rect 2310 1138 2318 1141
rect 2286 952 2289 1128
rect 2310 992 2313 1138
rect 2342 1102 2345 1138
rect 2326 1072 2329 1088
rect 2334 1062 2337 1068
rect 2374 1062 2377 1188
rect 2414 1152 2417 1278
rect 2422 1262 2425 1278
rect 2446 1272 2449 1278
rect 2462 1272 2465 1318
rect 2486 1312 2489 1348
rect 2550 1342 2553 1348
rect 2558 1342 2561 1368
rect 2570 1348 2574 1351
rect 2498 1338 2502 1341
rect 2494 1282 2497 1318
rect 2454 1252 2457 1258
rect 2462 1212 2465 1268
rect 2478 1252 2481 1258
rect 2486 1252 2489 1258
rect 2422 1192 2425 1198
rect 2382 1072 2385 1098
rect 2414 1072 2417 1148
rect 2446 1142 2449 1208
rect 2454 1162 2457 1168
rect 2482 1158 2486 1161
rect 2494 1152 2497 1188
rect 2454 1142 2457 1148
rect 2446 1092 2449 1138
rect 2430 1072 2433 1078
rect 2346 1058 2350 1061
rect 2322 1038 2326 1041
rect 2334 962 2337 1058
rect 2382 1052 2385 1068
rect 2410 1058 2414 1061
rect 2462 1052 2465 1059
rect 2426 1048 2430 1051
rect 2358 1042 2361 1048
rect 2298 948 2302 951
rect 2326 942 2329 948
rect 2334 942 2337 948
rect 2358 922 2361 1038
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2397 1003 2400 1007
rect 2430 952 2433 958
rect 2470 951 2473 1148
rect 2502 1142 2505 1338
rect 2558 1332 2561 1338
rect 2530 1288 2534 1291
rect 2542 1272 2545 1328
rect 2582 1322 2585 1358
rect 2590 1342 2593 1378
rect 2598 1352 2601 1448
rect 2606 1272 2609 1468
rect 2614 1462 2617 1528
rect 2614 1362 2617 1368
rect 2614 1342 2617 1348
rect 2638 1322 2641 1648
rect 2646 1552 2649 1648
rect 2678 1562 2681 1568
rect 2710 1542 2713 1668
rect 2726 1663 2729 1668
rect 2726 1658 2729 1659
rect 2774 1642 2777 1738
rect 2774 1602 2777 1638
rect 2654 1492 2657 1508
rect 2654 1472 2657 1488
rect 2662 1352 2665 1538
rect 2710 1532 2713 1538
rect 2726 1522 2729 1547
rect 2694 1492 2697 1518
rect 2710 1492 2713 1518
rect 2742 1482 2745 1518
rect 2702 1472 2705 1478
rect 2694 1462 2697 1468
rect 2686 1422 2689 1458
rect 2670 1402 2673 1418
rect 2670 1342 2673 1348
rect 2618 1318 2622 1321
rect 2702 1282 2705 1468
rect 2726 1462 2729 1478
rect 2750 1472 2753 1588
rect 2782 1552 2785 1738
rect 2806 1732 2809 1738
rect 2794 1718 2798 1721
rect 2814 1702 2817 1748
rect 2838 1742 2841 1758
rect 2914 1748 2918 1751
rect 2974 1742 2977 1768
rect 2990 1752 2993 1758
rect 2922 1738 2926 1741
rect 2830 1732 2833 1738
rect 2888 1703 2890 1707
rect 2894 1703 2897 1707
rect 2901 1703 2904 1707
rect 2802 1668 2806 1671
rect 2814 1662 2817 1688
rect 2830 1682 2833 1688
rect 2882 1678 2886 1681
rect 2814 1642 2817 1658
rect 2822 1631 2825 1678
rect 2854 1672 2857 1678
rect 2934 1672 2937 1688
rect 2838 1662 2841 1668
rect 2878 1662 2881 1668
rect 2850 1658 2854 1661
rect 2814 1628 2825 1631
rect 2862 1632 2865 1658
rect 2902 1652 2905 1658
rect 2814 1552 2817 1628
rect 2846 1592 2849 1608
rect 2902 1592 2905 1648
rect 2878 1582 2881 1588
rect 2822 1562 2825 1568
rect 2846 1552 2849 1568
rect 2794 1538 2798 1541
rect 2790 1522 2793 1528
rect 2806 1502 2809 1548
rect 2854 1542 2857 1548
rect 2902 1532 2905 1538
rect 2826 1528 2830 1531
rect 2754 1458 2758 1461
rect 2766 1442 2769 1458
rect 2774 1452 2777 1458
rect 2806 1442 2809 1459
rect 2746 1388 2750 1391
rect 2738 1348 2742 1351
rect 2726 1332 2729 1338
rect 2734 1302 2737 1328
rect 2734 1272 2737 1298
rect 2766 1292 2769 1398
rect 2802 1348 2806 1351
rect 2522 1258 2526 1261
rect 2554 1258 2558 1261
rect 2646 1262 2649 1268
rect 2694 1262 2697 1268
rect 2718 1262 2721 1268
rect 2782 1262 2785 1318
rect 2798 1282 2801 1338
rect 2830 1272 2833 1458
rect 2862 1442 2865 1518
rect 2870 1492 2873 1528
rect 2888 1503 2890 1507
rect 2894 1503 2897 1507
rect 2901 1503 2904 1507
rect 2910 1472 2913 1598
rect 2934 1572 2937 1668
rect 2958 1642 2961 1738
rect 2982 1722 2985 1748
rect 2998 1722 3001 1858
rect 3006 1842 3009 1858
rect 3022 1852 3025 1858
rect 3006 1762 3009 1778
rect 3022 1752 3025 1838
rect 2974 1672 2977 1678
rect 2934 1552 2937 1558
rect 2942 1552 2945 1578
rect 2958 1572 2961 1578
rect 2922 1548 2926 1551
rect 2974 1542 2977 1558
rect 2982 1552 2985 1718
rect 3006 1711 3009 1748
rect 3022 1722 3025 1748
rect 3030 1742 3033 1868
rect 3054 1862 3057 1928
rect 3062 1892 3065 1908
rect 3070 1872 3073 1938
rect 3094 1892 3097 1918
rect 3102 1892 3105 1928
rect 3110 1892 3113 1928
rect 3142 1922 3145 1958
rect 3158 1952 3161 1958
rect 3150 1932 3153 1938
rect 3038 1852 3041 1858
rect 3038 1842 3041 1848
rect 3054 1802 3057 1848
rect 3070 1822 3073 1868
rect 3078 1862 3081 1868
rect 3094 1852 3097 1858
rect 3038 1762 3041 1768
rect 3070 1752 3073 1788
rect 3050 1748 3054 1751
rect 3062 1742 3065 1748
rect 2998 1708 3009 1711
rect 2990 1542 2993 1608
rect 2998 1592 3001 1708
rect 3030 1702 3033 1738
rect 3046 1732 3049 1738
rect 3006 1642 3009 1659
rect 3014 1542 3017 1598
rect 3022 1582 3025 1668
rect 3038 1662 3041 1698
rect 3070 1692 3073 1738
rect 3070 1672 3073 1678
rect 3046 1662 3049 1668
rect 3078 1662 3081 1798
rect 3102 1782 3105 1878
rect 3090 1738 3094 1741
rect 3094 1682 3097 1728
rect 3102 1692 3105 1748
rect 3110 1732 3113 1738
rect 3118 1692 3121 1858
rect 3126 1822 3129 1868
rect 3134 1862 3137 1878
rect 3158 1872 3161 1888
rect 3150 1862 3153 1868
rect 3166 1862 3169 2058
rect 3174 2042 3177 2058
rect 3222 2051 3225 2108
rect 3238 2092 3241 2118
rect 3246 2102 3249 2118
rect 3254 2092 3257 2268
rect 3270 2252 3273 2258
rect 3262 2192 3265 2248
rect 3242 2058 3246 2061
rect 3218 2048 3225 2051
rect 3190 2028 3198 2031
rect 3190 1962 3193 2028
rect 3178 1958 3182 1961
rect 3198 1942 3201 2018
rect 3198 1932 3201 1938
rect 3182 1862 3185 1898
rect 3206 1892 3209 2048
rect 3238 1992 3241 2018
rect 3254 1992 3257 2048
rect 3262 1972 3265 2118
rect 3270 2092 3273 2218
rect 3294 2192 3297 2318
rect 3310 2292 3313 2318
rect 3350 2312 3353 2338
rect 3314 2268 3318 2271
rect 3302 2212 3305 2248
rect 3326 2242 3329 2268
rect 3334 2192 3337 2288
rect 3374 2192 3377 2308
rect 3382 2292 3385 2338
rect 3398 2302 3401 2328
rect 3406 2302 3409 2358
rect 3414 2292 3417 2378
rect 3422 2362 3425 2388
rect 3422 2342 3425 2358
rect 3438 2352 3441 2398
rect 3462 2352 3465 2448
rect 3478 2402 3481 2458
rect 3498 2448 3502 2451
rect 3510 2442 3513 2458
rect 3518 2422 3521 2458
rect 3486 2368 3494 2371
rect 3486 2352 3489 2368
rect 3510 2352 3513 2368
rect 3518 2352 3521 2418
rect 3526 2402 3529 2458
rect 3558 2451 3561 2518
rect 3606 2472 3609 2478
rect 3554 2448 3561 2451
rect 3434 2348 3438 2351
rect 3446 2342 3449 2348
rect 3430 2312 3433 2338
rect 3462 2332 3465 2348
rect 3518 2342 3521 2348
rect 3526 2342 3529 2368
rect 3542 2352 3545 2368
rect 3478 2322 3481 2338
rect 3494 2322 3497 2338
rect 3550 2332 3553 2348
rect 3522 2318 3526 2321
rect 3446 2282 3449 2308
rect 3458 2288 3462 2291
rect 3490 2288 3494 2291
rect 3478 2282 3481 2288
rect 3446 2272 3449 2278
rect 3426 2266 3430 2269
rect 3466 2268 3478 2271
rect 3486 2268 3494 2271
rect 3382 2242 3385 2248
rect 3400 2203 3402 2207
rect 3406 2203 3409 2207
rect 3413 2203 3416 2207
rect 3438 2202 3441 2268
rect 3502 2262 3505 2308
rect 3522 2268 3526 2271
rect 3510 2262 3513 2268
rect 3470 2222 3473 2258
rect 3534 2252 3537 2278
rect 3558 2272 3561 2438
rect 3574 2421 3577 2468
rect 3582 2452 3585 2468
rect 3582 2432 3585 2448
rect 3598 2442 3601 2458
rect 3614 2452 3617 2508
rect 3626 2458 3630 2461
rect 3646 2452 3649 2538
rect 3654 2482 3657 2498
rect 3574 2418 3585 2421
rect 3582 2412 3585 2418
rect 3574 2352 3577 2358
rect 3590 2352 3593 2378
rect 3550 2252 3553 2268
rect 3566 2262 3569 2288
rect 3598 2282 3601 2288
rect 3594 2268 3598 2271
rect 3582 2262 3585 2268
rect 3526 2212 3529 2248
rect 3434 2178 3438 2181
rect 3278 2152 3281 2168
rect 3306 2158 3310 2161
rect 3358 2152 3361 2158
rect 3322 2148 3326 2151
rect 3294 2142 3297 2148
rect 3350 2142 3353 2148
rect 3282 2138 3286 2141
rect 3346 2088 3350 2091
rect 3286 2062 3289 2088
rect 3326 2062 3329 2068
rect 3278 1992 3281 2008
rect 3222 1932 3225 1958
rect 3274 1948 3281 1951
rect 3230 1912 3233 1948
rect 3266 1938 3270 1941
rect 3278 1912 3281 1948
rect 3286 1932 3289 2058
rect 3294 2052 3297 2058
rect 3294 1952 3297 1998
rect 3318 1982 3321 2058
rect 3334 2022 3337 2078
rect 3358 2072 3361 2098
rect 3366 2062 3369 2088
rect 3346 2058 3350 2061
rect 3382 2052 3385 2158
rect 3390 2152 3393 2168
rect 3470 2152 3473 2168
rect 3534 2152 3537 2168
rect 3542 2152 3545 2218
rect 3494 2132 3497 2138
rect 3398 2092 3401 2108
rect 3454 2102 3457 2118
rect 3390 2082 3393 2088
rect 3518 2082 3521 2118
rect 3550 2072 3553 2238
rect 3558 2192 3561 2248
rect 3582 2222 3585 2248
rect 3570 2218 3574 2221
rect 3598 2152 3601 2168
rect 3466 2068 3470 2071
rect 3406 2062 3409 2068
rect 3414 2062 3417 2068
rect 3478 2062 3481 2068
rect 3450 2058 3454 2061
rect 3554 2058 3558 2061
rect 3370 2038 3374 2041
rect 3400 2003 3402 2007
rect 3406 2003 3409 2007
rect 3413 2003 3416 2007
rect 3438 1982 3441 2058
rect 3430 1962 3433 1968
rect 3294 1902 3297 1948
rect 3442 1948 3446 1951
rect 3366 1942 3369 1947
rect 3418 1938 3422 1941
rect 3450 1938 3454 1941
rect 3462 1932 3465 1938
rect 3306 1918 3310 1921
rect 3290 1888 3294 1891
rect 3262 1882 3265 1888
rect 3366 1882 3369 1928
rect 3398 1922 3401 1928
rect 3470 1922 3473 2058
rect 3502 1952 3505 2028
rect 3510 1962 3513 2048
rect 3494 1922 3497 1948
rect 3414 1882 3417 1918
rect 3454 1892 3457 1908
rect 3246 1878 3254 1881
rect 3190 1862 3193 1868
rect 3238 1862 3241 1868
rect 3226 1858 3230 1861
rect 3246 1861 3249 1878
rect 3366 1872 3369 1878
rect 3258 1868 3262 1871
rect 3326 1862 3329 1868
rect 3246 1858 3262 1861
rect 3274 1858 3278 1861
rect 3126 1792 3129 1808
rect 3142 1762 3145 1818
rect 3142 1752 3145 1758
rect 3166 1752 3169 1858
rect 3214 1852 3217 1858
rect 3178 1848 3182 1851
rect 3182 1822 3185 1848
rect 3238 1802 3241 1858
rect 3186 1758 3190 1761
rect 3126 1732 3129 1748
rect 3134 1742 3137 1748
rect 3170 1738 3174 1741
rect 3122 1678 3126 1681
rect 3142 1672 3145 1678
rect 3150 1672 3153 1688
rect 3090 1668 3094 1671
rect 3158 1662 3161 1698
rect 3198 1692 3201 1788
rect 3238 1742 3241 1748
rect 3206 1682 3209 1718
rect 3222 1672 3225 1688
rect 3210 1668 3214 1671
rect 3082 1658 3086 1661
rect 3138 1658 3142 1661
rect 3038 1652 3041 1658
rect 3054 1642 3057 1658
rect 3174 1652 3177 1668
rect 3106 1648 3110 1651
rect 3118 1592 3121 1648
rect 3046 1552 3049 1568
rect 3070 1562 3073 1568
rect 2994 1528 2998 1531
rect 2934 1522 2937 1528
rect 2934 1492 2937 1508
rect 2914 1468 2921 1471
rect 2882 1458 2886 1461
rect 2894 1452 2897 1458
rect 2878 1432 2881 1438
rect 2878 1412 2881 1428
rect 2870 1312 2873 1347
rect 2878 1291 2881 1408
rect 2898 1328 2902 1331
rect 2918 1322 2921 1468
rect 2926 1422 2929 1458
rect 2942 1452 2945 1478
rect 2950 1462 2953 1468
rect 2888 1303 2890 1307
rect 2894 1303 2897 1307
rect 2901 1303 2904 1307
rect 2878 1288 2889 1291
rect 2794 1268 2798 1271
rect 2858 1268 2862 1271
rect 2870 1262 2873 1268
rect 2886 1262 2889 1288
rect 2918 1271 2921 1318
rect 2914 1268 2921 1271
rect 2534 1181 2537 1248
rect 2542 1192 2545 1258
rect 2566 1252 2569 1258
rect 2598 1252 2601 1259
rect 2738 1258 2742 1261
rect 2770 1258 2774 1261
rect 2914 1258 2918 1261
rect 2714 1248 2718 1251
rect 2566 1192 2569 1218
rect 2534 1178 2542 1181
rect 2514 1148 2518 1151
rect 2534 1142 2537 1158
rect 2550 1142 2553 1168
rect 2566 1152 2569 1158
rect 2582 1152 2585 1158
rect 2590 1152 2593 1178
rect 2654 1142 2657 1148
rect 2610 1138 2614 1141
rect 2502 1102 2505 1138
rect 2518 1082 2521 1118
rect 2526 1092 2529 1128
rect 2494 1062 2497 1068
rect 2466 948 2473 951
rect 2350 912 2353 918
rect 2302 862 2305 908
rect 2350 872 2353 908
rect 2330 838 2334 841
rect 2218 768 2222 771
rect 2278 752 2281 758
rect 2286 752 2289 838
rect 2342 832 2345 868
rect 2234 748 2238 751
rect 2258 748 2262 751
rect 2246 742 2249 748
rect 2294 742 2297 798
rect 2302 762 2305 768
rect 2342 762 2345 828
rect 2358 792 2361 898
rect 2374 892 2377 948
rect 2462 942 2465 948
rect 2442 938 2446 941
rect 2406 932 2409 938
rect 2430 872 2433 878
rect 2378 858 2382 861
rect 2402 858 2406 861
rect 2390 842 2393 848
rect 2414 812 2417 868
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2397 803 2400 807
rect 2322 758 2326 761
rect 2306 748 2310 751
rect 2330 748 2334 751
rect 2258 738 2262 741
rect 2282 738 2286 741
rect 2234 688 2238 691
rect 2226 668 2230 671
rect 2190 641 2193 668
rect 2218 658 2222 661
rect 2206 642 2209 648
rect 2238 642 2241 648
rect 2246 642 2249 728
rect 2262 672 2265 698
rect 2270 692 2273 738
rect 2254 662 2257 668
rect 2270 652 2273 658
rect 2190 638 2201 641
rect 2198 572 2201 638
rect 2222 632 2225 638
rect 2182 562 2185 568
rect 2278 562 2281 678
rect 2294 672 2297 738
rect 2318 728 2326 731
rect 2318 682 2321 728
rect 2342 662 2345 758
rect 2398 752 2401 778
rect 2422 752 2425 818
rect 2446 792 2449 868
rect 2454 862 2457 938
rect 2478 932 2481 948
rect 2494 942 2497 1058
rect 2430 752 2433 768
rect 2446 752 2449 758
rect 2418 748 2422 751
rect 2362 738 2366 741
rect 2358 662 2361 718
rect 2366 682 2369 738
rect 2238 552 2241 558
rect 2278 552 2281 558
rect 2178 548 2185 551
rect 2102 538 2110 541
rect 2154 538 2158 541
rect 2170 538 2174 541
rect 2102 532 2105 538
rect 2110 522 2113 528
rect 2038 382 2041 398
rect 2038 342 2041 348
rect 2046 332 2049 518
rect 2054 482 2057 518
rect 2074 478 2078 481
rect 2074 468 2078 471
rect 2054 462 2057 468
rect 2086 452 2089 458
rect 2070 442 2073 448
rect 2070 352 2073 418
rect 2086 362 2089 368
rect 2094 351 2097 468
rect 2102 462 2105 508
rect 2110 472 2113 478
rect 2102 422 2105 458
rect 2118 432 2121 458
rect 2134 452 2137 458
rect 2142 452 2145 458
rect 2094 348 2105 351
rect 2058 338 2062 341
rect 2094 332 2097 338
rect 2034 328 2038 331
rect 2058 328 2062 331
rect 2026 318 2030 321
rect 2090 318 2094 321
rect 2102 302 2105 348
rect 2114 348 2118 351
rect 1998 282 2001 298
rect 2110 272 2113 348
rect 2134 342 2137 348
rect 2126 312 2129 318
rect 2126 292 2129 298
rect 2142 292 2145 428
rect 2150 352 2153 498
rect 2166 492 2169 508
rect 2182 502 2185 548
rect 2282 538 2286 541
rect 2262 522 2265 538
rect 2178 488 2182 491
rect 2262 472 2265 518
rect 2294 512 2297 658
rect 2342 652 2345 658
rect 2302 562 2305 568
rect 2366 552 2369 668
rect 2382 622 2385 748
rect 2402 718 2406 721
rect 2438 702 2441 738
rect 2454 692 2457 848
rect 2438 672 2441 678
rect 2418 668 2422 671
rect 2450 668 2454 671
rect 2410 648 2414 651
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2397 603 2400 607
rect 2406 592 2409 638
rect 2430 602 2433 658
rect 2454 592 2457 658
rect 2438 562 2441 568
rect 2302 542 2305 548
rect 2334 542 2337 547
rect 2366 542 2369 548
rect 2318 522 2321 538
rect 2278 472 2281 498
rect 2162 458 2166 461
rect 2174 412 2177 468
rect 2242 459 2246 462
rect 2150 302 2153 348
rect 2158 332 2161 338
rect 2166 292 2169 408
rect 2206 392 2209 408
rect 2174 352 2177 368
rect 2182 352 2185 358
rect 2214 352 2217 368
rect 2246 362 2249 368
rect 2262 362 2265 468
rect 2294 462 2297 468
rect 2278 392 2281 448
rect 2286 442 2289 458
rect 2310 452 2313 488
rect 2310 352 2313 358
rect 2266 338 2270 341
rect 2190 322 2193 338
rect 2210 328 2214 331
rect 2230 322 2233 338
rect 2158 282 2161 288
rect 2162 278 2166 281
rect 1962 268 1966 271
rect 2018 268 2022 271
rect 1830 152 1833 158
rect 1886 152 1889 208
rect 1690 148 1694 151
rect 1770 147 1774 150
rect 1810 148 1814 151
rect 1850 148 1854 151
rect 1822 142 1825 148
rect 1894 142 1897 168
rect 1910 142 1913 148
rect 1926 142 1929 268
rect 1982 262 1985 268
rect 2010 258 2014 261
rect 1974 192 1977 238
rect 1982 202 1985 258
rect 2030 212 2033 258
rect 2062 252 2065 259
rect 2062 192 2065 218
rect 2002 188 2006 191
rect 1942 151 1945 158
rect 1974 152 1977 168
rect 2038 152 2041 158
rect 2018 148 2022 151
rect 2030 142 2033 148
rect 1790 132 1793 138
rect 1686 92 1689 118
rect 1710 112 1713 118
rect 1790 72 1793 128
rect 1806 112 1809 128
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1885 103 1888 107
rect 1866 88 1870 91
rect 1642 68 1646 71
rect 1678 62 1681 68
rect 1750 63 1753 68
rect 1410 58 1414 61
rect 1814 62 1817 68
rect 1894 62 1897 138
rect 1926 132 1929 138
rect 1902 128 1910 131
rect 1902 92 1905 128
rect 1910 82 1913 88
rect 1942 82 1945 128
rect 1950 62 1953 118
rect 1974 82 1977 128
rect 2014 112 2017 128
rect 2006 92 2009 98
rect 2046 72 2049 168
rect 2062 152 2065 188
rect 2094 172 2097 258
rect 2110 212 2113 268
rect 2182 262 2185 298
rect 2230 282 2233 318
rect 2246 292 2249 328
rect 2254 282 2257 338
rect 2270 292 2273 328
rect 2126 258 2134 261
rect 2102 162 2105 208
rect 2102 152 2105 158
rect 2126 152 2129 258
rect 2174 252 2177 258
rect 2190 152 2193 268
rect 2222 262 2225 268
rect 2230 262 2233 278
rect 2214 252 2217 258
rect 2198 152 2201 168
rect 2238 152 2241 268
rect 2278 262 2281 278
rect 2286 262 2289 348
rect 2302 272 2305 278
rect 2258 258 2262 261
rect 2246 192 2249 248
rect 2270 152 2273 178
rect 2310 162 2313 338
rect 2318 332 2321 508
rect 2330 468 2334 471
rect 2358 462 2361 528
rect 2366 472 2369 478
rect 2390 472 2393 558
rect 2446 552 2449 588
rect 2418 468 2422 471
rect 2330 458 2334 461
rect 2338 448 2342 451
rect 2342 351 2345 368
rect 2358 362 2361 418
rect 2374 352 2377 468
rect 2430 462 2433 528
rect 2418 458 2422 461
rect 2398 442 2401 458
rect 2418 448 2422 451
rect 2430 442 2433 448
rect 2402 438 2409 441
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2397 403 2400 407
rect 2386 358 2390 361
rect 2398 352 2401 368
rect 2406 352 2409 438
rect 2430 352 2433 358
rect 2318 292 2321 328
rect 2310 152 2313 158
rect 2090 148 2094 151
rect 2122 148 2126 151
rect 2258 148 2262 151
rect 2282 148 2286 151
rect 2134 142 2137 148
rect 2078 132 2081 138
rect 2054 82 2057 118
rect 2062 62 2065 108
rect 2094 92 2097 138
rect 2106 88 2110 91
rect 2118 62 2121 68
rect 2142 62 2145 68
rect 2150 62 2153 98
rect 2190 82 2193 138
rect 2318 132 2321 258
rect 2334 152 2337 208
rect 2366 182 2369 268
rect 2374 152 2377 348
rect 2410 338 2414 341
rect 2382 263 2385 318
rect 2422 312 2425 348
rect 2438 312 2441 548
rect 2446 532 2449 538
rect 2462 492 2465 838
rect 2470 762 2473 878
rect 2494 842 2497 938
rect 2510 892 2513 948
rect 2518 942 2521 948
rect 2526 892 2529 1078
rect 2534 1062 2537 1068
rect 2550 1032 2553 1138
rect 2558 1082 2561 1138
rect 2646 1082 2649 1128
rect 2658 1088 2662 1091
rect 2574 1072 2577 1078
rect 2658 1068 2662 1071
rect 2670 1062 2673 1188
rect 2722 1168 2726 1171
rect 2730 1148 2734 1151
rect 2738 1138 2742 1141
rect 2678 1068 2694 1071
rect 2678 1062 2681 1068
rect 2710 1062 2713 1078
rect 2730 1068 2734 1071
rect 2718 1062 2721 1068
rect 2602 1058 2606 1061
rect 2558 1052 2561 1058
rect 2670 1042 2673 1058
rect 2686 1052 2689 1058
rect 2734 1042 2737 1058
rect 2750 1052 2753 1068
rect 2758 1041 2761 1258
rect 2766 1152 2769 1168
rect 2782 1162 2785 1208
rect 2774 1102 2777 1148
rect 2790 1132 2793 1138
rect 2798 1092 2801 1148
rect 2806 1142 2809 1148
rect 2830 1142 2833 1168
rect 2846 1162 2849 1178
rect 2854 1152 2857 1258
rect 2870 1192 2873 1258
rect 2926 1252 2929 1418
rect 2958 1402 2961 1458
rect 2974 1372 2977 1518
rect 3014 1512 3017 1538
rect 3034 1528 3038 1531
rect 3046 1522 3049 1538
rect 3070 1532 3073 1558
rect 3078 1512 3081 1578
rect 3110 1572 3113 1578
rect 3090 1548 3094 1551
rect 3098 1538 3102 1541
rect 3086 1532 3089 1538
rect 2990 1472 2993 1498
rect 2998 1472 3001 1478
rect 2982 1392 2985 1458
rect 2998 1442 3001 1458
rect 3014 1452 3017 1478
rect 3030 1392 3033 1498
rect 3078 1462 3081 1508
rect 3110 1492 3113 1498
rect 3118 1462 3121 1468
rect 3126 1462 3129 1548
rect 3150 1542 3153 1548
rect 3190 1542 3193 1648
rect 3198 1642 3201 1648
rect 3230 1642 3233 1658
rect 3254 1652 3257 1738
rect 3270 1672 3273 1678
rect 3270 1652 3273 1658
rect 3214 1592 3217 1638
rect 3230 1592 3233 1628
rect 3222 1562 3225 1568
rect 3238 1552 3241 1568
rect 3278 1562 3281 1858
rect 3298 1748 3302 1751
rect 3318 1742 3321 1758
rect 3326 1752 3329 1758
rect 3374 1751 3377 1758
rect 3382 1752 3385 1858
rect 3390 1832 3393 1868
rect 3438 1842 3441 1858
rect 3486 1852 3489 1858
rect 3502 1852 3505 1948
rect 3518 1882 3521 2038
rect 3526 1992 3529 2008
rect 3542 1952 3545 1978
rect 3582 1972 3585 2118
rect 3606 2092 3609 2408
rect 3614 2372 3617 2448
rect 3630 2362 3633 2418
rect 3646 2352 3649 2368
rect 3634 2348 3638 2351
rect 3614 2292 3617 2348
rect 3622 2322 3625 2348
rect 3638 2312 3641 2338
rect 3654 2332 3657 2468
rect 3678 2462 3681 2528
rect 3686 2472 3689 2518
rect 3694 2472 3697 2798
rect 3702 2692 3705 2958
rect 3758 2952 3761 2968
rect 3766 2952 3769 2958
rect 3798 2952 3801 2958
rect 3746 2948 3750 2951
rect 3718 2942 3721 2948
rect 3734 2882 3737 2888
rect 3782 2882 3785 2918
rect 3750 2862 3753 2868
rect 3782 2862 3785 2868
rect 3798 2862 3801 2948
rect 3806 2892 3809 2978
rect 3854 2942 3857 3138
rect 3870 3072 3873 3158
rect 3902 3152 3905 3248
rect 3910 3152 3913 3178
rect 3890 3138 3902 3141
rect 3878 3128 3886 3131
rect 3878 3022 3881 3128
rect 3890 3078 3902 3081
rect 3890 3068 3894 3071
rect 3902 3062 3905 3068
rect 3898 3048 3902 3051
rect 3886 3042 3889 3048
rect 3910 3011 3913 3118
rect 3920 3103 3922 3107
rect 3926 3103 3929 3107
rect 3933 3103 3936 3107
rect 3934 3082 3937 3088
rect 3918 3011 3921 3058
rect 3910 3008 3921 3011
rect 3862 2922 3865 2948
rect 3838 2892 3841 2908
rect 3830 2862 3833 2868
rect 3854 2862 3857 2888
rect 3850 2858 3854 2861
rect 3782 2792 3785 2838
rect 3790 2822 3793 2858
rect 3798 2762 3801 2858
rect 3806 2762 3809 2818
rect 3710 2751 3713 2758
rect 3766 2752 3769 2758
rect 3798 2752 3801 2758
rect 3806 2732 3809 2738
rect 3750 2722 3753 2728
rect 3718 2662 3721 2688
rect 3730 2668 3734 2671
rect 3702 2612 3705 2618
rect 3742 2552 3745 2708
rect 3754 2668 3758 2671
rect 3790 2662 3793 2668
rect 3814 2662 3817 2668
rect 3822 2662 3825 2698
rect 3830 2672 3833 2678
rect 3846 2662 3849 2848
rect 3870 2752 3873 2868
rect 3902 2862 3905 2878
rect 3910 2872 3913 3008
rect 3926 2992 3929 3068
rect 3926 2962 3929 2968
rect 3934 2932 3937 3048
rect 3942 2952 3945 3258
rect 4022 3242 4025 3248
rect 3962 3158 3966 3161
rect 3982 3082 3985 3098
rect 3990 3092 3993 3238
rect 4030 3202 4033 3338
rect 4038 3332 4041 3348
rect 4062 3342 4065 3378
rect 4078 3362 4081 3418
rect 4094 3372 4097 3418
rect 4110 3382 4113 3438
rect 4126 3392 4129 3448
rect 4078 3342 4081 3358
rect 4094 3352 4097 3358
rect 4046 3272 4049 3328
rect 4094 3302 4097 3338
rect 4102 3322 4105 3348
rect 4110 3342 4113 3368
rect 4134 3352 4137 3608
rect 4190 3582 4193 3618
rect 4158 3552 4161 3558
rect 4182 3552 4185 3568
rect 4222 3562 4225 3668
rect 4230 3662 4233 3698
rect 4254 3662 4257 3818
rect 4270 3762 4273 3858
rect 4278 3832 4281 3918
rect 4302 3882 4305 3918
rect 4302 3862 4305 3878
rect 4310 3862 4313 3878
rect 4318 3872 4321 3918
rect 4334 3882 4337 3898
rect 4342 3872 4345 3988
rect 4374 3962 4377 3968
rect 4350 3942 4353 3958
rect 4346 3858 4350 3861
rect 4294 3852 4297 3858
rect 4310 3851 4313 3858
rect 4302 3848 4313 3851
rect 4278 3751 4281 3818
rect 4274 3748 4281 3751
rect 4262 3672 4265 3678
rect 4302 3672 4305 3848
rect 4318 3792 4321 3848
rect 4334 3761 4337 3818
rect 4330 3758 4337 3761
rect 4342 3752 4345 3798
rect 4334 3732 4337 3738
rect 4310 3722 4313 3728
rect 4326 3722 4329 3728
rect 4318 3682 4321 3718
rect 4330 3668 4334 3671
rect 4350 3671 4353 3818
rect 4358 3802 4361 3948
rect 4446 3942 4449 3947
rect 4462 3942 4465 4068
rect 4562 4058 4566 4061
rect 4486 4052 4489 4058
rect 4518 3972 4521 4018
rect 4490 3958 4494 3961
rect 4506 3948 4510 3951
rect 4382 3861 4385 3918
rect 4446 3912 4449 3928
rect 4398 3892 4401 3898
rect 4390 3862 4393 3868
rect 4414 3862 4417 3878
rect 4422 3872 4425 3878
rect 4430 3862 4433 3878
rect 4382 3858 4390 3861
rect 4370 3848 4374 3851
rect 4358 3752 4361 3758
rect 4374 3752 4377 3828
rect 4374 3742 4377 3748
rect 4358 3722 4361 3728
rect 4366 3692 4369 3738
rect 4382 3692 4385 3848
rect 4398 3772 4401 3848
rect 4424 3803 4426 3807
rect 4430 3803 4433 3807
rect 4437 3803 4440 3807
rect 4406 3762 4409 3768
rect 4390 3732 4393 3758
rect 4446 3752 4449 3908
rect 4478 3892 4481 3948
rect 4518 3942 4521 3948
rect 4550 3932 4553 4058
rect 4494 3882 4497 3918
rect 4502 3872 4505 3898
rect 4486 3862 4489 3868
rect 4510 3862 4513 3878
rect 4534 3872 4537 3898
rect 4542 3862 4545 3908
rect 4558 3891 4561 3948
rect 4566 3942 4569 4018
rect 4646 3952 4649 4168
rect 4654 4142 4657 4158
rect 4678 4152 4681 4698
rect 4686 4682 4689 4688
rect 4694 4652 4697 4718
rect 4710 4702 4713 4748
rect 4750 4742 4753 4778
rect 4726 4722 4729 4728
rect 4722 4688 4726 4691
rect 4710 4662 4713 4668
rect 4702 4652 4705 4658
rect 4718 4592 4721 4658
rect 4726 4571 4729 4618
rect 4718 4568 4729 4571
rect 4690 4558 4694 4561
rect 4694 4552 4697 4558
rect 4718 4552 4721 4568
rect 4726 4552 4729 4558
rect 4734 4552 4737 4558
rect 4742 4552 4745 4718
rect 4758 4712 4761 4748
rect 4766 4741 4769 5059
rect 4782 4992 4785 5028
rect 4806 4972 4809 5018
rect 4806 4952 4809 4958
rect 4778 4948 4782 4951
rect 4798 4942 4801 4948
rect 4790 4862 4793 4868
rect 4798 4782 4801 4938
rect 4806 4872 4809 4948
rect 4822 4942 4825 4948
rect 4838 4912 4841 4947
rect 4862 4942 4865 5068
rect 4902 5052 4905 5058
rect 4926 5052 4929 5058
rect 4982 5052 4985 5068
rect 4994 5058 4998 5061
rect 5050 5058 5054 5061
rect 4962 5018 4966 5021
rect 4870 4952 4873 4958
rect 4914 4948 4918 4951
rect 4870 4882 4873 4948
rect 4974 4942 4977 4948
rect 4970 4938 4974 4941
rect 4898 4918 4902 4921
rect 4936 4903 4938 4907
rect 4942 4903 4945 4907
rect 4949 4903 4952 4907
rect 4970 4888 4974 4891
rect 4878 4862 4881 4878
rect 4974 4872 4977 4878
rect 4806 4752 4809 4758
rect 4766 4738 4774 4741
rect 4770 4718 4774 4721
rect 4854 4682 4857 4688
rect 4894 4681 4897 4848
rect 4910 4742 4913 4748
rect 4918 4722 4921 4748
rect 4974 4732 4977 4848
rect 4990 4822 4993 5018
rect 5006 4972 5009 5038
rect 5014 4942 5017 5048
rect 5022 4952 5025 5058
rect 5014 4932 5017 4938
rect 5006 4922 5009 4928
rect 5022 4922 5025 4948
rect 4998 4812 5001 4918
rect 5030 4892 5033 5038
rect 5038 4952 5041 4958
rect 5006 4862 5009 4868
rect 5014 4862 5017 4868
rect 5022 4862 5025 4888
rect 5006 4782 5009 4858
rect 5014 4812 5017 4858
rect 5030 4851 5033 4868
rect 5022 4848 5033 4851
rect 4998 4752 5001 4768
rect 5006 4762 5009 4768
rect 5022 4752 5025 4848
rect 4970 4728 4974 4731
rect 4936 4703 4938 4707
rect 4942 4703 4945 4707
rect 4949 4703 4952 4707
rect 4906 4688 4910 4691
rect 4894 4678 4905 4681
rect 4758 4552 4761 4668
rect 4894 4662 4897 4668
rect 4902 4662 4905 4678
rect 4966 4672 4969 4718
rect 4866 4658 4870 4661
rect 4686 4512 4689 4548
rect 4758 4542 4761 4548
rect 4698 4538 4702 4541
rect 4722 4538 4726 4541
rect 4686 4472 4689 4498
rect 4694 4342 4697 4488
rect 4702 4392 4705 4528
rect 4718 4502 4721 4538
rect 4750 4528 4758 4531
rect 4750 4522 4753 4528
rect 4766 4521 4769 4658
rect 4774 4552 4777 4658
rect 4782 4652 4785 4658
rect 4846 4622 4849 4658
rect 4886 4652 4889 4658
rect 4902 4642 4905 4658
rect 4806 4552 4809 4578
rect 4814 4552 4817 4608
rect 4830 4552 4833 4618
rect 4974 4602 4977 4728
rect 4990 4722 4993 4728
rect 4982 4682 4985 4718
rect 4990 4682 4993 4718
rect 4998 4702 5001 4738
rect 4982 4652 4985 4658
rect 4774 4542 4777 4548
rect 4794 4538 4798 4541
rect 4758 4518 4769 4521
rect 4726 4482 4729 4518
rect 4742 4462 4745 4508
rect 4758 4472 4761 4518
rect 4790 4512 4793 4518
rect 4790 4472 4793 4498
rect 4822 4492 4825 4548
rect 4838 4541 4841 4558
rect 4854 4552 4857 4568
rect 4974 4562 4977 4568
rect 4994 4558 4998 4561
rect 4830 4538 4841 4541
rect 4846 4542 4849 4548
rect 4754 4468 4758 4471
rect 4802 4458 4806 4461
rect 4814 4452 4817 4478
rect 4822 4462 4825 4488
rect 4830 4482 4833 4538
rect 4854 4492 4857 4548
rect 4862 4532 4865 4538
rect 4878 4522 4881 4548
rect 4910 4542 4913 4547
rect 4862 4472 4865 4518
rect 4858 4458 4862 4461
rect 4834 4448 4838 4451
rect 4726 4392 4729 4448
rect 4798 4392 4801 4418
rect 4846 4402 4849 4458
rect 4870 4412 4873 4518
rect 4894 4472 4897 4538
rect 4936 4503 4938 4507
rect 4942 4503 4945 4507
rect 4949 4503 4952 4507
rect 4902 4462 4905 4488
rect 4930 4468 4934 4471
rect 4942 4462 4945 4478
rect 4702 4352 4705 4388
rect 4766 4362 4769 4388
rect 4686 4262 4689 4318
rect 4702 4262 4705 4348
rect 4710 4342 4713 4348
rect 4750 4342 4753 4348
rect 4730 4338 4734 4341
rect 4758 4282 4761 4338
rect 4766 4292 4769 4348
rect 4774 4322 4777 4328
rect 4702 4152 4705 4258
rect 4714 4158 4718 4161
rect 4678 4142 4681 4148
rect 4698 4138 4702 4141
rect 4654 4102 4657 4138
rect 4710 4132 4713 4148
rect 4726 4122 4729 4268
rect 4742 4262 4745 4278
rect 4782 4262 4785 4368
rect 4878 4362 4881 4418
rect 4810 4348 4814 4351
rect 4790 4282 4793 4318
rect 4806 4292 4809 4338
rect 4830 4272 4833 4348
rect 4854 4342 4857 4358
rect 4882 4348 4886 4351
rect 4870 4312 4873 4348
rect 4866 4288 4870 4291
rect 4790 4262 4793 4268
rect 4894 4262 4897 4358
rect 4902 4352 4905 4458
rect 4958 4442 4961 4478
rect 4974 4472 4977 4518
rect 4990 4501 4993 4518
rect 5006 4512 5009 4718
rect 5022 4702 5025 4748
rect 5030 4742 5033 4758
rect 5038 4751 5041 4918
rect 5046 4902 5049 5018
rect 5078 4942 5081 4948
rect 5046 4852 5049 4878
rect 5054 4842 5057 4878
rect 5078 4872 5081 4928
rect 5086 4892 5089 4958
rect 5066 4868 5070 4871
rect 5082 4858 5086 4861
rect 5094 4852 5097 5058
rect 5046 4772 5049 4818
rect 5054 4802 5057 4818
rect 5038 4748 5046 4751
rect 5042 4718 5046 4721
rect 5022 4652 5025 4678
rect 5038 4662 5041 4698
rect 5070 4692 5073 4738
rect 5046 4672 5049 4678
rect 5062 4662 5065 4668
rect 5078 4661 5081 4838
rect 5086 4702 5089 4818
rect 5102 4772 5105 4948
rect 5110 4942 5113 5058
rect 5146 5018 5150 5021
rect 5150 4932 5153 4938
rect 5166 4892 5169 5018
rect 5174 4922 5177 4948
rect 5166 4872 5169 4878
rect 5134 4752 5137 4778
rect 5086 4672 5089 4678
rect 5102 4672 5105 4747
rect 5118 4732 5121 4738
rect 5134 4662 5137 4738
rect 5142 4712 5145 4858
rect 5150 4662 5153 4808
rect 5158 4742 5161 4748
rect 5166 4742 5169 4748
rect 5182 4722 5185 4868
rect 5222 4842 5225 5068
rect 5242 5058 5246 5061
rect 5302 5042 5305 5048
rect 5230 4912 5233 4918
rect 5238 4862 5241 5018
rect 5246 4882 5249 4918
rect 5254 4882 5257 5038
rect 5302 4942 5305 4948
rect 5250 4868 5254 4871
rect 5262 4852 5265 4858
rect 5278 4852 5281 4858
rect 5286 4822 5289 4858
rect 5302 4842 5305 4848
rect 5238 4792 5241 4818
rect 5262 4792 5265 4818
rect 5190 4762 5193 4768
rect 5242 4748 5246 4751
rect 5222 4732 5225 4738
rect 5166 4662 5169 4688
rect 5270 4682 5273 4738
rect 5194 4668 5198 4671
rect 5246 4662 5249 4668
rect 5078 4658 5089 4661
rect 5038 4652 5041 4658
rect 5054 4642 5057 4658
rect 5038 4551 5041 4618
rect 5054 4552 5057 4618
rect 5078 4552 5081 4648
rect 5038 4548 5049 4551
rect 5014 4532 5017 4548
rect 5034 4538 5038 4541
rect 5022 4532 5025 4538
rect 4990 4498 4998 4501
rect 4998 4482 5001 4488
rect 4986 4478 4990 4481
rect 5014 4472 5017 4528
rect 5030 4522 5033 4538
rect 4982 4442 4985 4458
rect 5006 4391 5009 4468
rect 5014 4452 5017 4458
rect 5014 4422 5017 4448
rect 5022 4442 5025 4448
rect 5006 4388 5017 4391
rect 4922 4348 4926 4351
rect 4910 4342 4913 4348
rect 5006 4342 5009 4348
rect 4936 4303 4938 4307
rect 4942 4303 4945 4307
rect 4949 4303 4952 4307
rect 4958 4282 4961 4288
rect 4754 4258 4758 4261
rect 4818 4258 4822 4261
rect 4850 4258 4854 4261
rect 4734 4172 4737 4178
rect 4734 4142 4737 4148
rect 4742 4142 4745 4178
rect 4766 4152 4769 4198
rect 4774 4152 4777 4228
rect 4782 4192 4785 4258
rect 4802 4248 4806 4251
rect 4798 4161 4801 4218
rect 4798 4158 4809 4161
rect 4754 4148 4758 4151
rect 4794 4148 4798 4151
rect 4806 4142 4809 4158
rect 4830 4151 4833 4258
rect 4926 4252 4929 4259
rect 4826 4148 4833 4151
rect 4694 4063 4697 4118
rect 4710 4082 4713 4118
rect 4726 4092 4729 4098
rect 4710 4072 4713 4078
rect 4670 3992 4673 4058
rect 4654 3952 4657 3988
rect 4726 3952 4729 3958
rect 4618 3948 4622 3951
rect 4642 3928 4646 3931
rect 4558 3888 4566 3891
rect 4598 3882 4601 3928
rect 4606 3872 4609 3878
rect 4550 3862 4553 3868
rect 4458 3858 4462 3861
rect 4494 3832 4497 3858
rect 4526 3852 4529 3858
rect 4510 3792 4513 3818
rect 4542 3772 4545 3858
rect 4402 3748 4406 3751
rect 4466 3748 4470 3751
rect 4494 3742 4497 3748
rect 4542 3742 4545 3748
rect 4506 3718 4510 3721
rect 4398 3682 4401 3718
rect 4414 3702 4417 3718
rect 4406 3682 4409 3688
rect 4414 3682 4417 3698
rect 4558 3692 4561 3748
rect 4574 3742 4577 3868
rect 4622 3862 4625 3908
rect 4606 3742 4609 3858
rect 4614 3762 4617 3818
rect 4630 3772 4633 3918
rect 4626 3758 4630 3761
rect 4618 3748 4622 3751
rect 4538 3688 4542 3691
rect 4446 3682 4449 3688
rect 4546 3678 4550 3681
rect 4342 3668 4353 3671
rect 4362 3668 4366 3671
rect 4242 3658 4246 3661
rect 4306 3658 4310 3661
rect 4242 3648 4246 3651
rect 4254 3642 4257 3658
rect 4270 3632 4273 3658
rect 4278 3652 4281 3658
rect 4318 3652 4321 3668
rect 4342 3662 4345 3668
rect 4354 3658 4358 3661
rect 4394 3658 4398 3661
rect 4170 3548 4174 3551
rect 4194 3548 4198 3551
rect 4162 3528 4166 3531
rect 4142 3502 4145 3518
rect 4190 3481 4193 3538
rect 4214 3532 4217 3548
rect 4222 3542 4225 3548
rect 4214 3512 4217 3518
rect 4262 3492 4265 3548
rect 4202 3488 4206 3491
rect 4190 3478 4201 3481
rect 4174 3472 4177 3478
rect 4146 3458 4150 3461
rect 4190 3432 4193 3468
rect 4130 3348 4134 3351
rect 4130 3328 4137 3331
rect 4078 3272 4081 3278
rect 4042 3268 4046 3271
rect 4042 3258 4046 3261
rect 4074 3258 4078 3261
rect 4054 3242 4057 3248
rect 3978 3068 3982 3071
rect 3998 3062 4001 3168
rect 4014 3132 4017 3147
rect 4030 3142 4033 3148
rect 4046 3132 4049 3158
rect 4042 3088 4046 3091
rect 4030 3072 4033 3088
rect 4038 3072 4041 3088
rect 3962 3058 3966 3061
rect 4026 3058 4030 3061
rect 3998 3042 4001 3058
rect 4006 3032 4009 3048
rect 4054 3032 4057 3238
rect 4062 3122 4065 3258
rect 4110 3162 4113 3188
rect 4102 3152 4105 3158
rect 4090 3148 4094 3151
rect 4118 3142 4121 3268
rect 4126 3262 4129 3268
rect 4134 3251 4137 3328
rect 4126 3248 4137 3251
rect 4126 3192 4129 3248
rect 4134 3152 4137 3228
rect 4142 3192 4145 3348
rect 4170 3338 4174 3341
rect 4178 3288 4182 3291
rect 4182 3232 4185 3258
rect 4142 3152 4145 3168
rect 4150 3152 4153 3198
rect 4130 3148 4134 3151
rect 4158 3141 4161 3148
rect 4138 3138 4161 3141
rect 4070 3132 4073 3138
rect 4118 3072 4121 3138
rect 4134 3082 4137 3088
rect 4166 3072 4169 3188
rect 4190 3171 4193 3328
rect 4198 3312 4201 3478
rect 4238 3472 4241 3488
rect 4270 3482 4273 3538
rect 4294 3482 4297 3508
rect 4310 3492 4313 3588
rect 4326 3552 4329 3558
rect 4350 3552 4353 3558
rect 4358 3542 4361 3618
rect 4366 3552 4369 3658
rect 4366 3542 4369 3548
rect 4398 3542 4401 3568
rect 4414 3552 4417 3658
rect 4424 3603 4426 3607
rect 4430 3603 4433 3607
rect 4437 3603 4440 3607
rect 4446 3592 4449 3648
rect 4462 3641 4465 3668
rect 4566 3662 4569 3668
rect 4574 3662 4577 3738
rect 4590 3682 4593 3688
rect 4622 3681 4625 3738
rect 4618 3678 4625 3681
rect 4638 3732 4641 3868
rect 4678 3832 4681 3948
rect 4734 3942 4737 4068
rect 4742 4022 4745 4128
rect 4750 4102 4753 4128
rect 4782 4062 4785 4118
rect 4822 4112 4825 4148
rect 4806 4072 4809 4078
rect 4830 4032 4833 4138
rect 4838 4132 4841 4158
rect 4846 4152 4849 4188
rect 4898 4158 4902 4161
rect 4870 4142 4873 4148
rect 4878 4142 4881 4148
rect 4918 4142 4921 4168
rect 4974 4152 4977 4268
rect 4914 4138 4918 4141
rect 4854 4042 4857 4138
rect 4894 4132 4897 4138
rect 4902 4132 4905 4138
rect 4936 4103 4938 4107
rect 4942 4103 4945 4107
rect 4949 4103 4952 4107
rect 4918 4072 4921 4078
rect 4890 4058 4894 4061
rect 4954 4028 4958 4031
rect 4742 3952 4745 4018
rect 4822 3992 4825 4018
rect 4786 3968 4790 3971
rect 4750 3952 4753 3968
rect 4686 3872 4689 3938
rect 4726 3872 4729 3918
rect 4686 3792 4689 3858
rect 4734 3832 4737 3858
rect 4654 3752 4657 3768
rect 4662 3742 4665 3748
rect 4650 3728 4654 3731
rect 4682 3728 4686 3731
rect 4630 3662 4633 3668
rect 4638 3662 4641 3728
rect 4702 3692 4705 3768
rect 4726 3752 4729 3758
rect 4714 3688 4718 3691
rect 4662 3682 4665 3688
rect 4678 3682 4681 3688
rect 4478 3652 4481 3659
rect 4606 3652 4609 3658
rect 4454 3638 4465 3641
rect 4378 3538 4382 3541
rect 4386 3528 4390 3531
rect 4334 3522 4337 3528
rect 4342 3522 4345 3528
rect 4394 3518 4398 3521
rect 4318 3512 4321 3518
rect 4338 3488 4342 3491
rect 4350 3482 4353 3518
rect 4406 3492 4409 3548
rect 4414 3542 4417 3548
rect 4454 3482 4457 3638
rect 4646 3632 4649 3658
rect 4462 3552 4465 3608
rect 4614 3592 4617 3618
rect 4558 3572 4561 3578
rect 4490 3558 4494 3561
rect 4506 3558 4510 3561
rect 4522 3558 4526 3561
rect 4534 3552 4537 3558
rect 4474 3548 4478 3551
rect 4250 3468 4254 3471
rect 4230 3452 4233 3458
rect 4214 3442 4217 3448
rect 4214 3432 4217 3438
rect 4198 3282 4201 3288
rect 4214 3282 4217 3428
rect 4238 3352 4241 3458
rect 4270 3451 4273 3478
rect 4366 3472 4369 3478
rect 4278 3462 4281 3468
rect 4270 3448 4281 3451
rect 4246 3342 4249 3348
rect 4226 3268 4230 3271
rect 4254 3262 4257 3348
rect 4278 3342 4281 3448
rect 4302 3392 4305 3468
rect 4326 3422 4329 3458
rect 4310 3362 4313 3418
rect 4298 3338 4302 3341
rect 4278 3332 4281 3338
rect 4270 3292 4273 3308
rect 4286 3262 4289 3278
rect 4294 3272 4297 3308
rect 4334 3292 4337 3468
rect 4382 3352 4385 3459
rect 4424 3403 4426 3407
rect 4430 3403 4433 3407
rect 4437 3403 4440 3407
rect 4446 3391 4449 3418
rect 4438 3388 4449 3391
rect 4406 3372 4409 3378
rect 4438 3372 4441 3388
rect 4390 3362 4393 3368
rect 4350 3348 4358 3351
rect 4350 3322 4353 3348
rect 4366 3342 4369 3348
rect 4358 3332 4361 3338
rect 4398 3332 4401 3338
rect 4202 3258 4206 3261
rect 4262 3252 4265 3258
rect 4270 3242 4273 3248
rect 4190 3168 4201 3171
rect 4178 3148 4182 3151
rect 4182 3132 4185 3138
rect 4190 3062 4193 3158
rect 4198 3072 4201 3168
rect 4238 3092 4241 3098
rect 4102 3052 4105 3059
rect 4202 3058 4206 3061
rect 4226 3058 4230 3061
rect 4170 3048 4174 3051
rect 3920 2903 3922 2907
rect 3926 2903 3929 2907
rect 3933 2903 3936 2907
rect 3910 2772 3913 2778
rect 3942 2761 3945 2948
rect 3954 2938 3958 2941
rect 3974 2932 3977 2958
rect 3986 2948 3990 2951
rect 3978 2928 3982 2931
rect 3958 2922 3961 2928
rect 3998 2902 4001 3018
rect 4006 2972 4009 2978
rect 4022 2962 4025 3018
rect 4062 2992 4065 3018
rect 4050 2958 4054 2961
rect 4086 2952 4089 3038
rect 4022 2942 4025 2948
rect 4078 2942 4081 2948
rect 4134 2942 4137 3028
rect 4158 2962 4161 2968
rect 3942 2758 3953 2761
rect 3950 2752 3953 2758
rect 3890 2748 3894 2751
rect 3750 2652 3753 2658
rect 3830 2652 3833 2658
rect 3750 2612 3753 2648
rect 3750 2562 3753 2568
rect 3702 2542 3705 2548
rect 3734 2542 3737 2548
rect 3750 2532 3753 2538
rect 3766 2521 3769 2618
rect 3778 2548 3782 2551
rect 3778 2528 3782 2531
rect 3766 2518 3777 2521
rect 3718 2492 3721 2518
rect 3766 2492 3769 2508
rect 3702 2472 3705 2478
rect 3710 2472 3713 2478
rect 3718 2452 3721 2488
rect 3742 2472 3745 2488
rect 3662 2432 3665 2448
rect 3694 2432 3697 2448
rect 3734 2442 3737 2458
rect 3750 2452 3753 2468
rect 3774 2451 3777 2518
rect 3770 2448 3777 2451
rect 3782 2452 3785 2458
rect 3662 2352 3665 2398
rect 3614 2252 3617 2268
rect 3622 2262 3625 2268
rect 3638 2242 3641 2268
rect 3662 2262 3665 2338
rect 3670 2302 3673 2338
rect 3630 2152 3633 2168
rect 3614 2112 3617 2118
rect 3614 2082 3617 2098
rect 3646 2092 3649 2218
rect 3654 2192 3657 2218
rect 3662 2092 3665 2198
rect 3678 2092 3681 2418
rect 3686 2392 3689 2408
rect 3694 2352 3697 2388
rect 3726 2362 3729 2418
rect 3734 2382 3737 2418
rect 3742 2402 3745 2428
rect 3742 2361 3745 2388
rect 3766 2382 3769 2388
rect 3734 2358 3745 2361
rect 3686 2342 3689 2348
rect 3734 2341 3737 2358
rect 3746 2348 3750 2351
rect 3758 2342 3761 2378
rect 3734 2338 3750 2341
rect 3690 2328 3710 2331
rect 3750 2292 3753 2318
rect 3766 2292 3769 2348
rect 3774 2312 3777 2448
rect 3790 2382 3793 2568
rect 3798 2542 3801 2618
rect 3846 2562 3849 2658
rect 3854 2652 3857 2668
rect 3862 2662 3865 2668
rect 3870 2662 3873 2748
rect 3942 2741 3945 2748
rect 3958 2742 3961 2758
rect 3966 2742 3969 2898
rect 4022 2892 4025 2938
rect 4030 2932 4033 2938
rect 4106 2928 4110 2931
rect 3990 2872 3993 2878
rect 3998 2862 4001 2868
rect 4018 2858 4022 2861
rect 4034 2858 4038 2861
rect 3982 2822 3985 2858
rect 4046 2852 4049 2918
rect 4054 2872 4057 2898
rect 4094 2882 4097 2918
rect 4118 2892 4121 2918
rect 4126 2902 4129 2928
rect 4034 2848 4038 2851
rect 3982 2742 3985 2818
rect 3942 2738 3953 2741
rect 3878 2732 3881 2738
rect 3906 2718 3910 2721
rect 3920 2703 3922 2707
rect 3926 2703 3929 2707
rect 3933 2703 3936 2707
rect 3942 2692 3945 2728
rect 3950 2692 3953 2738
rect 3882 2668 3886 2671
rect 3862 2592 3865 2648
rect 3870 2561 3873 2658
rect 3878 2642 3881 2658
rect 3870 2558 3881 2561
rect 3810 2548 3814 2551
rect 3870 2542 3873 2548
rect 3878 2542 3881 2558
rect 3806 2472 3809 2538
rect 3814 2512 3817 2518
rect 3790 2362 3793 2368
rect 3806 2352 3809 2378
rect 3814 2352 3817 2358
rect 3814 2332 3817 2338
rect 3778 2288 3782 2291
rect 3722 2268 3726 2271
rect 3734 2270 3737 2288
rect 3782 2282 3785 2288
rect 3754 2278 3758 2281
rect 3778 2258 3782 2261
rect 3702 2142 3705 2148
rect 3710 2142 3713 2238
rect 3718 2202 3721 2218
rect 3766 2171 3769 2188
rect 3774 2182 3777 2188
rect 3766 2168 3777 2171
rect 3710 2092 3713 2118
rect 3734 2092 3737 2108
rect 3774 2092 3777 2168
rect 3814 2161 3817 2298
rect 3822 2182 3825 2518
rect 3830 2482 3833 2508
rect 3834 2468 3838 2471
rect 3846 2362 3849 2418
rect 3838 2352 3841 2358
rect 3830 2322 3833 2348
rect 3846 2281 3849 2348
rect 3854 2332 3857 2528
rect 3870 2502 3873 2528
rect 3870 2452 3873 2498
rect 3862 2432 3865 2448
rect 3878 2372 3881 2538
rect 3894 2482 3897 2678
rect 3934 2672 3937 2678
rect 3902 2492 3905 2508
rect 3894 2472 3897 2478
rect 3890 2458 3894 2461
rect 3890 2448 3902 2451
rect 3854 2302 3857 2328
rect 3838 2278 3849 2281
rect 3862 2292 3865 2368
rect 3878 2352 3881 2358
rect 3870 2342 3873 2348
rect 3886 2332 3889 2438
rect 3910 2402 3913 2668
rect 3950 2662 3953 2678
rect 3958 2672 3961 2688
rect 3966 2682 3969 2738
rect 3978 2728 3982 2731
rect 3966 2572 3969 2678
rect 3974 2672 3977 2718
rect 3978 2548 3982 2551
rect 3958 2542 3961 2548
rect 3926 2522 3929 2528
rect 3920 2503 3922 2507
rect 3926 2503 3929 2507
rect 3933 2503 3936 2507
rect 3930 2468 3934 2471
rect 3918 2452 3921 2458
rect 3894 2352 3897 2398
rect 3910 2352 3913 2398
rect 3918 2382 3921 2448
rect 3958 2362 3961 2418
rect 3954 2348 3958 2351
rect 3838 2252 3841 2278
rect 3862 2272 3865 2288
rect 3878 2262 3881 2268
rect 3846 2242 3849 2259
rect 3886 2251 3889 2298
rect 3894 2262 3897 2268
rect 3882 2248 3889 2251
rect 3862 2172 3865 2198
rect 3902 2192 3905 2338
rect 3910 2302 3913 2348
rect 3954 2338 3958 2341
rect 3930 2328 3934 2331
rect 3920 2303 3922 2307
rect 3926 2303 3929 2307
rect 3933 2303 3936 2307
rect 3926 2288 3945 2291
rect 3926 2281 3929 2288
rect 3910 2278 3929 2281
rect 3910 2272 3913 2278
rect 3922 2268 3926 2271
rect 3910 2192 3913 2258
rect 3806 2158 3817 2161
rect 3786 2138 3790 2141
rect 3622 2072 3625 2078
rect 3602 2058 3606 2061
rect 3526 1902 3529 1948
rect 3538 1938 3542 1941
rect 3582 1932 3585 1938
rect 3518 1872 3521 1878
rect 3526 1862 3529 1868
rect 3454 1822 3457 1848
rect 3400 1803 3402 1807
rect 3406 1803 3409 1807
rect 3413 1803 3416 1807
rect 3438 1752 3441 1768
rect 3470 1752 3473 1818
rect 3502 1792 3505 1838
rect 3518 1762 3521 1778
rect 3490 1758 3494 1761
rect 3342 1742 3345 1748
rect 3506 1748 3510 1751
rect 3514 1748 3518 1751
rect 3294 1732 3297 1738
rect 3358 1732 3361 1738
rect 3302 1663 3305 1688
rect 3334 1672 3337 1678
rect 3342 1672 3345 1728
rect 3390 1692 3393 1738
rect 3362 1688 3366 1691
rect 3302 1658 3305 1659
rect 3334 1592 3337 1658
rect 3350 1652 3353 1658
rect 3374 1652 3377 1668
rect 3414 1662 3417 1708
rect 3462 1692 3465 1738
rect 3470 1682 3473 1748
rect 3526 1732 3529 1828
rect 3534 1742 3537 1858
rect 3550 1761 3553 1918
rect 3558 1902 3561 1918
rect 3582 1872 3585 1888
rect 3598 1882 3601 1948
rect 3606 1942 3609 1948
rect 3614 1931 3617 2038
rect 3630 1982 3633 2058
rect 3646 2052 3649 2058
rect 3642 2048 3646 2051
rect 3654 2042 3657 2078
rect 3638 1942 3641 1948
rect 3606 1928 3617 1931
rect 3634 1928 3638 1931
rect 3606 1892 3609 1928
rect 3614 1882 3617 1888
rect 3622 1872 3625 1878
rect 3598 1862 3601 1868
rect 3590 1851 3593 1858
rect 3590 1848 3601 1851
rect 3550 1758 3561 1761
rect 3558 1752 3561 1758
rect 3566 1752 3569 1838
rect 3546 1748 3550 1751
rect 3542 1732 3545 1738
rect 3486 1682 3489 1688
rect 3422 1662 3425 1668
rect 3446 1662 3449 1668
rect 3478 1662 3481 1668
rect 3402 1658 3406 1661
rect 3254 1552 3257 1558
rect 3222 1548 3230 1551
rect 3338 1548 3342 1551
rect 3190 1512 3193 1538
rect 3066 1458 3070 1461
rect 2958 1352 2961 1368
rect 3054 1362 3057 1368
rect 3070 1352 3073 1378
rect 3010 1348 3014 1351
rect 3050 1348 3054 1351
rect 3078 1351 3081 1428
rect 3102 1392 3105 1448
rect 3118 1392 3121 1458
rect 3126 1402 3129 1458
rect 3134 1442 3137 1458
rect 3150 1452 3153 1498
rect 3166 1452 3169 1458
rect 3174 1392 3177 1468
rect 3158 1362 3161 1368
rect 3174 1362 3177 1368
rect 3146 1358 3150 1361
rect 3078 1348 3086 1351
rect 3130 1348 3134 1351
rect 2966 1342 2969 1348
rect 2990 1332 2993 1348
rect 3038 1342 3041 1348
rect 3058 1338 3062 1341
rect 3070 1312 3073 1348
rect 3078 1302 3081 1338
rect 2958 1262 2961 1278
rect 2966 1272 2969 1288
rect 2982 1262 2985 1268
rect 2946 1258 2950 1261
rect 3086 1262 3089 1348
rect 3142 1342 3145 1348
rect 3102 1292 3105 1298
rect 3118 1292 3121 1338
rect 3150 1322 3153 1338
rect 3094 1262 3097 1268
rect 3150 1262 3153 1268
rect 3158 1262 3161 1348
rect 3190 1342 3193 1508
rect 3206 1502 3209 1528
rect 3222 1412 3225 1548
rect 3286 1542 3289 1548
rect 3258 1538 3262 1541
rect 3354 1538 3358 1541
rect 3302 1532 3305 1538
rect 3230 1462 3233 1518
rect 3206 1342 3209 1347
rect 3182 1263 3185 1288
rect 3214 1272 3217 1338
rect 3238 1321 3241 1458
rect 3234 1318 3241 1321
rect 3234 1288 3238 1291
rect 3254 1272 3257 1498
rect 3262 1472 3265 1528
rect 3270 1512 3273 1518
rect 3294 1492 3297 1498
rect 3310 1492 3313 1528
rect 3326 1482 3329 1508
rect 3342 1492 3345 1528
rect 3278 1462 3281 1478
rect 3366 1472 3369 1608
rect 3382 1582 3385 1658
rect 3390 1652 3393 1658
rect 3400 1603 3402 1607
rect 3406 1603 3409 1607
rect 3413 1603 3416 1607
rect 3374 1562 3377 1568
rect 3382 1502 3385 1578
rect 3430 1532 3433 1548
rect 3354 1458 3358 1461
rect 3310 1442 3313 1458
rect 3366 1442 3369 1468
rect 3270 1362 3273 1368
rect 3270 1342 3273 1358
rect 3294 1352 3297 1358
rect 3302 1332 3305 1358
rect 3270 1328 3278 1331
rect 3002 1259 3006 1261
rect 2998 1258 3006 1259
rect 3074 1258 3078 1261
rect 3222 1262 3225 1268
rect 3246 1262 3249 1268
rect 2938 1248 2942 1251
rect 2878 1162 2881 1218
rect 2862 1152 2865 1158
rect 2842 1148 2846 1151
rect 2894 1142 2897 1148
rect 2818 1138 2822 1141
rect 2906 1138 2910 1141
rect 2810 1128 2814 1131
rect 2766 1088 2785 1091
rect 2766 1072 2769 1088
rect 2782 1082 2785 1088
rect 2750 1038 2761 1041
rect 2774 1062 2777 1078
rect 2782 1062 2785 1068
rect 2814 1063 2817 1078
rect 2774 1042 2777 1058
rect 2586 968 2590 971
rect 2606 962 2609 1028
rect 2750 992 2753 1038
rect 2838 1032 2841 1058
rect 2514 878 2518 881
rect 2530 868 2534 871
rect 2494 771 2497 838
rect 2494 768 2505 771
rect 2502 742 2505 768
rect 2542 752 2545 868
rect 2558 862 2561 958
rect 2606 952 2609 958
rect 2630 952 2633 968
rect 2670 962 2673 978
rect 2718 972 2721 978
rect 2638 952 2641 958
rect 2650 948 2654 951
rect 2598 942 2601 948
rect 2650 938 2654 941
rect 2590 862 2593 868
rect 2550 842 2553 858
rect 2582 812 2585 858
rect 2590 772 2593 858
rect 2598 832 2601 868
rect 2606 862 2609 918
rect 2638 892 2641 918
rect 2618 848 2622 851
rect 2598 792 2601 808
rect 2486 732 2489 738
rect 2486 682 2489 718
rect 2510 682 2513 688
rect 2506 678 2510 681
rect 2566 681 2569 768
rect 2606 732 2609 848
rect 2630 792 2633 848
rect 2646 812 2649 868
rect 2654 862 2657 938
rect 2654 832 2657 858
rect 2614 752 2617 758
rect 2630 752 2633 788
rect 2638 762 2641 768
rect 2642 748 2646 751
rect 2626 738 2630 741
rect 2606 722 2609 728
rect 2566 678 2574 681
rect 2486 662 2489 678
rect 2574 663 2577 668
rect 2474 658 2478 661
rect 2494 592 2497 658
rect 2502 592 2505 628
rect 2482 558 2486 561
rect 2502 552 2505 588
rect 2510 572 2513 598
rect 2470 492 2473 528
rect 2502 512 2505 538
rect 2510 532 2513 568
rect 2570 547 2574 550
rect 2558 472 2561 538
rect 2574 492 2577 508
rect 2574 482 2577 488
rect 2534 462 2537 468
rect 2458 448 2462 451
rect 2446 442 2449 448
rect 2474 438 2478 441
rect 2462 352 2465 358
rect 2450 348 2454 351
rect 2458 338 2462 341
rect 2470 292 2473 428
rect 2426 268 2430 271
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2397 203 2400 207
rect 2398 172 2401 178
rect 2358 142 2361 148
rect 2430 142 2433 258
rect 2454 252 2457 288
rect 2478 272 2481 298
rect 2474 268 2478 271
rect 2486 262 2489 278
rect 2518 272 2521 458
rect 2558 442 2561 468
rect 2542 342 2545 348
rect 2566 342 2569 438
rect 2590 392 2593 698
rect 2606 672 2609 678
rect 2654 672 2657 748
rect 2662 742 2665 958
rect 2682 948 2686 951
rect 2694 942 2697 968
rect 2738 958 2742 961
rect 2714 948 2718 951
rect 2758 951 2761 1008
rect 2806 992 2809 1018
rect 2830 962 2833 978
rect 2754 948 2761 951
rect 2786 958 2790 961
rect 2702 942 2705 948
rect 2750 942 2753 948
rect 2710 922 2713 938
rect 2726 882 2729 898
rect 2698 878 2702 881
rect 2714 858 2718 861
rect 2726 742 2729 878
rect 2742 822 2745 938
rect 2758 852 2761 918
rect 2766 892 2769 958
rect 2806 952 2809 958
rect 2778 938 2782 941
rect 2790 931 2793 938
rect 2782 928 2793 931
rect 2774 872 2777 878
rect 2782 752 2785 928
rect 2790 751 2793 918
rect 2838 902 2841 1028
rect 2846 932 2849 1128
rect 2870 1122 2873 1138
rect 2886 1131 2889 1138
rect 2886 1128 2910 1131
rect 2854 942 2857 958
rect 2846 892 2849 928
rect 2818 868 2822 871
rect 2798 862 2801 868
rect 2810 858 2814 861
rect 2830 832 2833 858
rect 2814 752 2817 828
rect 2822 752 2825 798
rect 2838 752 2841 758
rect 2854 752 2857 878
rect 2862 872 2865 1118
rect 2888 1103 2890 1107
rect 2894 1103 2897 1107
rect 2901 1103 2904 1107
rect 2870 952 2873 1098
rect 2882 1088 2886 1091
rect 2878 1072 2881 1088
rect 2910 1062 2913 1068
rect 2918 972 2921 1148
rect 2926 1062 2929 1198
rect 2950 1192 2953 1238
rect 2958 1222 2961 1258
rect 3050 1248 3054 1251
rect 2986 1158 2990 1161
rect 3014 1152 3017 1208
rect 3030 1192 3033 1218
rect 3046 1162 3049 1168
rect 3070 1162 3073 1188
rect 3078 1162 3081 1228
rect 3126 1182 3129 1188
rect 3106 1158 3110 1161
rect 3002 1148 3006 1151
rect 3026 1148 3030 1151
rect 3138 1148 3142 1151
rect 2958 1142 2961 1148
rect 2950 1122 2953 1128
rect 2966 1092 2969 1148
rect 2982 1062 2985 1148
rect 3014 1142 3017 1148
rect 3050 1138 3054 1141
rect 2938 1058 2942 1061
rect 2914 958 2918 961
rect 2870 942 2873 948
rect 2898 938 2902 941
rect 2890 928 2894 931
rect 2888 903 2890 907
rect 2894 903 2897 907
rect 2901 903 2904 907
rect 2862 862 2865 868
rect 2910 832 2913 948
rect 2926 892 2929 1058
rect 2966 1032 2969 1058
rect 2942 972 2945 1028
rect 2958 972 2961 1018
rect 2934 862 2937 888
rect 2942 862 2945 968
rect 2966 932 2969 948
rect 2974 942 2977 1058
rect 2982 932 2985 1058
rect 2990 1022 2993 1058
rect 3006 1032 3009 1138
rect 3022 1122 3025 1138
rect 3038 1072 3041 1078
rect 3022 1062 3025 1068
rect 3022 992 3025 1028
rect 3054 962 3057 1138
rect 3082 1118 3086 1121
rect 3070 1092 3073 1118
rect 3094 1112 3097 1148
rect 3070 952 3073 1068
rect 3082 1058 3086 1061
rect 3102 972 3105 1138
rect 3126 1061 3129 1148
rect 3150 1142 3153 1208
rect 3158 1142 3161 1258
rect 3214 1212 3217 1258
rect 3262 1242 3265 1278
rect 3270 1252 3273 1328
rect 3298 1318 3305 1321
rect 3278 1262 3281 1268
rect 3286 1262 3289 1298
rect 3302 1292 3305 1318
rect 3294 1252 3297 1258
rect 3230 1192 3233 1198
rect 3246 1162 3249 1178
rect 3278 1152 3281 1158
rect 3250 1148 3254 1151
rect 3266 1148 3270 1151
rect 3134 1122 3137 1138
rect 3166 1132 3169 1148
rect 3286 1141 3289 1148
rect 3282 1138 3289 1141
rect 3174 1132 3177 1138
rect 3270 1132 3273 1138
rect 3158 1112 3161 1118
rect 3230 1112 3233 1118
rect 3146 1088 3150 1091
rect 3134 1082 3137 1088
rect 3206 1082 3209 1108
rect 3206 1063 3209 1068
rect 3126 1058 3137 1061
rect 3134 992 3137 1058
rect 3238 1032 3241 1068
rect 3246 1062 3249 1068
rect 3254 1062 3257 1068
rect 3262 1062 3265 1078
rect 3270 1052 3273 1088
rect 3286 1062 3289 1118
rect 3294 1072 3297 1218
rect 3310 1212 3313 1438
rect 3318 1332 3321 1358
rect 3326 1342 3329 1378
rect 3354 1358 3358 1361
rect 3366 1352 3369 1398
rect 3390 1392 3393 1518
rect 3430 1462 3433 1488
rect 3438 1462 3441 1538
rect 3470 1492 3473 1498
rect 3478 1472 3481 1558
rect 3502 1552 3505 1598
rect 3518 1562 3521 1728
rect 3558 1672 3561 1748
rect 3566 1682 3569 1748
rect 3586 1738 3590 1741
rect 3598 1692 3601 1848
rect 3630 1762 3633 1928
rect 3646 1912 3649 1918
rect 3638 1872 3641 1878
rect 3654 1872 3657 1938
rect 3670 1932 3673 2068
rect 3678 2062 3681 2078
rect 3726 2072 3729 2088
rect 3758 2072 3761 2078
rect 3686 2052 3689 2068
rect 3718 2062 3721 2068
rect 3706 2058 3710 2061
rect 3738 2058 3742 2061
rect 3694 2032 3697 2058
rect 3670 1902 3673 1918
rect 3678 1891 3681 1918
rect 3670 1888 3681 1891
rect 3646 1862 3649 1868
rect 3670 1862 3673 1888
rect 3686 1882 3689 1898
rect 3678 1871 3681 1878
rect 3678 1868 3686 1871
rect 3694 1862 3697 1868
rect 3678 1852 3681 1858
rect 3670 1832 3673 1848
rect 3606 1732 3609 1738
rect 3630 1691 3633 1758
rect 3650 1748 3654 1751
rect 3670 1742 3673 1748
rect 3622 1688 3633 1691
rect 3638 1692 3641 1698
rect 3614 1672 3617 1688
rect 3622 1662 3625 1688
rect 3630 1672 3633 1678
rect 3646 1672 3649 1678
rect 3662 1662 3665 1678
rect 3554 1658 3558 1661
rect 3650 1658 3654 1661
rect 3666 1658 3670 1661
rect 3546 1548 3550 1551
rect 3490 1538 3494 1541
rect 3486 1512 3489 1518
rect 3490 1488 3494 1491
rect 3474 1458 3478 1461
rect 3438 1452 3441 1458
rect 3400 1403 3402 1407
rect 3406 1403 3409 1407
rect 3413 1403 3416 1407
rect 3378 1358 3382 1361
rect 3334 1342 3337 1348
rect 3390 1342 3393 1388
rect 3398 1352 3401 1368
rect 3438 1362 3441 1428
rect 3454 1362 3457 1368
rect 3418 1358 3422 1361
rect 3406 1352 3409 1358
rect 3362 1338 3366 1341
rect 3378 1338 3382 1341
rect 3318 1282 3321 1288
rect 3334 1252 3337 1258
rect 3310 1192 3313 1208
rect 3350 1162 3353 1318
rect 3306 1158 3310 1161
rect 3358 1152 3361 1158
rect 3366 1152 3369 1208
rect 3374 1202 3377 1268
rect 3382 1262 3385 1268
rect 3390 1222 3393 1338
rect 3434 1328 3438 1331
rect 3462 1282 3465 1288
rect 3478 1282 3481 1458
rect 3502 1382 3505 1548
rect 3526 1542 3529 1548
rect 3534 1522 3537 1528
rect 3558 1512 3561 1528
rect 3526 1482 3529 1498
rect 3510 1462 3513 1468
rect 3542 1452 3545 1468
rect 3502 1342 3505 1348
rect 3542 1342 3545 1448
rect 3566 1432 3569 1558
rect 3574 1552 3577 1618
rect 3598 1592 3601 1648
rect 3622 1592 3625 1658
rect 3670 1592 3673 1648
rect 3678 1642 3681 1848
rect 3694 1812 3697 1858
rect 3702 1851 3705 1908
rect 3710 1862 3713 1868
rect 3718 1852 3721 1948
rect 3730 1947 3734 1950
rect 3750 1921 3753 2058
rect 3790 2052 3793 2058
rect 3782 2002 3785 2048
rect 3750 1918 3761 1921
rect 3750 1872 3753 1878
rect 3726 1862 3729 1868
rect 3702 1848 3710 1851
rect 3694 1662 3697 1758
rect 3718 1692 3721 1848
rect 3734 1842 3737 1868
rect 3730 1818 3734 1821
rect 3750 1742 3753 1748
rect 3742 1682 3745 1738
rect 3710 1672 3713 1678
rect 3706 1658 3710 1661
rect 3622 1562 3625 1588
rect 3650 1558 3654 1561
rect 3590 1542 3593 1548
rect 3574 1532 3577 1538
rect 3582 1531 3585 1538
rect 3606 1532 3609 1548
rect 3622 1542 3625 1558
rect 3582 1528 3593 1531
rect 3582 1452 3585 1458
rect 3590 1432 3593 1528
rect 3638 1502 3641 1548
rect 3646 1522 3649 1538
rect 3654 1492 3657 1558
rect 3678 1552 3681 1618
rect 3694 1562 3697 1658
rect 3742 1592 3745 1668
rect 3750 1662 3753 1668
rect 3758 1632 3761 1918
rect 3774 1892 3777 1948
rect 3798 1922 3801 2108
rect 3806 2092 3809 2158
rect 3838 2152 3841 2158
rect 3834 2148 3838 2151
rect 3814 2112 3817 2148
rect 3822 2122 3825 2148
rect 3862 2142 3865 2148
rect 3834 2138 3838 2141
rect 3806 2072 3809 2088
rect 3818 2078 3822 2081
rect 3838 2062 3841 2068
rect 3870 2062 3873 2188
rect 3934 2182 3937 2278
rect 3942 2272 3945 2288
rect 3966 2262 3969 2368
rect 3974 2352 3977 2528
rect 3990 2492 3993 2798
rect 3998 2752 4001 2838
rect 4022 2762 4025 2768
rect 3998 2702 4001 2748
rect 4022 2742 4025 2748
rect 4038 2742 4041 2768
rect 4046 2762 4049 2818
rect 4062 2772 4065 2818
rect 4090 2758 4094 2761
rect 4050 2748 4054 2751
rect 4090 2748 4094 2751
rect 4078 2732 4081 2748
rect 4094 2722 4097 2728
rect 4062 2712 4065 2718
rect 4014 2662 4017 2668
rect 3998 2652 4001 2658
rect 4022 2552 4025 2618
rect 4038 2592 4041 2678
rect 4102 2662 4105 2858
rect 4126 2802 4129 2859
rect 4142 2821 4145 2948
rect 4182 2941 4185 3058
rect 4222 3012 4225 3048
rect 4198 2962 4201 2998
rect 4218 2968 4222 2971
rect 4202 2948 4206 2951
rect 4182 2938 4190 2941
rect 4194 2938 4198 2941
rect 4174 2932 4177 2938
rect 4190 2892 4193 2898
rect 4170 2888 4174 2891
rect 4158 2882 4161 2888
rect 4174 2872 4177 2878
rect 4162 2868 4166 2871
rect 4178 2858 4182 2861
rect 4134 2818 4145 2821
rect 4110 2752 4113 2758
rect 4118 2742 4121 2788
rect 4126 2762 4129 2768
rect 4134 2692 4137 2818
rect 4146 2758 4158 2761
rect 4166 2752 4169 2798
rect 4174 2752 4177 2758
rect 4182 2752 4185 2858
rect 4194 2788 4198 2791
rect 4206 2762 4209 2918
rect 4222 2862 4225 2868
rect 4230 2862 4233 2888
rect 4142 2702 4145 2748
rect 4182 2742 4185 2748
rect 4102 2652 4105 2658
rect 4062 2642 4065 2648
rect 4062 2592 4065 2628
rect 4102 2592 4105 2618
rect 4062 2502 4065 2518
rect 4070 2482 4073 2548
rect 4058 2468 4062 2471
rect 4034 2458 4038 2461
rect 3982 2452 3985 2458
rect 4006 2452 4009 2458
rect 4046 2422 4049 2468
rect 4078 2462 4081 2548
rect 4094 2472 4097 2508
rect 4110 2492 4113 2588
rect 4118 2532 4121 2688
rect 4150 2682 4153 2738
rect 4198 2732 4201 2758
rect 4134 2663 4137 2668
rect 4150 2602 4153 2678
rect 4166 2662 4169 2668
rect 4198 2662 4201 2678
rect 4214 2662 4217 2668
rect 4222 2662 4225 2758
rect 4230 2752 4233 2768
rect 4238 2762 4241 2848
rect 4254 2752 4257 3208
rect 4286 3162 4289 3258
rect 4302 3232 4305 3268
rect 4262 3132 4265 3148
rect 4286 3142 4289 3148
rect 4262 3072 4265 3078
rect 4270 3062 4273 3098
rect 4302 3062 4305 3148
rect 4310 3102 4313 3258
rect 4326 3251 4329 3268
rect 4334 3262 4337 3288
rect 4342 3262 4345 3268
rect 4350 3262 4353 3318
rect 4362 3288 4366 3291
rect 4326 3248 4334 3251
rect 4318 3192 4321 3248
rect 4350 3172 4353 3258
rect 4358 3202 4361 3268
rect 4398 3232 4401 3328
rect 4406 3252 4409 3348
rect 4462 3272 4465 3548
rect 4478 3532 4481 3538
rect 4470 3472 4473 3498
rect 4486 3472 4489 3548
rect 4494 3462 4497 3518
rect 4510 3512 4513 3538
rect 4518 3502 4521 3548
rect 4494 3452 4497 3458
rect 4470 3392 4473 3398
rect 4486 3362 4489 3368
rect 4494 3362 4497 3448
rect 4502 3382 4505 3418
rect 4542 3382 4545 3558
rect 4554 3548 4558 3551
rect 4566 3542 4569 3568
rect 4578 3558 4582 3561
rect 4598 3552 4601 3558
rect 4630 3552 4633 3598
rect 4646 3582 4649 3618
rect 4662 3592 4665 3648
rect 4686 3642 4689 3658
rect 4670 3552 4673 3618
rect 4690 3558 4694 3561
rect 4650 3548 4654 3551
rect 4606 3542 4609 3548
rect 4638 3542 4641 3548
rect 4618 3538 4622 3541
rect 4626 3538 4633 3541
rect 4574 3522 4577 3528
rect 4590 3502 4593 3538
rect 4582 3472 4585 3478
rect 4606 3472 4609 3528
rect 4566 3392 4569 3459
rect 4610 3458 4614 3461
rect 4598 3442 4601 3448
rect 4518 3372 4521 3378
rect 4538 3358 4550 3361
rect 4566 3352 4569 3378
rect 4610 3368 4614 3371
rect 4502 3342 4505 3348
rect 4550 3342 4553 3348
rect 4590 3342 4593 3348
rect 4478 3302 4481 3338
rect 4478 3292 4481 3298
rect 4486 3292 4489 3308
rect 4482 3268 4486 3271
rect 4418 3258 4422 3261
rect 4424 3203 4426 3207
rect 4430 3203 4433 3207
rect 4437 3203 4440 3207
rect 4358 3162 4361 3168
rect 4346 3158 4350 3161
rect 4334 3142 4337 3158
rect 4374 3152 4377 3188
rect 4382 3142 4385 3188
rect 4430 3152 4433 3158
rect 4438 3152 4441 3158
rect 4418 3148 4422 3151
rect 4446 3142 4449 3268
rect 4482 3258 4486 3261
rect 4494 3261 4497 3338
rect 4530 3288 4534 3291
rect 4518 3272 4521 3288
rect 4542 3282 4545 3338
rect 4542 3272 4545 3278
rect 4510 3262 4513 3268
rect 4494 3258 4502 3261
rect 4470 3222 4473 3228
rect 4462 3152 4465 3208
rect 4470 3142 4473 3218
rect 4494 3172 4497 3198
rect 4518 3182 4521 3268
rect 4550 3262 4553 3338
rect 4574 3262 4577 3338
rect 4582 3332 4585 3338
rect 4582 3282 4585 3328
rect 4542 3258 4550 3261
rect 4534 3252 4537 3258
rect 4542 3252 4545 3258
rect 4566 3242 4569 3248
rect 4582 3202 4585 3278
rect 4590 3262 4593 3268
rect 4598 3262 4601 3268
rect 4614 3262 4617 3318
rect 4622 3282 4625 3468
rect 4630 3442 4633 3538
rect 4638 3352 4641 3418
rect 4630 3322 4633 3348
rect 4638 3342 4641 3348
rect 4646 3342 4649 3498
rect 4694 3492 4697 3528
rect 4702 3512 4705 3618
rect 4734 3552 4737 3828
rect 4742 3772 4745 3948
rect 4766 3872 4769 3968
rect 4822 3962 4825 3968
rect 4802 3958 4806 3961
rect 4802 3948 4806 3951
rect 4790 3922 4793 3938
rect 4838 3872 4841 3948
rect 4846 3942 4849 4008
rect 4846 3932 4849 3938
rect 4854 3932 4857 3958
rect 4870 3952 4873 3978
rect 4906 3958 4910 3961
rect 4950 3952 4953 4028
rect 4966 3952 4969 4088
rect 4982 3971 4985 4278
rect 5014 4272 5017 4388
rect 5030 4362 5033 4518
rect 5046 4501 5049 4548
rect 5038 4498 5049 4501
rect 5038 4382 5041 4498
rect 5046 4362 5049 4368
rect 5030 4342 5033 4348
rect 5046 4322 5049 4328
rect 5054 4282 5057 4548
rect 5078 4542 5081 4548
rect 5062 4372 5065 4478
rect 5078 4462 5081 4488
rect 5062 4352 5065 4358
rect 5062 4272 5065 4348
rect 5070 4322 5073 4338
rect 5078 4282 5081 4318
rect 5010 4268 5014 4271
rect 4990 4262 4993 4268
rect 5022 4262 5025 4268
rect 5054 4262 5057 4268
rect 5062 4262 5065 4268
rect 5010 4258 5014 4261
rect 5022 4232 5025 4258
rect 5030 4212 5033 4248
rect 5046 4242 5049 4258
rect 4994 4148 4998 4151
rect 5006 4072 5009 4128
rect 5046 4122 5049 4218
rect 5070 4172 5073 4218
rect 5074 4148 5078 4151
rect 5046 4072 5049 4078
rect 5014 4052 5017 4059
rect 5050 4058 5054 4061
rect 5054 4042 5057 4048
rect 5078 4032 5081 4038
rect 5086 4021 5089 4658
rect 5094 4532 5097 4598
rect 5102 4531 5105 4658
rect 5118 4642 5121 4658
rect 5142 4652 5145 4658
rect 5142 4582 5145 4588
rect 5118 4552 5121 4568
rect 5150 4562 5153 4658
rect 5190 4592 5193 4658
rect 5190 4572 5193 4588
rect 5206 4562 5209 4618
rect 5114 4538 5118 4541
rect 5102 4528 5113 4531
rect 5102 4482 5105 4518
rect 5110 4492 5113 4528
rect 5126 4512 5129 4558
rect 5138 4548 5142 4551
rect 5142 4542 5145 4548
rect 5158 4542 5161 4558
rect 5182 4542 5185 4548
rect 5190 4542 5193 4558
rect 5170 4538 5174 4541
rect 5190 4532 5193 4538
rect 5162 4528 5166 4531
rect 5134 4492 5137 4518
rect 5166 4512 5169 4518
rect 5126 4472 5129 4488
rect 5198 4482 5201 4518
rect 5206 4492 5209 4548
rect 5214 4522 5217 4528
rect 5254 4522 5257 4548
rect 5262 4542 5265 4668
rect 5146 4478 5150 4481
rect 5278 4472 5281 4528
rect 5130 4468 5137 4471
rect 5102 4452 5105 4468
rect 5118 4462 5121 4468
rect 5134 4451 5137 4468
rect 5150 4468 5158 4471
rect 5186 4468 5190 4471
rect 5150 4462 5153 4468
rect 5254 4462 5257 4468
rect 5162 4458 5166 4461
rect 5186 4458 5190 4461
rect 5126 4448 5137 4451
rect 5230 4452 5233 4458
rect 5102 4441 5105 4448
rect 5102 4438 5113 4441
rect 5110 4352 5113 4438
rect 5110 4342 5113 4348
rect 5118 4292 5121 4348
rect 5126 4272 5129 4448
rect 5202 4418 5206 4421
rect 5126 4262 5129 4268
rect 5134 4262 5137 4418
rect 5142 4301 5145 4358
rect 5174 4352 5177 4358
rect 5190 4321 5193 4348
rect 5198 4332 5201 4338
rect 5182 4318 5193 4321
rect 5174 4312 5177 4318
rect 5142 4298 5153 4301
rect 5150 4292 5153 4298
rect 5142 4272 5145 4278
rect 5150 4262 5153 4288
rect 5106 4258 5110 4261
rect 5110 4192 5113 4218
rect 5110 4162 5113 4178
rect 5110 4072 5113 4128
rect 5078 4018 5089 4021
rect 4974 3968 4985 3971
rect 4890 3948 4894 3951
rect 4910 3942 4913 3948
rect 4846 3921 4849 3928
rect 4846 3918 4857 3921
rect 4854 3872 4857 3918
rect 4894 3912 4897 3938
rect 4918 3932 4921 3940
rect 4958 3932 4961 3938
rect 4926 3918 4934 3921
rect 4894 3882 4897 3888
rect 4926 3881 4929 3918
rect 4936 3903 4938 3907
rect 4942 3903 4945 3907
rect 4949 3903 4952 3907
rect 4926 3878 4934 3881
rect 4750 3862 4753 3868
rect 4750 3832 4753 3848
rect 4766 3752 4769 3868
rect 4786 3859 4790 3861
rect 4782 3858 4790 3859
rect 4846 3852 4849 3858
rect 4854 3841 4857 3868
rect 4862 3862 4865 3868
rect 4886 3852 4889 3878
rect 4918 3872 4921 3878
rect 4898 3858 4902 3861
rect 4874 3848 4878 3851
rect 4846 3838 4857 3841
rect 4822 3792 4825 3808
rect 4786 3788 4790 3791
rect 4822 3772 4825 3788
rect 4798 3762 4801 3768
rect 4838 3752 4841 3758
rect 4782 3748 4790 3751
rect 4750 3742 4753 3748
rect 4766 3672 4769 3748
rect 4674 3488 4678 3491
rect 4714 3488 4718 3491
rect 4714 3468 4718 3471
rect 4654 3462 4657 3468
rect 4662 3432 4665 3468
rect 4726 3462 4729 3518
rect 4698 3458 4702 3461
rect 4678 3431 4681 3448
rect 4686 3442 4689 3448
rect 4678 3428 4689 3431
rect 4686 3392 4689 3428
rect 4654 3352 4657 3368
rect 4666 3358 4670 3361
rect 4702 3352 4705 3418
rect 4734 3382 4737 3538
rect 4742 3502 4745 3548
rect 4718 3352 4721 3358
rect 4734 3352 4737 3378
rect 4758 3372 4761 3548
rect 4766 3482 4769 3668
rect 4774 3652 4777 3658
rect 4782 3612 4785 3748
rect 4838 3742 4841 3748
rect 4846 3742 4849 3838
rect 4862 3822 4865 3828
rect 4910 3812 4913 3858
rect 4854 3742 4857 3788
rect 4910 3752 4913 3768
rect 4918 3752 4921 3868
rect 4958 3802 4961 3868
rect 4942 3762 4945 3768
rect 4926 3752 4929 3758
rect 4862 3742 4865 3748
rect 4902 3742 4905 3748
rect 4790 3722 4793 3738
rect 4846 3732 4849 3738
rect 4918 3732 4921 3738
rect 4878 3728 4886 3731
rect 4862 3692 4865 3728
rect 4878 3722 4881 3728
rect 4814 3642 4817 3678
rect 4838 3672 4841 3688
rect 4878 3662 4881 3668
rect 4834 3658 4838 3661
rect 4894 3661 4897 3718
rect 4936 3703 4938 3707
rect 4942 3703 4945 3707
rect 4949 3703 4952 3707
rect 4890 3658 4897 3661
rect 4958 3662 4961 3668
rect 4790 3542 4793 3548
rect 4814 3542 4817 3618
rect 4766 3472 4769 3478
rect 4814 3472 4817 3518
rect 4846 3512 4849 3658
rect 4798 3462 4801 3468
rect 4846 3462 4849 3468
rect 4770 3458 4774 3461
rect 4766 3392 4769 3448
rect 4758 3352 4761 3368
rect 4746 3348 4750 3351
rect 4802 3348 4806 3351
rect 4638 3272 4641 3338
rect 4646 3312 4649 3338
rect 4594 3248 4598 3251
rect 4602 3238 4606 3241
rect 4494 3162 4497 3168
rect 4514 3148 4518 3151
rect 4526 3142 4529 3198
rect 4586 3178 4590 3181
rect 4550 3172 4553 3178
rect 4538 3168 4542 3171
rect 4558 3162 4561 3168
rect 4534 3152 4537 3158
rect 4578 3148 4582 3151
rect 4590 3142 4593 3148
rect 4334 3122 4337 3138
rect 4342 3101 4345 3118
rect 4334 3098 4345 3101
rect 4310 3062 4313 3068
rect 4262 3052 4265 3058
rect 4290 3048 4294 3051
rect 4310 3032 4313 3038
rect 4318 2992 4321 3068
rect 4278 2932 4281 2948
rect 4302 2912 4305 2938
rect 4318 2922 4321 2928
rect 4294 2862 4297 2878
rect 4318 2862 4321 2898
rect 4326 2872 4329 3028
rect 4334 2971 4337 3098
rect 4350 3082 4353 3138
rect 4366 3132 4369 3138
rect 4406 3132 4409 3138
rect 4470 3132 4473 3138
rect 4518 3132 4521 3138
rect 4566 3132 4569 3138
rect 4386 3128 4390 3131
rect 4398 3122 4401 3128
rect 4422 3122 4425 3128
rect 4350 3042 4353 3059
rect 4334 2968 4345 2971
rect 4342 2962 4345 2968
rect 4334 2952 4337 2958
rect 4358 2952 4361 2958
rect 4366 2942 4369 3118
rect 4478 3112 4481 3118
rect 4438 3062 4441 3088
rect 4494 3072 4497 3088
rect 4482 3058 4486 3061
rect 4502 3052 4505 3098
rect 4518 3072 4521 3108
rect 4526 3072 4529 3078
rect 4530 3068 4537 3071
rect 4458 3048 4462 3051
rect 4414 3032 4417 3048
rect 4418 3028 4422 3031
rect 4374 2962 4377 2968
rect 4334 2892 4337 2928
rect 4334 2872 4337 2878
rect 4326 2862 4329 2868
rect 4286 2858 4294 2861
rect 4314 2858 4318 2861
rect 4278 2752 4281 2818
rect 4230 2732 4233 2738
rect 4174 2642 4177 2658
rect 4158 2562 4161 2628
rect 4182 2562 4185 2588
rect 4130 2548 4134 2551
rect 4162 2548 4166 2551
rect 4174 2542 4177 2558
rect 4190 2552 4193 2648
rect 4198 2552 4201 2658
rect 4206 2612 4209 2658
rect 4230 2592 4233 2618
rect 4238 2572 4241 2718
rect 4246 2662 4249 2738
rect 4254 2582 4257 2748
rect 4262 2722 4265 2738
rect 4270 2712 4273 2738
rect 4278 2702 4281 2748
rect 4286 2732 4289 2858
rect 4334 2851 4337 2858
rect 4310 2848 4337 2851
rect 4310 2842 4313 2848
rect 4350 2812 4353 2938
rect 4374 2922 4377 2928
rect 4334 2762 4337 2768
rect 4298 2758 4302 2761
rect 4314 2748 4318 2751
rect 4310 2732 4313 2738
rect 4326 2722 4329 2738
rect 4278 2682 4281 2688
rect 4262 2662 4265 2668
rect 4326 2662 4329 2698
rect 4334 2662 4337 2738
rect 4374 2732 4377 2748
rect 4382 2742 4385 3018
rect 4390 2952 4393 3008
rect 4424 3003 4426 3007
rect 4430 3003 4433 3007
rect 4437 3003 4440 3007
rect 4418 2958 4425 2961
rect 4382 2682 4385 2718
rect 4390 2682 4393 2948
rect 4398 2942 4401 2958
rect 4422 2952 4425 2958
rect 4406 2932 4409 2938
rect 4414 2932 4417 2948
rect 4430 2922 4433 2958
rect 4414 2872 4417 2908
rect 4446 2892 4449 2928
rect 4402 2858 4406 2861
rect 4414 2752 4417 2868
rect 4424 2803 4426 2807
rect 4430 2803 4433 2807
rect 4437 2803 4440 2807
rect 4414 2742 4417 2748
rect 4378 2668 4382 2671
rect 4342 2662 4345 2668
rect 4398 2662 4401 2688
rect 4266 2658 4273 2661
rect 4306 2658 4310 2661
rect 4354 2658 4358 2661
rect 4262 2592 4265 2648
rect 4270 2582 4273 2658
rect 4338 2648 4342 2651
rect 4306 2628 4310 2631
rect 4318 2602 4321 2628
rect 4310 2552 4313 2578
rect 4318 2552 4321 2598
rect 4346 2578 4350 2581
rect 4382 2562 4385 2578
rect 4146 2538 4150 2541
rect 4130 2528 4134 2531
rect 4154 2518 4158 2521
rect 4142 2492 4145 2498
rect 4122 2478 4126 2481
rect 4102 2462 4105 2478
rect 4126 2462 4129 2468
rect 4090 2458 4094 2461
rect 4058 2448 4062 2451
rect 4066 2428 4070 2431
rect 3990 2362 3993 2418
rect 4022 2372 4025 2418
rect 3974 2342 3977 2348
rect 3982 2342 3985 2348
rect 3990 2331 3993 2348
rect 3998 2342 4001 2348
rect 3990 2328 4001 2331
rect 3974 2272 3977 2298
rect 3982 2272 3985 2308
rect 3946 2248 3950 2251
rect 3966 2201 3969 2258
rect 3966 2198 3974 2201
rect 3970 2188 3974 2191
rect 3926 2152 3929 2178
rect 3950 2162 3953 2168
rect 3890 2148 3894 2151
rect 3914 2148 3918 2151
rect 3882 2138 3886 2141
rect 3886 2092 3889 2108
rect 3920 2103 3922 2107
rect 3926 2103 3929 2107
rect 3933 2103 3936 2107
rect 3910 2072 3913 2098
rect 3846 2042 3849 2048
rect 3822 1952 3825 2028
rect 3870 2022 3873 2058
rect 3878 2042 3881 2068
rect 3902 2062 3905 2068
rect 3902 1952 3905 1968
rect 3798 1872 3801 1918
rect 3806 1912 3809 1948
rect 3910 1942 3913 2068
rect 3950 1982 3953 2148
rect 3878 1932 3881 1938
rect 3866 1928 3870 1931
rect 3858 1918 3862 1921
rect 3862 1892 3865 1908
rect 3810 1868 3814 1871
rect 3822 1868 3830 1871
rect 3790 1852 3793 1858
rect 3770 1848 3774 1851
rect 3766 1652 3769 1848
rect 3798 1682 3801 1868
rect 3806 1852 3809 1858
rect 3822 1692 3825 1868
rect 3830 1852 3833 1858
rect 3830 1812 3833 1848
rect 3838 1762 3841 1868
rect 3870 1862 3873 1918
rect 3846 1842 3849 1858
rect 3878 1852 3881 1928
rect 3886 1872 3889 1918
rect 3920 1903 3922 1907
rect 3926 1903 3929 1907
rect 3933 1903 3936 1907
rect 3942 1892 3945 1908
rect 3950 1882 3953 1898
rect 3958 1872 3961 2168
rect 3982 2152 3985 2258
rect 3990 2252 3993 2258
rect 3998 2252 4001 2328
rect 4006 2242 4009 2318
rect 4014 2281 4017 2358
rect 4038 2352 4041 2358
rect 4046 2352 4049 2418
rect 4078 2392 4081 2458
rect 4054 2382 4057 2388
rect 4078 2352 4081 2388
rect 4094 2362 4097 2428
rect 4102 2362 4105 2418
rect 4110 2392 4113 2458
rect 4102 2341 4105 2358
rect 4118 2352 4121 2418
rect 4134 2392 4137 2438
rect 4166 2402 4169 2538
rect 4118 2342 4121 2348
rect 4102 2338 4110 2341
rect 4022 2312 4025 2328
rect 4014 2278 4022 2281
rect 4022 2262 4025 2278
rect 4014 2242 4017 2258
rect 3990 2212 3993 2218
rect 3998 2192 4001 2208
rect 4014 2152 4017 2198
rect 4022 2152 4025 2248
rect 4006 2148 4014 2151
rect 3966 2142 3969 2148
rect 3978 2138 3982 2141
rect 3966 2102 3969 2138
rect 4006 2122 4009 2148
rect 4014 2092 4017 2118
rect 4022 2062 4025 2148
rect 4030 2122 4033 2338
rect 4038 2252 4041 2258
rect 4054 2192 4057 2318
rect 4070 2292 4073 2328
rect 4078 2322 4081 2338
rect 4070 2282 4073 2288
rect 4078 2272 4081 2288
rect 4082 2258 4086 2261
rect 4046 2142 4049 2148
rect 4058 2138 4062 2141
rect 4058 2078 4062 2081
rect 4030 2062 4033 2078
rect 4042 2068 4046 2071
rect 4086 2062 4089 2188
rect 4002 2058 4006 2061
rect 4046 2052 4049 2058
rect 3982 2032 3985 2038
rect 3982 1962 3985 1978
rect 3998 1962 4001 2008
rect 3998 1952 4001 1958
rect 4014 1942 4017 1958
rect 3966 1912 3969 1918
rect 3982 1882 3985 1918
rect 4006 1892 4009 1928
rect 3966 1872 3969 1878
rect 3926 1862 3929 1868
rect 3914 1858 3918 1861
rect 3870 1842 3873 1848
rect 3862 1752 3865 1828
rect 3878 1752 3881 1798
rect 3910 1792 3913 1818
rect 3886 1758 3894 1761
rect 3834 1748 3838 1751
rect 3846 1748 3854 1751
rect 3834 1738 3838 1741
rect 3830 1662 3833 1668
rect 3734 1552 3737 1558
rect 3674 1538 3678 1541
rect 3686 1532 3689 1548
rect 3702 1542 3705 1548
rect 3722 1538 3726 1541
rect 3730 1538 3737 1541
rect 3686 1492 3689 1528
rect 3630 1462 3633 1468
rect 3638 1462 3641 1478
rect 3622 1442 3625 1448
rect 3594 1358 3598 1361
rect 3630 1352 3633 1458
rect 3638 1352 3641 1358
rect 3646 1352 3649 1468
rect 3654 1462 3657 1468
rect 3662 1452 3665 1478
rect 3678 1452 3681 1468
rect 3686 1392 3689 1428
rect 3654 1352 3657 1358
rect 3610 1348 3614 1351
rect 3694 1351 3697 1518
rect 3718 1461 3721 1518
rect 3718 1458 3726 1461
rect 3690 1348 3697 1351
rect 3734 1352 3737 1538
rect 3750 1482 3753 1528
rect 3782 1472 3785 1578
rect 3830 1572 3833 1648
rect 3846 1582 3849 1748
rect 3870 1742 3873 1748
rect 3854 1661 3857 1678
rect 3870 1662 3873 1698
rect 3854 1658 3862 1661
rect 3854 1592 3857 1628
rect 3838 1552 3841 1558
rect 3794 1548 3798 1551
rect 3846 1542 3849 1548
rect 3822 1532 3825 1538
rect 3854 1492 3857 1568
rect 3862 1562 3865 1658
rect 3886 1572 3889 1758
rect 3898 1748 3902 1751
rect 3918 1742 3921 1748
rect 3934 1742 3937 1868
rect 4014 1862 4017 1868
rect 3954 1858 3958 1861
rect 3986 1858 3990 1861
rect 4022 1852 4025 1858
rect 3986 1848 3990 1851
rect 3974 1752 3977 1778
rect 3990 1772 3993 1818
rect 4006 1792 4009 1818
rect 3990 1752 3993 1768
rect 4006 1762 4009 1768
rect 3946 1748 3950 1751
rect 3982 1742 3985 1748
rect 4030 1742 4033 2028
rect 4038 1862 4041 1978
rect 4062 1952 4065 2058
rect 4078 1962 4081 1988
rect 4086 1982 4089 2058
rect 4094 1992 4097 2318
rect 4102 2202 4105 2318
rect 4126 2161 4129 2358
rect 4150 2352 4153 2388
rect 4166 2382 4169 2388
rect 4182 2352 4185 2528
rect 4190 2462 4193 2548
rect 4198 2502 4201 2548
rect 4278 2532 4281 2548
rect 4346 2538 4350 2541
rect 4294 2532 4297 2538
rect 4330 2528 4334 2531
rect 4342 2528 4350 2531
rect 4190 2362 4193 2368
rect 4178 2348 4182 2351
rect 4198 2332 4201 2468
rect 4206 2462 4209 2518
rect 4238 2491 4241 2528
rect 4238 2488 4246 2491
rect 4250 2468 4254 2471
rect 4254 2452 4257 2458
rect 4262 2432 4265 2518
rect 4326 2502 4329 2518
rect 4326 2472 4329 2478
rect 4282 2468 4286 2471
rect 4294 2462 4297 2468
rect 4318 2462 4321 2468
rect 4282 2458 4286 2461
rect 4310 2452 4313 2458
rect 4298 2448 4302 2451
rect 4262 2412 4265 2418
rect 4294 2382 4297 2388
rect 4134 2282 4137 2318
rect 4134 2242 4137 2248
rect 4126 2158 4137 2161
rect 4122 2148 4126 2151
rect 4102 2062 4105 2078
rect 4134 2062 4137 2158
rect 4142 2122 4145 2268
rect 4150 2262 4153 2268
rect 4190 2262 4193 2318
rect 4206 2272 4209 2368
rect 4254 2351 4257 2378
rect 4222 2332 4225 2348
rect 4290 2348 4294 2351
rect 4286 2332 4289 2338
rect 4226 2288 4230 2291
rect 4250 2288 4254 2291
rect 4222 2278 4230 2281
rect 4162 2258 4166 2261
rect 4174 2242 4177 2248
rect 4174 2172 4177 2238
rect 4198 2212 4201 2268
rect 4206 2152 4209 2258
rect 4222 2152 4225 2278
rect 4238 2272 4241 2278
rect 4262 2272 4265 2298
rect 4254 2252 4257 2258
rect 4262 2212 4265 2268
rect 4270 2262 4273 2318
rect 4274 2258 4278 2261
rect 4286 2242 4289 2248
rect 4302 2192 4305 2448
rect 4310 2402 4313 2448
rect 4314 2358 4318 2361
rect 4334 2352 4337 2528
rect 4342 2492 4345 2528
rect 4382 2522 4385 2528
rect 4358 2482 4361 2488
rect 4354 2468 4358 2471
rect 4358 2442 4361 2458
rect 4342 2392 4345 2438
rect 4310 2272 4313 2348
rect 4318 2272 4321 2278
rect 4310 2262 4313 2268
rect 4334 2262 4337 2348
rect 4342 2302 4345 2338
rect 4350 2282 4353 2378
rect 4366 2362 4369 2498
rect 4374 2462 4377 2488
rect 4382 2472 4385 2478
rect 4390 2452 4393 2648
rect 4398 2552 4401 2558
rect 4374 2352 4377 2438
rect 4398 2422 4401 2538
rect 4406 2462 4409 2678
rect 4414 2652 4417 2718
rect 4438 2692 4441 2748
rect 4446 2722 4449 2728
rect 4454 2671 4457 2988
rect 4470 2982 4473 3048
rect 4510 3032 4513 3038
rect 4486 2972 4489 3018
rect 4462 2822 4465 2918
rect 4470 2791 4473 2968
rect 4478 2952 4481 2958
rect 4486 2932 4489 2958
rect 4482 2918 4486 2921
rect 4494 2882 4497 3028
rect 4518 3012 4521 3068
rect 4502 2942 4505 2948
rect 4510 2942 4513 2958
rect 4518 2942 4521 2948
rect 4526 2942 4529 2948
rect 4518 2892 4521 2928
rect 4534 2922 4537 3068
rect 4582 3012 4585 3138
rect 4590 3072 4593 3138
rect 4598 3072 4601 3198
rect 4638 3152 4641 3258
rect 4646 3232 4649 3308
rect 4654 3302 4657 3348
rect 4686 3332 4689 3348
rect 4722 3338 4726 3341
rect 4714 3328 4718 3331
rect 4738 3328 4742 3331
rect 4662 3252 4665 3258
rect 4710 3192 4713 3308
rect 4730 3259 4734 3262
rect 4782 3232 4785 3348
rect 4802 3338 4806 3341
rect 4814 3332 4817 3418
rect 4830 3352 4833 3408
rect 4802 3328 4806 3331
rect 4826 3328 4830 3331
rect 4842 3328 4846 3331
rect 4790 3292 4793 3298
rect 4794 3268 4798 3271
rect 4814 3252 4817 3298
rect 4830 3272 4833 3278
rect 4842 3258 4846 3261
rect 4854 3252 4857 3658
rect 4906 3648 4910 3651
rect 4886 3622 4889 3628
rect 4926 3622 4929 3628
rect 4866 3548 4870 3551
rect 4870 3452 4873 3458
rect 4894 3441 4897 3538
rect 4910 3522 4913 3558
rect 4926 3552 4929 3618
rect 4930 3538 4934 3541
rect 4910 3462 4913 3508
rect 4894 3438 4905 3441
rect 4878 3352 4881 3368
rect 4870 3342 4873 3348
rect 4886 3341 4889 3388
rect 4902 3372 4905 3438
rect 4910 3402 4913 3458
rect 4878 3338 4889 3341
rect 4866 3318 4870 3321
rect 4878 3272 4881 3338
rect 4886 3322 4889 3328
rect 4874 3268 4878 3271
rect 4894 3271 4897 3358
rect 4890 3268 4897 3271
rect 4902 3272 4905 3278
rect 4918 3272 4921 3538
rect 4946 3528 4950 3531
rect 4936 3503 4938 3507
rect 4942 3503 4945 3507
rect 4949 3503 4952 3507
rect 4926 3482 4929 3488
rect 4950 3462 4953 3468
rect 4942 3362 4945 3418
rect 4934 3322 4937 3348
rect 4950 3332 4953 3458
rect 4966 3422 4969 3818
rect 4974 3802 4977 3968
rect 4998 3962 5001 3968
rect 5014 3962 5017 3968
rect 4986 3958 4990 3961
rect 4986 3948 4990 3951
rect 4998 3942 5001 3948
rect 4990 3932 4993 3938
rect 4990 3872 4993 3888
rect 4998 3862 5001 3898
rect 4982 3852 4985 3858
rect 4998 3822 5001 3828
rect 4990 3752 4993 3778
rect 4998 3772 5001 3778
rect 4982 3742 4985 3748
rect 4974 3732 4977 3738
rect 4974 3552 4977 3718
rect 4990 3692 4993 3738
rect 4990 3652 4993 3659
rect 4982 3552 4985 3608
rect 5006 3592 5009 3948
rect 5014 3852 5017 3948
rect 5050 3947 5054 3950
rect 5038 3882 5041 3888
rect 5026 3858 5030 3861
rect 5070 3842 5073 3948
rect 5078 3942 5081 4018
rect 5094 4012 5097 4058
rect 5110 4002 5113 4068
rect 5106 3968 5110 3971
rect 5118 3962 5121 4218
rect 5126 3992 5129 4258
rect 5134 4182 5137 4258
rect 5166 4252 5169 4268
rect 5174 4262 5177 4298
rect 5182 4281 5185 4318
rect 5238 4302 5241 4348
rect 5246 4342 5249 4348
rect 5190 4292 5193 4298
rect 5202 4288 5206 4291
rect 5182 4278 5193 4281
rect 5182 4262 5185 4268
rect 5166 4222 5169 4248
rect 5134 4092 5137 4178
rect 5150 4162 5153 4218
rect 5182 4152 5185 4228
rect 5190 4212 5193 4278
rect 5198 4272 5201 4278
rect 5246 4262 5249 4338
rect 5278 4322 5281 4328
rect 5250 4258 5257 4261
rect 5198 4192 5201 4198
rect 5150 4142 5153 4148
rect 5158 4142 5161 4148
rect 5174 4142 5177 4148
rect 5182 4092 5185 4148
rect 5190 4142 5193 4168
rect 5198 4122 5201 4148
rect 5166 4072 5169 4088
rect 5186 4078 5190 4081
rect 5162 4058 5166 4061
rect 5134 4032 5137 4048
rect 5150 4042 5153 4058
rect 5134 3952 5137 4028
rect 5190 4022 5193 4028
rect 5174 3962 5177 4018
rect 5146 3958 5150 3961
rect 5162 3948 5166 3951
rect 5182 3942 5185 4018
rect 5190 3992 5193 4008
rect 5190 3942 5193 3948
rect 5014 3722 5017 3798
rect 5054 3792 5057 3818
rect 5070 3791 5073 3838
rect 5110 3802 5113 3918
rect 5118 3902 5121 3918
rect 5142 3892 5145 3938
rect 5150 3932 5153 3938
rect 5118 3863 5121 3868
rect 5118 3858 5121 3859
rect 5134 3842 5137 3868
rect 5166 3862 5169 3938
rect 5174 3892 5177 3938
rect 5174 3872 5177 3878
rect 5154 3858 5158 3861
rect 5186 3858 5190 3861
rect 5166 3852 5169 3858
rect 5062 3788 5073 3791
rect 5054 3782 5057 3788
rect 5038 3732 5041 3748
rect 5062 3742 5065 3788
rect 5110 3782 5113 3788
rect 5078 3672 5081 3768
rect 5094 3762 5097 3778
rect 5110 3752 5113 3758
rect 5006 3562 5009 3568
rect 5022 3552 5025 3668
rect 5030 3642 5033 3658
rect 5038 3652 5041 3658
rect 5078 3652 5081 3658
rect 5054 3632 5057 3648
rect 4974 3532 4977 3538
rect 4974 3482 4977 3498
rect 4990 3492 4993 3538
rect 5010 3528 5014 3531
rect 5030 3492 5033 3548
rect 5038 3522 5041 3528
rect 5038 3472 5041 3478
rect 5010 3468 5014 3471
rect 4982 3452 4985 3468
rect 4990 3372 4993 3458
rect 5018 3448 5022 3451
rect 4966 3342 4969 3348
rect 4936 3303 4938 3307
rect 4942 3303 4945 3307
rect 4949 3303 4952 3307
rect 4966 3292 4969 3328
rect 4998 3312 5001 3318
rect 4946 3278 4950 3281
rect 4946 3268 4950 3271
rect 4966 3262 4969 3288
rect 4982 3282 4985 3308
rect 4862 3258 4870 3261
rect 4914 3258 4918 3261
rect 4938 3258 4942 3261
rect 4862 3252 4865 3258
rect 4850 3248 4854 3251
rect 4878 3251 4881 3258
rect 4874 3248 4881 3251
rect 4782 3192 4785 3228
rect 4806 3192 4809 3218
rect 4686 3182 4689 3188
rect 4730 3158 4734 3161
rect 4646 3132 4649 3148
rect 4622 3078 4638 3081
rect 4622 3062 4625 3078
rect 4646 3071 4649 3118
rect 4670 3092 4673 3138
rect 4694 3132 4697 3158
rect 4806 3152 4809 3178
rect 4818 3158 4822 3161
rect 4762 3148 4766 3151
rect 4726 3142 4729 3148
rect 4750 3142 4753 3148
rect 4830 3142 4833 3218
rect 4854 3162 4857 3168
rect 4894 3162 4897 3168
rect 4866 3148 4870 3151
rect 4882 3148 4886 3151
rect 4794 3138 4798 3141
rect 4662 3088 4670 3091
rect 4642 3068 4649 3071
rect 4602 3058 4606 3061
rect 4638 3052 4641 3058
rect 4654 3042 4657 3078
rect 4558 2952 4561 2998
rect 4582 2952 4585 3008
rect 4550 2932 4553 2938
rect 4558 2902 4561 2948
rect 4570 2938 4574 2941
rect 4562 2878 4566 2881
rect 4478 2852 4481 2858
rect 4486 2812 4489 2868
rect 4510 2842 4513 2878
rect 4526 2862 4529 2868
rect 4534 2862 4537 2878
rect 4578 2868 4582 2871
rect 4542 2862 4545 2868
rect 4590 2862 4593 2898
rect 4598 2882 4601 2888
rect 4578 2858 4582 2861
rect 4506 2818 4510 2821
rect 4614 2801 4617 3018
rect 4622 2932 4625 2948
rect 4662 2942 4665 3088
rect 4694 3082 4697 3128
rect 4734 3112 4737 3118
rect 4758 3102 4761 3138
rect 4678 2952 4681 2958
rect 4686 2932 4689 2988
rect 4694 2982 4697 3058
rect 4710 2992 4713 3098
rect 4742 3072 4745 3088
rect 4774 3068 4782 3071
rect 4722 3059 4726 3061
rect 4774 3062 4777 3068
rect 4722 3058 4729 3059
rect 4762 3058 4766 3061
rect 4762 3048 4766 3051
rect 4694 2952 4697 2978
rect 4694 2872 4697 2918
rect 4678 2862 4681 2868
rect 4642 2858 4646 2861
rect 4462 2788 4473 2791
rect 4606 2798 4617 2801
rect 4462 2692 4465 2788
rect 4558 2762 4561 2768
rect 4606 2762 4609 2798
rect 4574 2752 4577 2758
rect 4614 2752 4617 2788
rect 4482 2748 4486 2751
rect 4478 2732 4481 2738
rect 4526 2692 4529 2738
rect 4454 2668 4462 2671
rect 4466 2658 4470 2661
rect 4506 2658 4510 2661
rect 4454 2652 4457 2658
rect 4424 2603 4426 2607
rect 4430 2603 4433 2607
rect 4437 2603 4440 2607
rect 4430 2542 4433 2548
rect 4418 2468 4422 2471
rect 4406 2452 4409 2458
rect 4430 2422 4433 2538
rect 4446 2471 4449 2548
rect 4454 2542 4457 2578
rect 4462 2542 4465 2548
rect 4462 2472 4465 2478
rect 4470 2472 4473 2598
rect 4478 2542 4481 2658
rect 4486 2532 4489 2558
rect 4494 2482 4497 2618
rect 4518 2591 4521 2678
rect 4534 2662 4537 2668
rect 4514 2588 4521 2591
rect 4510 2492 4513 2498
rect 4478 2472 4481 2478
rect 4446 2470 4457 2471
rect 4446 2468 4454 2470
rect 4506 2468 4510 2471
rect 4442 2458 4446 2461
rect 4474 2458 4478 2461
rect 4370 2348 4374 2351
rect 4382 2342 4385 2418
rect 4424 2403 4426 2407
rect 4430 2403 4433 2407
rect 4437 2403 4440 2407
rect 4398 2362 4401 2398
rect 4406 2352 4409 2368
rect 4394 2318 4398 2321
rect 4358 2272 4361 2318
rect 4350 2252 4353 2259
rect 4314 2248 4318 2251
rect 4358 2222 4361 2268
rect 4406 2262 4409 2348
rect 4454 2342 4457 2428
rect 4462 2392 4465 2448
rect 4478 2352 4481 2418
rect 4494 2412 4497 2458
rect 4486 2352 4489 2358
rect 4502 2332 4505 2388
rect 4510 2362 4513 2368
rect 4518 2351 4521 2548
rect 4526 2381 4529 2648
rect 4542 2552 4545 2748
rect 4582 2742 4585 2748
rect 4590 2742 4593 2748
rect 4586 2738 4590 2741
rect 4550 2682 4553 2738
rect 4554 2668 4558 2671
rect 4566 2662 4569 2728
rect 4582 2672 4585 2688
rect 4550 2552 4553 2658
rect 4582 2591 4585 2668
rect 4598 2602 4601 2718
rect 4574 2588 4585 2591
rect 4566 2462 4569 2528
rect 4538 2388 4542 2391
rect 4574 2382 4577 2588
rect 4606 2572 4609 2578
rect 4614 2552 4617 2748
rect 4622 2742 4625 2768
rect 4646 2742 4649 2818
rect 4670 2762 4673 2778
rect 4654 2742 4657 2748
rect 4622 2692 4625 2738
rect 4630 2681 4633 2718
rect 4638 2712 4641 2728
rect 4622 2678 4633 2681
rect 4622 2662 4625 2678
rect 4670 2672 4673 2708
rect 4630 2662 4633 2668
rect 4622 2562 4625 2578
rect 4638 2552 4641 2588
rect 4646 2542 4649 2648
rect 4590 2502 4593 2538
rect 4614 2532 4617 2538
rect 4650 2518 4654 2521
rect 4590 2472 4593 2498
rect 4622 2472 4625 2518
rect 4638 2482 4641 2518
rect 4654 2462 4657 2468
rect 4626 2458 4630 2461
rect 4626 2448 4630 2451
rect 4526 2378 4537 2381
rect 4534 2352 4537 2378
rect 4510 2348 4521 2351
rect 4398 2242 4401 2248
rect 4414 2202 4417 2238
rect 4424 2203 4426 2207
rect 4430 2203 4433 2207
rect 4437 2203 4440 2207
rect 4234 2158 4238 2161
rect 4270 2152 4273 2188
rect 4294 2181 4297 2188
rect 4294 2178 4310 2181
rect 4438 2152 4441 2158
rect 4210 2148 4214 2151
rect 4290 2148 4294 2151
rect 4306 2148 4310 2151
rect 4146 2068 4150 2071
rect 4146 2058 4150 2061
rect 4126 2042 4129 2058
rect 4134 2002 4137 2058
rect 4158 2052 4161 2138
rect 4166 2072 4169 2078
rect 4174 2052 4177 2148
rect 4246 2142 4249 2148
rect 4186 2138 4190 2141
rect 4198 2112 4201 2118
rect 4210 2088 4214 2091
rect 4190 2072 4193 2078
rect 4202 2068 4206 2071
rect 4110 1962 4113 1968
rect 4142 1952 4145 2048
rect 4050 1948 4054 1951
rect 4046 1762 4049 1868
rect 4054 1862 4057 1938
rect 4062 1852 4065 1948
rect 4070 1942 4073 1948
rect 4094 1942 4097 1948
rect 4082 1938 4086 1941
rect 4106 1938 4110 1941
rect 4062 1772 4065 1848
rect 4062 1742 4065 1748
rect 3898 1728 3902 1731
rect 3902 1682 3905 1708
rect 3920 1703 3922 1707
rect 3926 1703 3929 1707
rect 3933 1703 3936 1707
rect 4030 1672 4033 1738
rect 4038 1672 4041 1698
rect 4070 1682 4073 1908
rect 4102 1892 4105 1918
rect 4102 1872 4105 1878
rect 4094 1862 4097 1868
rect 4110 1862 4113 1878
rect 4110 1701 4113 1768
rect 4118 1732 4121 1738
rect 4110 1698 4121 1701
rect 3950 1662 3953 1668
rect 4014 1662 4017 1668
rect 3938 1658 3942 1661
rect 4030 1652 4033 1658
rect 4002 1648 4006 1651
rect 4038 1641 4041 1668
rect 4094 1662 4097 1668
rect 4030 1638 4041 1641
rect 3910 1552 3913 1568
rect 3874 1548 3878 1551
rect 3966 1542 3969 1638
rect 3982 1612 3985 1618
rect 4030 1582 4033 1638
rect 4038 1592 4041 1598
rect 3982 1542 3985 1548
rect 3966 1532 3969 1538
rect 3898 1518 3902 1521
rect 3790 1462 3793 1478
rect 3818 1468 3825 1471
rect 3790 1452 3793 1458
rect 3810 1448 3814 1451
rect 3750 1362 3753 1368
rect 3766 1352 3769 1398
rect 3778 1358 3782 1361
rect 3790 1352 3793 1438
rect 3822 1412 3825 1468
rect 3838 1432 3841 1468
rect 3854 1462 3857 1478
rect 3866 1468 3870 1471
rect 3850 1448 3854 1451
rect 3582 1342 3585 1348
rect 3662 1342 3665 1348
rect 3474 1268 3478 1271
rect 3502 1262 3505 1278
rect 3542 1272 3545 1338
rect 3558 1332 3561 1338
rect 3510 1262 3513 1268
rect 3510 1222 3513 1258
rect 3400 1203 3402 1207
rect 3406 1203 3409 1207
rect 3413 1203 3416 1207
rect 3418 1158 3422 1161
rect 3374 1152 3377 1158
rect 3402 1148 3406 1151
rect 3310 1142 3313 1148
rect 3354 1138 3358 1141
rect 3310 1122 3313 1138
rect 3326 1122 3329 1128
rect 3334 1122 3337 1128
rect 3302 1112 3305 1118
rect 3302 1072 3305 1078
rect 3298 1058 3302 1061
rect 3318 1022 3321 1118
rect 3334 1102 3337 1118
rect 3334 1072 3337 1078
rect 3342 1062 3345 1118
rect 3366 1102 3369 1148
rect 3374 1142 3377 1148
rect 3366 1082 3369 1088
rect 3350 1062 3353 1068
rect 3390 1062 3393 1118
rect 3430 1082 3433 1188
rect 3526 1162 3529 1198
rect 3542 1192 3545 1268
rect 3554 1258 3558 1261
rect 3550 1192 3553 1228
rect 3566 1202 3569 1318
rect 3590 1302 3593 1328
rect 3606 1311 3609 1338
rect 3678 1332 3681 1338
rect 3598 1308 3609 1311
rect 3662 1318 3670 1321
rect 3598 1262 3601 1308
rect 3606 1292 3609 1298
rect 3622 1272 3625 1278
rect 3662 1262 3665 1318
rect 3686 1192 3689 1348
rect 3798 1342 3801 1408
rect 3822 1352 3825 1388
rect 3722 1328 3726 1331
rect 3474 1158 3478 1161
rect 3514 1158 3518 1161
rect 3538 1158 3542 1161
rect 3550 1152 3553 1178
rect 3566 1152 3569 1158
rect 3514 1148 3521 1151
rect 3438 1102 3441 1128
rect 3430 1063 3433 1068
rect 3326 1052 3329 1058
rect 3142 982 3145 998
rect 3094 952 3097 968
rect 3174 962 3177 968
rect 3074 948 3078 951
rect 3006 942 3009 948
rect 3146 938 3150 941
rect 2982 892 2985 918
rect 2986 858 2998 861
rect 2926 792 2929 858
rect 2878 772 2881 778
rect 2862 762 2865 768
rect 2790 748 2801 751
rect 2734 742 2737 747
rect 2786 738 2790 741
rect 2702 732 2705 738
rect 2626 668 2630 671
rect 2646 662 2649 668
rect 2662 662 2665 708
rect 2626 658 2630 661
rect 2646 602 2649 658
rect 2654 552 2657 658
rect 2662 572 2665 578
rect 2606 532 2609 538
rect 2622 532 2625 548
rect 2630 542 2633 548
rect 2646 532 2649 538
rect 2654 522 2657 548
rect 2670 532 2673 618
rect 2670 512 2673 528
rect 2678 482 2681 678
rect 2686 672 2689 698
rect 2726 672 2729 738
rect 2770 728 2774 731
rect 2710 662 2713 668
rect 2742 663 2745 668
rect 2698 658 2702 661
rect 2710 642 2713 648
rect 2778 548 2782 551
rect 2726 542 2729 547
rect 2670 472 2673 478
rect 2686 472 2689 508
rect 2718 472 2721 518
rect 2730 488 2734 491
rect 2706 468 2710 471
rect 2634 459 2638 462
rect 2686 462 2689 468
rect 2694 462 2697 468
rect 2718 462 2721 468
rect 2606 452 2609 458
rect 2742 452 2745 538
rect 2758 402 2761 548
rect 2770 538 2774 541
rect 2790 532 2793 568
rect 2798 502 2801 748
rect 2886 742 2889 758
rect 2902 752 2905 778
rect 2914 768 2918 771
rect 2934 762 2937 818
rect 2958 792 2961 848
rect 2974 842 2977 848
rect 2982 842 2985 848
rect 2922 748 2926 751
rect 2830 732 2833 738
rect 2838 682 2841 688
rect 2814 672 2817 678
rect 2814 662 2817 668
rect 2846 662 2849 668
rect 2822 652 2825 658
rect 2830 648 2838 651
rect 2806 552 2809 598
rect 2822 552 2825 558
rect 2806 542 2809 548
rect 2766 452 2769 458
rect 2782 452 2785 458
rect 2822 452 2825 488
rect 2706 378 2710 381
rect 2614 352 2617 378
rect 2702 352 2705 358
rect 2642 348 2646 351
rect 2614 342 2617 348
rect 2670 342 2673 348
rect 2634 338 2638 341
rect 2682 338 2686 341
rect 2598 332 2601 338
rect 2694 332 2697 338
rect 2658 328 2662 331
rect 2582 292 2585 328
rect 2630 322 2633 328
rect 2462 142 2465 208
rect 2254 92 2257 128
rect 2350 122 2353 128
rect 2286 112 2289 118
rect 2302 62 2305 108
rect 2366 92 2369 128
rect 2326 62 2329 68
rect 2374 62 2377 68
rect 2414 62 2417 78
rect 2438 62 2441 138
rect 2478 82 2481 228
rect 2518 192 2521 268
rect 2526 262 2529 268
rect 2590 262 2593 318
rect 2638 282 2641 288
rect 2646 282 2649 288
rect 2602 268 2606 271
rect 2630 262 2633 268
rect 2618 258 2622 261
rect 2598 252 2601 258
rect 2646 252 2649 278
rect 2678 272 2681 308
rect 2714 288 2718 291
rect 2714 268 2718 271
rect 2670 262 2673 268
rect 2698 258 2702 261
rect 2674 248 2678 251
rect 2682 248 2686 251
rect 2706 248 2710 251
rect 2542 142 2545 148
rect 2566 142 2569 148
rect 2522 138 2526 141
rect 2494 62 2497 98
rect 2614 82 2617 238
rect 2646 152 2649 218
rect 2726 172 2729 348
rect 2758 342 2761 348
rect 2766 342 2769 448
rect 2814 392 2817 438
rect 2774 252 2777 258
rect 2654 152 2657 158
rect 2634 148 2638 151
rect 2674 148 2678 151
rect 2514 78 2518 81
rect 2646 72 2649 148
rect 2742 142 2745 148
rect 2750 142 2753 168
rect 2782 152 2785 268
rect 2814 252 2817 358
rect 2830 302 2833 648
rect 2846 642 2849 648
rect 2854 572 2857 738
rect 2888 703 2890 707
rect 2894 703 2897 707
rect 2901 703 2904 707
rect 2890 688 2894 691
rect 2878 682 2881 688
rect 2870 672 2873 678
rect 2862 662 2865 668
rect 2910 662 2913 718
rect 2926 672 2929 728
rect 2934 712 2937 758
rect 2954 748 2958 751
rect 2974 732 2977 748
rect 2982 712 2985 748
rect 2990 741 2993 758
rect 2990 738 3001 741
rect 2990 722 2993 728
rect 2958 672 2961 678
rect 2898 658 2902 661
rect 2862 592 2865 648
rect 2898 568 2902 571
rect 2846 552 2849 568
rect 2882 548 2886 551
rect 2838 532 2841 538
rect 2854 532 2857 548
rect 2894 542 2897 558
rect 2838 462 2841 478
rect 2838 442 2841 448
rect 2846 372 2849 468
rect 2854 442 2857 448
rect 2862 431 2865 528
rect 2870 472 2873 528
rect 2888 503 2890 507
rect 2894 503 2897 507
rect 2901 503 2904 507
rect 2878 472 2881 498
rect 2870 462 2873 468
rect 2870 442 2873 448
rect 2854 428 2865 431
rect 2878 432 2881 468
rect 2910 462 2913 658
rect 2918 512 2921 668
rect 2966 662 2969 668
rect 2934 572 2937 618
rect 2898 458 2902 461
rect 2942 461 2945 658
rect 2954 648 2958 651
rect 2966 642 2969 648
rect 2982 642 2985 648
rect 2966 492 2969 618
rect 2998 612 3001 738
rect 3006 721 3009 938
rect 3086 892 3089 938
rect 3046 882 3049 888
rect 3070 872 3073 878
rect 3086 872 3089 888
rect 3094 882 3097 888
rect 3014 852 3017 858
rect 3022 852 3025 858
rect 3030 772 3033 858
rect 3038 842 3041 868
rect 3046 852 3049 858
rect 3062 792 3065 858
rect 3022 762 3025 768
rect 3042 748 3046 751
rect 3054 742 3057 748
rect 3042 738 3046 741
rect 3014 732 3017 738
rect 3006 718 3017 721
rect 3014 672 3017 718
rect 3014 621 3017 668
rect 3026 658 3030 661
rect 3006 618 3017 621
rect 3046 622 3049 738
rect 3062 702 3065 748
rect 3070 692 3073 868
rect 3102 862 3105 928
rect 3134 922 3137 928
rect 3134 862 3137 868
rect 3142 862 3145 888
rect 3114 858 3118 861
rect 3178 859 3182 861
rect 3174 858 3182 859
rect 3078 852 3081 858
rect 3118 842 3121 858
rect 3078 762 3081 808
rect 3078 732 3081 738
rect 3078 692 3081 698
rect 3006 552 3009 618
rect 3078 592 3081 648
rect 3034 558 3038 561
rect 3062 552 3065 578
rect 2982 542 2985 548
rect 3006 542 3009 548
rect 3038 542 3041 548
rect 3022 492 3025 538
rect 2978 478 3001 481
rect 2998 472 3001 478
rect 2978 468 2982 471
rect 2950 462 2953 468
rect 2942 458 2950 461
rect 2910 452 2913 458
rect 2846 312 2849 368
rect 2822 272 2825 278
rect 2838 272 2841 298
rect 2854 292 2857 428
rect 2870 342 2873 388
rect 2926 352 2929 418
rect 2942 362 2945 458
rect 2958 402 2961 468
rect 2990 462 2993 468
rect 3014 462 3017 488
rect 3054 462 3057 508
rect 3026 458 3030 461
rect 2990 392 2993 398
rect 3006 352 3009 448
rect 3030 442 3033 458
rect 3014 438 3022 441
rect 3054 441 3057 458
rect 3054 438 3065 441
rect 3014 392 3017 438
rect 3038 402 3041 418
rect 3062 392 3065 438
rect 3054 362 3057 378
rect 3038 352 3041 358
rect 3050 348 3054 351
rect 2902 342 2905 348
rect 2862 302 2865 328
rect 2846 272 2849 278
rect 2862 272 2865 298
rect 2830 232 2833 258
rect 2870 212 2873 338
rect 2982 322 2985 338
rect 2998 332 3001 338
rect 3006 332 3009 348
rect 2814 151 2817 158
rect 2830 142 2833 178
rect 2846 152 2849 168
rect 2854 142 2857 198
rect 2862 152 2865 158
rect 2878 142 2881 318
rect 2888 303 2890 307
rect 2894 303 2897 307
rect 2901 303 2904 307
rect 3022 302 3025 328
rect 3030 322 3033 338
rect 2926 282 2929 288
rect 2958 282 2961 298
rect 2886 252 2889 278
rect 2918 272 2921 278
rect 2906 258 2910 261
rect 2918 222 2921 268
rect 2942 262 2945 268
rect 2894 152 2897 198
rect 2942 152 2945 228
rect 2938 148 2942 151
rect 2706 138 2710 141
rect 2930 138 2934 141
rect 2662 132 2665 138
rect 2702 102 2705 138
rect 2722 128 2726 131
rect 2710 112 2713 118
rect 2742 82 2745 138
rect 2878 132 2881 138
rect 2886 121 2889 128
rect 2878 118 2889 121
rect 2782 92 2785 118
rect 2878 92 2881 118
rect 2888 103 2890 107
rect 2894 103 2897 107
rect 2901 103 2904 107
rect 2894 82 2897 88
rect 2910 82 2913 118
rect 2918 92 2921 128
rect 2926 102 2929 118
rect 2554 68 2558 71
rect 2738 68 2742 71
rect 2834 68 2838 71
rect 2502 62 2505 68
rect 2566 62 2569 68
rect 2574 62 2577 68
rect 2886 62 2889 78
rect 2958 72 2961 268
rect 2990 263 2993 278
rect 3022 262 3025 268
rect 3006 182 3009 218
rect 3006 152 3009 178
rect 3046 152 3049 338
rect 3062 302 3065 368
rect 3070 342 3073 538
rect 3078 512 3081 518
rect 3086 312 3089 788
rect 3094 762 3097 768
rect 3166 742 3169 747
rect 3182 742 3185 848
rect 3110 672 3113 678
rect 3142 672 3145 688
rect 3150 682 3153 718
rect 3114 668 3118 671
rect 3122 658 3126 661
rect 3138 658 3142 661
rect 3102 642 3105 648
rect 3094 472 3097 528
rect 3110 482 3113 658
rect 3166 652 3169 658
rect 3118 642 3121 648
rect 3182 632 3185 658
rect 3190 652 3193 668
rect 3198 662 3201 1018
rect 3310 952 3313 958
rect 3318 952 3321 958
rect 3282 948 3286 951
rect 3246 942 3249 947
rect 3282 938 3286 941
rect 3262 921 3265 938
rect 3262 918 3273 921
rect 3254 882 3257 888
rect 3270 872 3273 918
rect 3270 862 3273 868
rect 3310 862 3313 888
rect 3206 852 3209 858
rect 3206 792 3209 828
rect 3206 752 3209 788
rect 3230 752 3233 758
rect 3238 752 3241 798
rect 3270 752 3273 858
rect 3318 802 3321 948
rect 3358 942 3361 948
rect 3334 842 3337 938
rect 3370 888 3374 891
rect 3382 882 3385 1058
rect 3400 1003 3402 1007
rect 3406 1003 3409 1007
rect 3413 1003 3416 1007
rect 3446 992 3449 1138
rect 3454 1112 3457 1148
rect 3506 1138 3510 1141
rect 3498 1128 3502 1131
rect 3486 1092 3489 1118
rect 3494 1092 3497 1098
rect 3462 1002 3465 1028
rect 3462 952 3465 998
rect 3490 948 3494 951
rect 3438 932 3441 938
rect 3446 892 3449 948
rect 3454 941 3457 948
rect 3470 942 3473 948
rect 3454 938 3465 941
rect 3482 938 3486 941
rect 3462 882 3465 938
rect 3502 912 3505 1068
rect 3510 952 3513 988
rect 3518 942 3521 1148
rect 3542 1148 3550 1151
rect 3578 1148 3585 1151
rect 3534 1072 3537 1078
rect 3542 1062 3545 1148
rect 3558 1122 3561 1138
rect 3574 1092 3577 1138
rect 3530 1058 3534 1061
rect 3566 1061 3569 1088
rect 3566 1058 3574 1061
rect 3526 1052 3529 1058
rect 3554 1048 3558 1051
rect 3582 1002 3585 1148
rect 3598 1142 3601 1148
rect 3606 1142 3609 1168
rect 3634 1158 3638 1161
rect 3654 1142 3657 1188
rect 3606 1082 3609 1138
rect 3622 1122 3625 1128
rect 3658 1118 3662 1121
rect 3630 1092 3633 1118
rect 3626 1078 3630 1081
rect 3590 1062 3593 1078
rect 3622 1062 3625 1068
rect 3646 1062 3649 1078
rect 3662 1072 3665 1088
rect 3694 1081 3697 1308
rect 3702 1292 3705 1328
rect 3710 1252 3713 1268
rect 3722 1258 3726 1261
rect 3734 1242 3737 1338
rect 3742 1272 3745 1328
rect 3742 1252 3745 1258
rect 3714 1148 3718 1151
rect 3718 1082 3721 1088
rect 3694 1078 3705 1081
rect 3670 1072 3673 1078
rect 3690 1068 3694 1071
rect 3642 1058 3646 1061
rect 3634 1048 3638 1051
rect 3542 952 3545 978
rect 3590 952 3593 1018
rect 3622 952 3625 998
rect 3590 942 3593 948
rect 3622 942 3625 948
rect 3610 938 3614 941
rect 3514 928 3518 931
rect 3494 882 3497 888
rect 3362 868 3366 871
rect 3390 862 3393 868
rect 3406 862 3409 878
rect 3438 872 3441 878
rect 3454 872 3457 878
rect 3462 872 3465 878
rect 3482 868 3486 871
rect 3430 862 3433 868
rect 3494 862 3497 868
rect 3466 858 3470 861
rect 3350 852 3353 858
rect 3358 842 3361 858
rect 3400 803 3402 807
rect 3406 803 3409 807
rect 3413 803 3416 807
rect 3314 778 3318 781
rect 3218 748 3222 751
rect 3306 748 3310 751
rect 3246 742 3249 748
rect 3206 692 3209 718
rect 3134 552 3137 568
rect 3174 542 3177 628
rect 3182 592 3185 608
rect 3198 572 3201 658
rect 3230 552 3233 588
rect 3126 532 3129 538
rect 3174 502 3177 538
rect 3182 492 3185 548
rect 3246 541 3249 738
rect 3270 682 3273 748
rect 3334 742 3337 768
rect 3462 762 3465 778
rect 3442 758 3446 761
rect 3354 748 3358 751
rect 3382 751 3385 758
rect 3442 748 3446 751
rect 3478 742 3481 748
rect 3242 538 3249 541
rect 3210 528 3214 531
rect 3154 488 3158 491
rect 3094 372 3097 468
rect 3102 462 3105 468
rect 3110 462 3113 478
rect 3170 468 3174 471
rect 3054 292 3057 298
rect 3062 272 3065 298
rect 3070 262 3073 278
rect 3086 242 3089 248
rect 3094 222 3097 368
rect 3102 261 3105 308
rect 3110 282 3113 458
rect 3158 432 3161 468
rect 3170 458 3177 461
rect 3118 282 3121 428
rect 3134 352 3137 398
rect 3174 352 3177 458
rect 3182 451 3185 488
rect 3210 468 3214 471
rect 3210 458 3214 461
rect 3182 448 3190 451
rect 3206 352 3209 358
rect 3214 352 3217 368
rect 3222 352 3225 538
rect 3238 392 3241 538
rect 3226 348 3230 351
rect 3158 332 3161 338
rect 3118 272 3121 278
rect 3158 272 3161 278
rect 3174 262 3177 348
rect 3198 332 3201 338
rect 3214 292 3217 348
rect 3222 272 3225 278
rect 3102 258 3110 261
rect 3062 152 3065 198
rect 3070 152 3073 158
rect 3086 152 3089 158
rect 3102 152 3105 258
rect 3182 252 3185 258
rect 3206 252 3209 268
rect 3114 248 3118 251
rect 3122 238 3126 241
rect 3110 152 3113 158
rect 2986 148 2990 151
rect 3050 148 3054 151
rect 3098 148 3102 151
rect 3062 142 3065 148
rect 3114 138 3118 141
rect 3014 92 3017 108
rect 3110 92 3113 98
rect 3122 88 3126 91
rect 3134 82 3137 148
rect 3142 132 3145 218
rect 3158 152 3161 188
rect 3214 152 3217 208
rect 3222 192 3225 248
rect 3230 232 3233 258
rect 3222 172 3225 188
rect 3230 162 3233 218
rect 3158 142 3161 148
rect 3170 138 3174 141
rect 3142 102 3145 128
rect 3030 72 3033 78
rect 3054 62 3057 78
rect 3198 72 3201 78
rect 3182 63 3185 68
rect 2162 58 2166 61
rect 2482 58 2486 61
rect 2546 58 2550 61
rect 2650 58 2654 61
rect 2730 58 2734 61
rect 2826 58 2830 61
rect 2890 58 2894 61
rect 2962 58 2966 61
rect 3214 62 3217 148
rect 3238 142 3241 388
rect 3246 302 3249 468
rect 3254 462 3257 638
rect 3262 632 3265 658
rect 3278 512 3281 558
rect 3278 472 3281 508
rect 3286 482 3289 688
rect 3302 662 3305 698
rect 3302 602 3305 618
rect 3306 548 3310 551
rect 3294 542 3297 548
rect 3310 532 3313 548
rect 3302 462 3305 488
rect 3310 472 3313 478
rect 3318 472 3321 728
rect 3334 692 3337 738
rect 3422 722 3425 738
rect 3430 732 3433 738
rect 3390 672 3393 678
rect 3406 662 3409 718
rect 3486 692 3489 848
rect 3494 752 3497 758
rect 3502 752 3505 908
rect 3526 892 3529 918
rect 3514 848 3518 851
rect 3534 802 3537 928
rect 3550 892 3553 938
rect 3574 932 3577 938
rect 3638 921 3641 938
rect 3630 918 3641 921
rect 3542 872 3545 878
rect 3542 782 3545 858
rect 3558 812 3561 918
rect 3606 862 3609 918
rect 3630 872 3633 918
rect 3654 902 3657 1068
rect 3702 1062 3705 1078
rect 3714 1068 3718 1071
rect 3726 1062 3729 1188
rect 3750 1172 3753 1318
rect 3758 1292 3761 1338
rect 3790 1331 3793 1338
rect 3790 1328 3814 1331
rect 3806 1312 3809 1318
rect 3774 1288 3793 1291
rect 3774 1272 3777 1288
rect 3790 1281 3793 1288
rect 3806 1282 3809 1288
rect 3790 1278 3798 1281
rect 3758 1262 3761 1268
rect 3782 1262 3785 1278
rect 3814 1272 3817 1318
rect 3822 1272 3825 1308
rect 3838 1302 3841 1318
rect 3854 1312 3857 1318
rect 3830 1272 3833 1288
rect 3850 1268 3854 1271
rect 3766 1242 3769 1248
rect 3766 1192 3769 1228
rect 3782 1192 3785 1258
rect 3790 1232 3793 1268
rect 3814 1202 3817 1268
rect 3822 1262 3825 1268
rect 3862 1262 3865 1458
rect 3886 1442 3889 1468
rect 3894 1452 3897 1478
rect 3902 1292 3905 1518
rect 3920 1503 3922 1507
rect 3926 1503 3929 1507
rect 3933 1503 3936 1507
rect 3910 1472 3913 1478
rect 3966 1472 3969 1528
rect 4030 1502 4033 1578
rect 4050 1538 4054 1541
rect 4050 1488 4054 1491
rect 3958 1442 3961 1459
rect 3958 1392 3961 1428
rect 3910 1332 3913 1348
rect 3920 1303 3922 1307
rect 3926 1303 3929 1307
rect 3933 1303 3936 1307
rect 3958 1272 3961 1338
rect 3974 1312 3977 1488
rect 3986 1478 3990 1481
rect 4034 1468 4049 1471
rect 3842 1258 3846 1261
rect 3862 1252 3865 1258
rect 3878 1242 3881 1268
rect 3894 1232 3897 1258
rect 3918 1252 3921 1258
rect 3846 1192 3849 1228
rect 3926 1222 3929 1258
rect 3742 1112 3745 1138
rect 3758 1092 3761 1158
rect 3838 1152 3841 1158
rect 3910 1152 3913 1218
rect 3958 1172 3961 1268
rect 3974 1263 3977 1268
rect 3974 1258 3977 1259
rect 3778 1148 3782 1151
rect 3766 1141 3769 1148
rect 3766 1138 3774 1141
rect 3802 1118 3806 1121
rect 3806 1082 3809 1088
rect 3754 1078 3758 1081
rect 3674 1058 3678 1061
rect 3714 1058 3718 1061
rect 3686 992 3689 1058
rect 3742 1022 3745 1078
rect 3758 962 3761 1068
rect 3822 1062 3825 1118
rect 3894 1111 3897 1148
rect 3958 1142 3961 1168
rect 3970 1148 3974 1151
rect 3886 1108 3897 1111
rect 3854 1072 3857 1108
rect 3886 1072 3889 1108
rect 3920 1103 3922 1107
rect 3926 1103 3929 1107
rect 3933 1103 3936 1107
rect 3902 1072 3905 1078
rect 3770 1058 3774 1061
rect 3802 1058 3806 1061
rect 3782 1002 3785 1018
rect 3734 952 3737 958
rect 3666 948 3670 951
rect 3746 948 3750 951
rect 3730 938 3734 941
rect 3722 918 3726 921
rect 3670 892 3673 918
rect 3718 892 3721 898
rect 3750 882 3753 918
rect 3766 882 3769 998
rect 3774 952 3777 988
rect 3782 972 3785 988
rect 3782 962 3785 968
rect 3798 952 3801 958
rect 3822 951 3825 1038
rect 3830 992 3833 1008
rect 3854 972 3857 1068
rect 3870 1063 3873 1068
rect 3918 1062 3921 1068
rect 3958 1062 3961 1098
rect 3982 1092 3985 1468
rect 4034 1458 4038 1461
rect 4006 1372 4009 1438
rect 4046 1412 4049 1468
rect 4054 1442 4057 1448
rect 4062 1422 4065 1518
rect 4006 1352 4009 1368
rect 4014 1352 4017 1408
rect 4062 1352 4065 1418
rect 4070 1352 4073 1558
rect 4086 1552 4089 1638
rect 4098 1558 4102 1561
rect 4078 1472 4081 1548
rect 4086 1512 4089 1548
rect 4106 1538 4110 1541
rect 4118 1532 4121 1698
rect 4126 1592 4129 1938
rect 4142 1912 4145 1948
rect 4150 1892 4153 2028
rect 4162 1948 4166 1951
rect 4174 1902 4177 2048
rect 4198 1982 4201 2058
rect 4222 2032 4225 2138
rect 4238 2082 4241 2088
rect 4234 2068 4238 2071
rect 4230 2052 4233 2058
rect 4202 1968 4206 1971
rect 4190 1942 4193 1948
rect 4182 1882 4185 1898
rect 4214 1882 4217 1888
rect 4190 1872 4193 1878
rect 4150 1852 4153 1868
rect 4162 1858 4166 1861
rect 4166 1812 4169 1858
rect 4174 1842 4177 1868
rect 4198 1792 4201 1868
rect 4206 1862 4209 1878
rect 4214 1862 4217 1868
rect 4182 1752 4185 1758
rect 4214 1752 4217 1818
rect 4222 1761 4225 1998
rect 4230 1832 4233 1868
rect 4246 1862 4249 1868
rect 4254 1862 4257 2148
rect 4382 2142 4385 2148
rect 4286 2132 4289 2138
rect 4286 2072 4289 2108
rect 4262 1942 4265 1948
rect 4270 1942 4273 1947
rect 4286 1942 4289 2068
rect 4302 2063 4305 2088
rect 4302 2058 4305 2059
rect 4334 2052 4337 2078
rect 4342 1971 4345 2118
rect 4374 2112 4377 2138
rect 4382 2108 4390 2111
rect 4362 2088 4366 2091
rect 4350 2062 4353 2068
rect 4350 2042 4353 2048
rect 4358 2002 4361 2068
rect 4382 2062 4385 2108
rect 4446 2102 4449 2268
rect 4454 2192 4457 2248
rect 4462 2172 4465 2318
rect 4470 2272 4473 2278
rect 4486 2272 4489 2298
rect 4510 2292 4513 2348
rect 4526 2342 4529 2348
rect 4502 2272 4505 2278
rect 4478 2262 4481 2268
rect 4462 2132 4465 2138
rect 4470 2132 4473 2148
rect 4402 2068 4406 2071
rect 4366 2042 4369 2048
rect 4342 1968 4353 1971
rect 4302 1942 4305 1968
rect 4314 1958 4318 1961
rect 4342 1952 4345 1958
rect 4318 1942 4321 1948
rect 4350 1942 4353 1968
rect 4362 1948 4366 1951
rect 4390 1942 4393 2068
rect 4402 2058 4406 2061
rect 4446 2052 4449 2088
rect 4462 2072 4465 2088
rect 4478 2081 4481 2258
rect 4494 2162 4497 2258
rect 4526 2252 4529 2278
rect 4494 2082 4497 2158
rect 4502 2152 4505 2158
rect 4518 2152 4521 2218
rect 4526 2152 4529 2238
rect 4534 2141 4537 2348
rect 4542 2272 4545 2278
rect 4550 2272 4553 2318
rect 4558 2262 4561 2368
rect 4574 2352 4577 2378
rect 4582 2352 4585 2358
rect 4606 2342 4609 2448
rect 4654 2372 4657 2458
rect 4638 2352 4641 2358
rect 4662 2352 4665 2668
rect 4678 2662 4681 2858
rect 4694 2772 4697 2868
rect 4686 2762 4689 2768
rect 4702 2762 4705 2958
rect 4710 2792 4713 2918
rect 4710 2752 4713 2788
rect 4690 2748 4697 2751
rect 4694 2692 4697 2748
rect 4702 2738 4710 2741
rect 4686 2662 4689 2688
rect 4686 2602 4689 2658
rect 4702 2632 4705 2738
rect 4718 2672 4721 3048
rect 4774 3032 4777 3058
rect 4782 3002 4785 3058
rect 4794 3038 4798 3041
rect 4782 2952 4785 2998
rect 4822 2962 4825 3118
rect 4838 3112 4841 3148
rect 4890 3138 4894 3141
rect 4838 3102 4841 3108
rect 4854 3063 4857 3098
rect 4870 3092 4873 3128
rect 4870 3072 4873 3088
rect 4886 3042 4889 3048
rect 4870 2952 4873 2958
rect 4734 2942 4737 2948
rect 4758 2932 4761 2948
rect 4826 2938 4830 2941
rect 4838 2922 4841 2948
rect 4846 2942 4849 2948
rect 4886 2942 4889 2998
rect 4894 2952 4897 3108
rect 4902 3062 4905 3088
rect 4910 3072 4913 3108
rect 4918 3092 4921 3098
rect 4910 3052 4913 3068
rect 4902 3042 4905 3048
rect 4918 3042 4921 3048
rect 4926 3032 4929 3258
rect 4966 3232 4969 3258
rect 4990 3212 4993 3218
rect 4938 3148 4942 3151
rect 4974 3132 4977 3138
rect 4936 3103 4938 3107
rect 4942 3103 4945 3107
rect 4949 3103 4952 3107
rect 4966 3072 4969 3098
rect 4990 3092 4993 3188
rect 5006 3152 5009 3378
rect 5014 3152 5017 3408
rect 5030 3402 5033 3458
rect 5038 3452 5041 3458
rect 5038 3282 5041 3448
rect 5030 3192 5033 3198
rect 5038 3152 5041 3208
rect 5046 3161 5049 3518
rect 5078 3482 5081 3648
rect 5094 3552 5097 3558
rect 5094 3472 5097 3538
rect 5086 3462 5089 3468
rect 5054 3332 5057 3348
rect 5062 3342 5065 3438
rect 5102 3382 5105 3688
rect 5110 3652 5113 3748
rect 5118 3742 5121 3768
rect 5126 3752 5129 3808
rect 5150 3792 5153 3848
rect 5158 3762 5161 3768
rect 5126 3732 5129 3738
rect 5134 3702 5137 3748
rect 5142 3722 5145 3738
rect 5150 3692 5153 3758
rect 5174 3752 5177 3858
rect 5162 3718 5166 3721
rect 5174 3702 5177 3748
rect 5182 3732 5185 3738
rect 5142 3672 5145 3678
rect 5130 3658 5134 3661
rect 5138 3648 5142 3651
rect 5114 3638 5118 3641
rect 5146 3638 5150 3641
rect 5118 3501 5121 3638
rect 5150 3592 5153 3618
rect 5158 3581 5161 3698
rect 5182 3662 5185 3668
rect 5166 3592 5169 3598
rect 5158 3578 5169 3581
rect 5134 3522 5137 3558
rect 5158 3552 5161 3558
rect 5110 3498 5121 3501
rect 5102 3352 5105 3368
rect 5062 3272 5065 3338
rect 5094 3321 5097 3348
rect 5086 3318 5097 3321
rect 5062 3202 5065 3258
rect 5046 3158 5054 3161
rect 4998 3072 5001 3148
rect 4934 3062 4937 3068
rect 4942 3062 4945 3068
rect 4882 2938 4886 2941
rect 4750 2872 4753 2878
rect 4738 2768 4742 2771
rect 4754 2758 4758 2761
rect 4766 2752 4769 2868
rect 4798 2862 4801 2878
rect 4846 2872 4849 2938
rect 4858 2928 4862 2931
rect 4806 2862 4809 2868
rect 4838 2862 4841 2868
rect 4854 2862 4857 2908
rect 4862 2872 4865 2878
rect 4778 2858 4782 2861
rect 4830 2852 4833 2858
rect 4794 2848 4798 2851
rect 4774 2832 4777 2838
rect 4794 2768 4798 2771
rect 4750 2748 4758 2751
rect 4786 2748 4790 2751
rect 4750 2741 4753 2748
rect 4738 2738 4753 2741
rect 4790 2732 4793 2738
rect 4770 2718 4774 2721
rect 4742 2692 4745 2708
rect 4670 2492 4673 2538
rect 4686 2481 4689 2598
rect 4702 2512 4705 2628
rect 4710 2622 4713 2658
rect 4718 2612 4721 2668
rect 4750 2662 4753 2718
rect 4758 2682 4761 2688
rect 4782 2672 4785 2688
rect 4806 2682 4809 2798
rect 4830 2662 4833 2788
rect 4854 2772 4857 2858
rect 4878 2852 4881 2898
rect 4890 2868 4894 2871
rect 4902 2862 4905 2978
rect 4910 2962 4913 2978
rect 4926 2958 4945 2961
rect 4926 2952 4929 2958
rect 4942 2952 4945 2958
rect 4934 2942 4937 2948
rect 4958 2942 4961 3028
rect 4966 3002 4969 3068
rect 4974 3052 4977 3058
rect 4998 3052 5001 3068
rect 4990 2982 4993 2988
rect 4966 2962 4969 2968
rect 4942 2922 4945 2938
rect 4982 2932 4985 2938
rect 4936 2903 4938 2907
rect 4942 2903 4945 2907
rect 4949 2903 4952 2907
rect 4942 2832 4945 2868
rect 4954 2858 4958 2861
rect 4974 2852 4977 2918
rect 4986 2888 4993 2891
rect 4990 2872 4993 2888
rect 4958 2842 4961 2848
rect 4854 2722 4857 2748
rect 4878 2742 4881 2778
rect 4918 2772 4921 2818
rect 4990 2772 4993 2868
rect 4926 2762 4929 2768
rect 4898 2758 4902 2761
rect 4906 2748 4910 2751
rect 4926 2742 4929 2748
rect 4918 2732 4921 2738
rect 4838 2672 4841 2678
rect 4862 2662 4865 2728
rect 4870 2672 4873 2708
rect 4894 2702 4897 2718
rect 4918 2712 4921 2728
rect 4958 2722 4961 2758
rect 4974 2752 4977 2768
rect 4966 2732 4969 2738
rect 4936 2703 4938 2707
rect 4942 2703 4945 2707
rect 4949 2703 4952 2707
rect 4898 2678 4902 2681
rect 4910 2672 4913 2688
rect 4998 2682 5001 3018
rect 5014 3012 5017 3148
rect 5070 3141 5073 3288
rect 5086 3222 5089 3318
rect 5102 3282 5105 3318
rect 5102 3192 5105 3248
rect 5110 3162 5113 3498
rect 5126 3452 5129 3468
rect 5142 3462 5145 3468
rect 5150 3462 5153 3548
rect 5158 3532 5161 3538
rect 5166 3471 5169 3578
rect 5190 3531 5193 3818
rect 5198 3542 5201 4108
rect 5206 3962 5209 4238
rect 5214 4142 5217 4148
rect 5222 4142 5225 4158
rect 5230 4152 5233 4188
rect 5222 3992 5225 4098
rect 5230 4042 5233 4058
rect 5206 3682 5209 3818
rect 5222 3752 5225 3838
rect 5238 3821 5241 4148
rect 5246 4132 5249 4138
rect 5254 4082 5257 4258
rect 5270 4192 5273 4259
rect 5262 4142 5265 4178
rect 5282 4158 5286 4161
rect 5254 3872 5257 4078
rect 5270 4072 5273 4148
rect 5274 3938 5278 3941
rect 5258 3858 5262 3861
rect 5230 3818 5241 3821
rect 5222 3732 5225 3738
rect 5222 3701 5225 3728
rect 5214 3698 5225 3701
rect 5206 3652 5209 3658
rect 5190 3528 5201 3531
rect 5186 3518 5190 3521
rect 5158 3468 5169 3471
rect 5178 3468 5182 3471
rect 5126 3352 5129 3438
rect 5118 3342 5121 3348
rect 5126 3342 5129 3348
rect 5126 3272 5129 3328
rect 5118 3262 5121 3268
rect 5118 3232 5121 3258
rect 5082 3158 5086 3161
rect 5094 3151 5097 3158
rect 5118 3152 5121 3218
rect 5126 3152 5129 3158
rect 5090 3148 5097 3151
rect 5070 3138 5078 3141
rect 5030 3072 5033 3138
rect 5038 3062 5041 3128
rect 5046 3082 5049 3138
rect 5078 3132 5081 3138
rect 5054 3122 5057 3128
rect 5078 3072 5081 3078
rect 5094 3031 5097 3108
rect 5086 3028 5097 3031
rect 5022 2882 5025 2998
rect 5086 2952 5089 3028
rect 5094 3012 5097 3018
rect 5102 3012 5105 3148
rect 5110 3132 5113 3138
rect 5118 3112 5121 3148
rect 5126 3072 5129 3078
rect 5094 2952 5097 2958
rect 5034 2948 5038 2951
rect 5046 2882 5049 2938
rect 5102 2892 5105 2998
rect 5110 2992 5113 3058
rect 5118 2892 5121 2948
rect 5078 2872 5081 2878
rect 5062 2862 5065 2868
rect 5014 2858 5022 2861
rect 5014 2792 5017 2858
rect 5038 2772 5041 2818
rect 5054 2792 5057 2808
rect 5042 2768 5049 2771
rect 5014 2752 5017 2758
rect 5038 2752 5041 2768
rect 4946 2668 4950 2671
rect 4770 2658 4774 2661
rect 4726 2652 4729 2658
rect 4834 2648 4838 2651
rect 4842 2648 4846 2651
rect 4710 2542 4713 2548
rect 4678 2478 4689 2481
rect 4678 2472 4681 2478
rect 4694 2472 4697 2478
rect 4710 2472 4713 2488
rect 4686 2462 4689 2468
rect 4718 2462 4721 2578
rect 4766 2562 4769 2608
rect 4790 2582 4793 2618
rect 4814 2591 4817 2638
rect 4862 2632 4865 2658
rect 4810 2588 4817 2591
rect 4806 2572 4809 2588
rect 4766 2552 4769 2558
rect 4790 2542 4793 2558
rect 4734 2502 4737 2538
rect 4782 2532 4785 2538
rect 4750 2522 4753 2528
rect 4782 2482 4785 2518
rect 4770 2478 4774 2481
rect 4790 2472 4793 2478
rect 4798 2472 4801 2548
rect 4814 2462 4817 2558
rect 4862 2552 4865 2618
rect 4870 2542 4873 2668
rect 4878 2662 4881 2668
rect 4910 2662 4913 2668
rect 4886 2562 4889 2618
rect 4902 2602 4905 2658
rect 4930 2648 4934 2651
rect 4942 2632 4945 2658
rect 5014 2572 5017 2748
rect 5022 2742 5025 2748
rect 5030 2732 5033 2738
rect 4902 2541 4905 2558
rect 4910 2552 4913 2558
rect 4918 2552 4921 2568
rect 4990 2552 4993 2558
rect 4902 2538 4913 2541
rect 4838 2502 4841 2538
rect 4838 2492 4841 2498
rect 4870 2492 4873 2538
rect 4886 2492 4889 2538
rect 4698 2458 4702 2461
rect 4686 2382 4689 2458
rect 4750 2452 4753 2458
rect 4734 2362 4737 2448
rect 4702 2342 4705 2348
rect 4710 2342 4713 2348
rect 4658 2338 4662 2341
rect 4546 2258 4550 2261
rect 4578 2258 4582 2261
rect 4566 2252 4569 2258
rect 4526 2138 4537 2141
rect 4526 2122 4529 2138
rect 4534 2122 4537 2128
rect 4478 2078 4486 2081
rect 4470 2072 4473 2078
rect 4510 2062 4513 2108
rect 4542 2072 4545 2158
rect 4550 2072 4553 2248
rect 4590 2222 4593 2258
rect 4578 2148 4582 2151
rect 4590 2102 4593 2218
rect 4598 2142 4601 2338
rect 4678 2332 4681 2338
rect 4670 2322 4673 2328
rect 4686 2322 4689 2328
rect 4718 2322 4721 2328
rect 4698 2318 4702 2321
rect 4610 2248 4614 2251
rect 4638 2161 4641 2318
rect 4686 2282 4689 2288
rect 4718 2262 4721 2268
rect 4726 2262 4729 2338
rect 4750 2282 4753 2338
rect 4758 2322 4761 2348
rect 4766 2322 4769 2458
rect 4790 2452 4793 2458
rect 4802 2448 4806 2451
rect 4782 2342 4785 2378
rect 4814 2362 4817 2368
rect 4822 2352 4825 2468
rect 4886 2382 4889 2488
rect 4894 2432 4897 2468
rect 4902 2452 4905 2518
rect 4910 2472 4913 2538
rect 4918 2442 4921 2548
rect 4926 2542 4929 2548
rect 4926 2512 4929 2528
rect 4938 2518 4942 2521
rect 4926 2472 4929 2508
rect 4936 2503 4938 2507
rect 4942 2503 4945 2507
rect 4949 2503 4952 2507
rect 4934 2472 4937 2478
rect 4938 2458 4942 2461
rect 4926 2452 4929 2458
rect 4958 2452 4961 2548
rect 4966 2522 4969 2538
rect 4974 2492 4977 2498
rect 4886 2352 4889 2378
rect 4766 2292 4769 2298
rect 4758 2272 4761 2288
rect 4774 2282 4777 2308
rect 4782 2282 4785 2318
rect 4798 2281 4801 2348
rect 4814 2292 4817 2328
rect 4830 2292 4833 2348
rect 4838 2322 4841 2338
rect 4902 2332 4905 2348
rect 4846 2312 4849 2318
rect 4838 2292 4841 2298
rect 4858 2288 4862 2291
rect 4822 2282 4825 2288
rect 4798 2278 4809 2281
rect 4730 2258 4734 2261
rect 4678 2252 4681 2258
rect 4634 2158 4641 2161
rect 4598 2132 4601 2138
rect 4614 2072 4617 2148
rect 4646 2142 4649 2148
rect 4654 2142 4657 2188
rect 4662 2162 4665 2168
rect 4670 2132 4673 2158
rect 4682 2148 4686 2151
rect 4678 2122 4681 2138
rect 4622 2082 4625 2118
rect 4630 2112 4633 2118
rect 4634 2068 4641 2071
rect 4566 2062 4569 2068
rect 4482 2058 4486 2061
rect 4522 2058 4526 2061
rect 4538 2058 4542 2061
rect 4490 2048 4494 2051
rect 4406 2042 4409 2048
rect 4424 2003 4426 2007
rect 4430 2003 4433 2007
rect 4437 2003 4440 2007
rect 4478 1982 4481 2018
rect 4286 1902 4289 1938
rect 4294 1882 4297 1888
rect 4282 1868 4286 1871
rect 4342 1862 4345 1898
rect 4390 1872 4393 1938
rect 4414 1902 4417 1938
rect 4430 1892 4433 1947
rect 4366 1862 4369 1868
rect 4414 1862 4417 1868
rect 4238 1832 4241 1858
rect 4254 1852 4257 1858
rect 4406 1852 4409 1858
rect 4222 1758 4230 1761
rect 4250 1758 4254 1761
rect 4138 1738 4142 1741
rect 4134 1692 4137 1708
rect 4166 1702 4169 1748
rect 4174 1682 4177 1748
rect 4198 1742 4201 1748
rect 4198 1722 4201 1728
rect 4206 1712 4209 1738
rect 4214 1692 4217 1748
rect 4238 1732 4241 1738
rect 4230 1692 4233 1718
rect 4222 1672 4225 1678
rect 4162 1668 4166 1671
rect 4194 1668 4198 1671
rect 4218 1668 4222 1671
rect 4178 1658 4182 1661
rect 4202 1658 4206 1661
rect 4158 1652 4161 1658
rect 4134 1542 4137 1608
rect 4190 1592 4193 1648
rect 4230 1602 4233 1658
rect 4238 1652 4241 1668
rect 4166 1562 4169 1588
rect 4174 1562 4177 1568
rect 4190 1552 4193 1578
rect 4222 1562 4225 1588
rect 4230 1562 4233 1568
rect 4246 1562 4249 1758
rect 4254 1682 4257 1688
rect 4262 1672 4265 1808
rect 4342 1792 4345 1838
rect 4278 1772 4281 1778
rect 4274 1748 4278 1751
rect 4278 1742 4281 1748
rect 4286 1742 4289 1748
rect 4294 1742 4297 1788
rect 4366 1762 4369 1788
rect 4270 1692 4273 1718
rect 4254 1662 4257 1668
rect 4262 1582 4265 1668
rect 4286 1662 4289 1668
rect 4274 1648 4278 1651
rect 4286 1631 4289 1658
rect 4278 1628 4289 1631
rect 4254 1552 4257 1568
rect 4154 1548 4158 1551
rect 4142 1542 4145 1548
rect 4166 1542 4169 1548
rect 4242 1538 4246 1541
rect 4250 1538 4257 1541
rect 4098 1518 4102 1521
rect 4094 1472 4097 1478
rect 4142 1472 4145 1478
rect 4122 1459 4126 1461
rect 4174 1462 4177 1498
rect 4186 1468 4190 1471
rect 4122 1458 4129 1459
rect 4162 1458 4166 1461
rect 4158 1442 4161 1448
rect 4182 1442 4185 1458
rect 4190 1452 4193 1458
rect 4198 1432 4201 1538
rect 4206 1522 4209 1538
rect 4222 1532 4225 1538
rect 4234 1518 4238 1521
rect 4238 1482 4241 1498
rect 4206 1462 4209 1468
rect 4214 1451 4217 1468
rect 4206 1448 4217 1451
rect 4062 1292 4065 1338
rect 4070 1282 4073 1288
rect 4050 1268 4054 1271
rect 4078 1262 4081 1378
rect 4098 1348 4102 1351
rect 4118 1342 4121 1368
rect 4134 1342 4137 1347
rect 4098 1338 4102 1341
rect 4094 1292 4097 1328
rect 4102 1262 4105 1268
rect 4130 1258 4134 1261
rect 4022 1242 4025 1248
rect 4150 1192 4153 1398
rect 4206 1332 4209 1448
rect 4214 1442 4217 1448
rect 4254 1392 4257 1538
rect 4246 1372 4249 1378
rect 4214 1352 4217 1358
rect 4226 1348 4230 1351
rect 4262 1351 4265 1508
rect 4270 1502 4273 1528
rect 4278 1482 4281 1628
rect 4286 1592 4289 1608
rect 4294 1572 4297 1738
rect 4302 1732 4305 1748
rect 4302 1682 4305 1728
rect 4318 1722 4321 1758
rect 4334 1752 4337 1758
rect 4382 1752 4385 1778
rect 4406 1762 4409 1848
rect 4424 1803 4426 1807
rect 4430 1803 4433 1807
rect 4437 1803 4440 1807
rect 4358 1722 4361 1738
rect 4390 1722 4393 1738
rect 4322 1688 4326 1691
rect 4322 1668 4326 1671
rect 4326 1642 4329 1668
rect 4334 1662 4337 1698
rect 4334 1592 4337 1648
rect 4286 1542 4289 1548
rect 4258 1348 4265 1351
rect 4270 1352 4273 1468
rect 4282 1459 4286 1461
rect 4282 1458 4289 1459
rect 4278 1362 4281 1398
rect 4302 1382 4305 1548
rect 4310 1542 4313 1568
rect 4330 1548 4334 1551
rect 4318 1542 4321 1548
rect 4318 1482 4321 1498
rect 4350 1482 4353 1548
rect 4306 1358 4310 1361
rect 4278 1352 4281 1358
rect 4246 1312 4249 1328
rect 4254 1322 4257 1348
rect 4286 1332 4289 1348
rect 4270 1322 4273 1328
rect 4166 1172 4169 1268
rect 4174 1262 4177 1268
rect 4034 1158 4038 1161
rect 4070 1152 4073 1168
rect 4026 1148 4030 1151
rect 4006 1142 4009 1148
rect 4014 1122 4017 1148
rect 4034 1118 4038 1121
rect 3990 1072 3993 1118
rect 4022 1082 4025 1118
rect 4078 1112 4081 1148
rect 4038 1092 4041 1108
rect 4086 1092 4089 1128
rect 3978 1068 3982 1071
rect 3958 1052 3961 1058
rect 3922 1048 3926 1051
rect 3822 948 3830 951
rect 3774 922 3777 938
rect 3806 882 3809 938
rect 3818 928 3822 931
rect 3814 892 3817 898
rect 3826 878 3830 881
rect 3646 862 3649 868
rect 3678 862 3681 868
rect 3658 858 3662 861
rect 3570 778 3574 781
rect 3510 742 3513 758
rect 3494 702 3497 738
rect 3510 732 3513 738
rect 3518 732 3521 778
rect 3590 772 3593 858
rect 3430 672 3433 688
rect 3454 682 3457 688
rect 3502 682 3505 718
rect 3526 692 3529 768
rect 3562 748 3566 751
rect 3534 742 3537 748
rect 3554 738 3558 741
rect 3526 682 3529 688
rect 3534 672 3537 738
rect 3554 728 3558 731
rect 3606 722 3609 748
rect 3614 732 3617 748
rect 3554 678 3558 681
rect 3418 668 3422 671
rect 3438 662 3441 668
rect 3362 658 3366 661
rect 3366 642 3369 658
rect 3400 603 3402 607
rect 3406 603 3409 607
rect 3413 603 3416 607
rect 3326 472 3329 518
rect 3346 468 3350 471
rect 3274 458 3278 461
rect 3266 448 3270 451
rect 3254 392 3257 438
rect 3246 281 3249 298
rect 3278 292 3281 458
rect 3290 448 3294 451
rect 3302 352 3305 418
rect 3294 342 3297 348
rect 3246 278 3257 281
rect 3254 272 3257 278
rect 3262 262 3265 288
rect 3282 268 3286 271
rect 3294 262 3297 288
rect 3250 248 3254 251
rect 3262 242 3265 248
rect 3278 202 3281 238
rect 3230 82 3233 88
rect 3230 62 3233 68
rect 3254 62 3257 68
rect 3262 62 3265 178
rect 3302 152 3305 328
rect 3310 252 3313 298
rect 3318 282 3321 468
rect 3358 462 3361 468
rect 3326 442 3329 458
rect 3346 448 3350 451
rect 3358 442 3361 448
rect 3326 422 3329 428
rect 3330 388 3334 391
rect 3366 352 3369 528
rect 3374 522 3377 548
rect 3382 462 3385 468
rect 3422 462 3425 638
rect 3446 632 3449 668
rect 3454 662 3457 668
rect 3502 662 3505 668
rect 3538 658 3542 661
rect 3478 652 3481 658
rect 3454 552 3457 568
rect 3462 552 3465 648
rect 3510 642 3513 658
rect 3566 642 3569 648
rect 3486 562 3489 618
rect 3518 592 3521 608
rect 3534 552 3537 618
rect 3498 548 3502 551
rect 3462 542 3465 548
rect 3526 542 3529 548
rect 3430 522 3433 538
rect 3486 532 3489 538
rect 3534 531 3537 538
rect 3526 528 3537 531
rect 3486 522 3489 528
rect 3502 522 3505 528
rect 3474 518 3478 521
rect 3526 482 3529 528
rect 3542 482 3545 488
rect 3550 482 3553 618
rect 3582 592 3585 628
rect 3614 592 3617 698
rect 3622 662 3625 668
rect 3630 592 3633 858
rect 3670 832 3673 848
rect 3694 812 3697 818
rect 3702 792 3705 798
rect 3710 781 3713 868
rect 3766 862 3769 878
rect 3798 862 3801 868
rect 3722 858 3726 861
rect 3738 858 3742 861
rect 3790 852 3793 858
rect 3806 842 3809 858
rect 3794 838 3798 841
rect 3702 778 3713 781
rect 3814 792 3817 868
rect 3838 852 3841 918
rect 3870 862 3873 928
rect 3886 892 3889 948
rect 3902 912 3905 1018
rect 3974 992 3977 1068
rect 3998 1062 4001 1068
rect 4046 1062 4049 1068
rect 4054 1062 4057 1078
rect 4094 1062 4097 1068
rect 4110 1062 4113 1108
rect 4118 1082 4121 1118
rect 4134 1092 4137 1158
rect 4182 1152 4185 1158
rect 4146 1148 4150 1151
rect 4162 1148 4166 1151
rect 4158 1092 4161 1138
rect 4174 1112 4177 1138
rect 4190 1132 4193 1288
rect 4262 1281 4265 1318
rect 4262 1278 4270 1281
rect 4250 1268 4254 1271
rect 4298 1268 4302 1271
rect 4262 1262 4265 1268
rect 4310 1262 4313 1288
rect 4286 1212 4289 1258
rect 4294 1252 4297 1258
rect 4318 1251 4321 1468
rect 4342 1462 4345 1468
rect 4358 1461 4361 1698
rect 4374 1682 4377 1718
rect 4390 1562 4393 1718
rect 4406 1682 4409 1738
rect 4438 1692 4441 1747
rect 4446 1742 4449 1898
rect 4470 1892 4473 1898
rect 4478 1882 4481 1928
rect 4486 1882 4489 2018
rect 4494 1892 4497 2038
rect 4502 1972 4505 2058
rect 4514 1938 4518 1941
rect 4526 1882 4529 1888
rect 4534 1882 4537 1888
rect 4542 1882 4545 2048
rect 4558 1932 4561 2058
rect 4598 2052 4601 2068
rect 4582 2042 4585 2048
rect 4566 1951 4569 1968
rect 4606 1962 4609 2068
rect 4614 2062 4617 2068
rect 4630 2052 4633 2058
rect 4638 2052 4641 2068
rect 4598 1942 4601 1948
rect 4522 1868 4526 1871
rect 4530 1868 4534 1871
rect 4406 1581 4409 1659
rect 4454 1652 4457 1818
rect 4502 1782 4505 1858
rect 4510 1772 4513 1858
rect 4542 1802 4545 1878
rect 4566 1862 4569 1928
rect 4582 1871 4585 1938
rect 4590 1882 4593 1888
rect 4582 1868 4593 1871
rect 4558 1852 4561 1858
rect 4574 1822 4577 1868
rect 4582 1852 4585 1858
rect 4574 1772 4577 1818
rect 4590 1772 4593 1868
rect 4598 1852 4601 1918
rect 4614 1912 4617 1958
rect 4630 1952 4633 1968
rect 4638 1912 4641 1948
rect 4646 1942 4649 2108
rect 4662 2072 4665 2098
rect 4694 2072 4697 2218
rect 4706 2158 4710 2161
rect 4714 2148 4718 2151
rect 4726 2142 4729 2148
rect 4734 2142 4737 2228
rect 4774 2182 4777 2258
rect 4782 2182 4785 2278
rect 4806 2272 4809 2278
rect 4910 2272 4913 2428
rect 4958 2352 4961 2358
rect 4990 2352 4993 2538
rect 5006 2492 5009 2538
rect 5030 2532 5033 2728
rect 5038 2652 5041 2658
rect 5046 2552 5049 2768
rect 5054 2762 5057 2788
rect 5062 2782 5065 2858
rect 5062 2742 5065 2778
rect 5070 2752 5073 2778
rect 5062 2672 5065 2738
rect 5078 2692 5081 2828
rect 5086 2822 5089 2858
rect 5110 2802 5113 2818
rect 5098 2788 5102 2791
rect 5126 2772 5129 2988
rect 5134 2982 5137 3428
rect 5150 3372 5153 3458
rect 5146 3318 5150 3321
rect 5158 3311 5161 3468
rect 5178 3458 5182 3461
rect 5190 3392 5193 3418
rect 5198 3362 5201 3528
rect 5214 3502 5217 3698
rect 5230 3512 5233 3818
rect 5290 3748 5294 3751
rect 5246 3682 5249 3698
rect 5254 3692 5257 3747
rect 5270 3671 5273 3748
rect 5298 3728 5302 3731
rect 5294 3702 5297 3718
rect 5278 3682 5281 3688
rect 5266 3668 5273 3671
rect 5238 3482 5241 3638
rect 5246 3551 5249 3558
rect 5246 3472 5249 3528
rect 5262 3501 5265 3668
rect 5278 3552 5281 3658
rect 5286 3562 5289 3618
rect 5294 3552 5297 3658
rect 5278 3542 5281 3548
rect 5294 3538 5297 3548
rect 5254 3498 5265 3501
rect 5230 3462 5233 3468
rect 5246 3452 5249 3468
rect 5246 3392 5249 3448
rect 5202 3348 5206 3351
rect 5222 3342 5225 3348
rect 5242 3338 5246 3341
rect 5158 3308 5169 3311
rect 5146 3268 5150 3271
rect 5158 3262 5161 3288
rect 5150 3252 5153 3258
rect 5166 3252 5169 3308
rect 5142 3162 5145 3168
rect 5150 3142 5153 3248
rect 5162 3238 5166 3241
rect 5174 3222 5177 3318
rect 5202 3288 5206 3291
rect 5182 3282 5185 3288
rect 5146 3058 5150 3061
rect 5150 2942 5153 2948
rect 5134 2932 5137 2938
rect 5142 2862 5145 2868
rect 5158 2802 5161 3218
rect 5166 3182 5169 3188
rect 5174 3142 5177 3148
rect 5174 3122 5177 3128
rect 5182 3111 5185 3268
rect 5202 3258 5206 3261
rect 5190 3152 5193 3218
rect 5198 3142 5201 3258
rect 5238 3151 5241 3158
rect 5174 3108 5185 3111
rect 5174 3022 5177 3108
rect 5190 3092 5193 3138
rect 5206 3132 5209 3138
rect 5198 3082 5201 3118
rect 5198 2992 5201 3068
rect 5214 3063 5217 3078
rect 5182 2952 5185 2958
rect 5170 2938 5174 2941
rect 5166 2902 5169 2918
rect 5182 2901 5185 2948
rect 5222 2901 5225 3148
rect 5238 3072 5241 3128
rect 5246 3092 5249 3268
rect 5254 3262 5257 3498
rect 5286 3492 5289 3538
rect 5298 3528 5302 3531
rect 5298 3518 5302 3521
rect 5182 2898 5193 2901
rect 5166 2862 5169 2878
rect 5086 2752 5089 2758
rect 5134 2752 5137 2778
rect 5190 2752 5193 2898
rect 5214 2898 5225 2901
rect 5214 2852 5217 2898
rect 5230 2863 5233 2898
rect 5214 2792 5217 2838
rect 5222 2792 5225 2818
rect 5194 2748 5198 2751
rect 5126 2742 5129 2748
rect 5086 2732 5089 2738
rect 5082 2678 5086 2681
rect 5126 2662 5129 2738
rect 5146 2658 5150 2661
rect 5046 2532 5049 2538
rect 5070 2502 5073 2558
rect 5078 2482 5081 2518
rect 5086 2492 5089 2658
rect 5098 2618 5102 2621
rect 5106 2618 5113 2621
rect 5094 2552 5097 2568
rect 5098 2538 5102 2541
rect 5110 2532 5113 2618
rect 5198 2612 5201 2738
rect 5214 2732 5217 2748
rect 5230 2732 5233 2848
rect 5238 2792 5241 3018
rect 5254 2942 5257 3018
rect 5262 2992 5265 3418
rect 5286 3342 5289 3478
rect 5298 3338 5302 3341
rect 5270 3282 5273 3338
rect 5270 3252 5273 3259
rect 5286 3022 5289 3338
rect 5298 3118 5302 3121
rect 5278 3012 5281 3018
rect 5254 2922 5257 2938
rect 5270 2932 5273 2948
rect 5290 2938 5294 2941
rect 5238 2742 5241 2748
rect 5238 2722 5241 2728
rect 5246 2661 5249 2828
rect 5278 2821 5281 2928
rect 5286 2832 5289 2918
rect 5294 2892 5297 2928
rect 5270 2818 5281 2821
rect 5254 2752 5257 2788
rect 5254 2742 5257 2748
rect 5242 2658 5249 2661
rect 5242 2648 5249 2651
rect 5162 2588 5166 2591
rect 5130 2558 5134 2561
rect 5158 2552 5161 2568
rect 5138 2548 5142 2551
rect 5118 2502 5121 2518
rect 5094 2482 5097 2498
rect 5038 2463 5041 2478
rect 5054 2442 5057 2468
rect 4986 2348 4990 2351
rect 4926 2322 4929 2338
rect 4842 2268 4846 2271
rect 4798 2262 4801 2268
rect 4806 2262 4809 2268
rect 4846 2262 4849 2268
rect 4818 2158 4822 2161
rect 4846 2152 4849 2258
rect 4854 2222 4857 2258
rect 4854 2192 4857 2208
rect 4910 2162 4913 2268
rect 4918 2262 4921 2298
rect 4926 2282 4929 2318
rect 4936 2303 4938 2307
rect 4942 2303 4945 2307
rect 4949 2303 4952 2307
rect 4958 2262 4961 2348
rect 4966 2342 4969 2348
rect 4998 2342 5001 2348
rect 4990 2332 4993 2338
rect 5014 2332 5017 2358
rect 5030 2322 5033 2338
rect 5046 2332 5049 2347
rect 5022 2282 5025 2288
rect 4982 2262 4985 2278
rect 5006 2252 5009 2258
rect 4942 2172 4945 2178
rect 4770 2148 4774 2151
rect 4834 2148 4838 2151
rect 4882 2148 4886 2151
rect 4910 2142 4913 2148
rect 4918 2142 4921 2148
rect 4726 2112 4729 2138
rect 4750 2132 4753 2138
rect 4862 2128 4870 2131
rect 4654 2062 4657 2068
rect 4734 2062 4737 2078
rect 4742 2062 4745 2068
rect 4830 2062 4833 2068
rect 4674 2058 4678 2061
rect 4802 2058 4806 2061
rect 4662 2051 4665 2058
rect 4658 2048 4665 2051
rect 4710 2042 4713 2058
rect 4750 2042 4753 2048
rect 4654 2032 4657 2038
rect 4654 1992 4657 2028
rect 4630 1872 4633 1898
rect 4638 1862 4641 1868
rect 4646 1862 4649 1938
rect 4686 1872 4689 2018
rect 4726 1952 4729 2018
rect 4782 1982 4785 1988
rect 4830 1962 4833 1978
rect 4854 1972 4857 2118
rect 4862 2092 4865 2128
rect 4862 2082 4865 2088
rect 4886 2062 4889 2068
rect 4902 2062 4905 2118
rect 4794 1958 4798 1961
rect 4766 1942 4769 1958
rect 4822 1942 4825 1958
rect 4850 1938 4854 1941
rect 4750 1932 4753 1938
rect 4790 1912 4793 1938
rect 4838 1892 4841 1938
rect 4754 1888 4758 1891
rect 4806 1872 4809 1888
rect 4846 1882 4849 1888
rect 4814 1872 4817 1878
rect 4754 1868 4758 1871
rect 4618 1858 4625 1861
rect 4614 1842 4617 1848
rect 4622 1812 4625 1858
rect 4862 1861 4865 2008
rect 4870 1992 4873 2018
rect 4870 1952 4873 1968
rect 4878 1892 4881 1898
rect 4874 1868 4881 1871
rect 4878 1862 4881 1868
rect 4862 1858 4870 1861
rect 4630 1822 4633 1858
rect 4654 1842 4657 1848
rect 4694 1842 4697 1858
rect 4538 1758 4542 1761
rect 4510 1752 4513 1758
rect 4614 1752 4617 1758
rect 4546 1748 4550 1751
rect 4466 1728 4470 1731
rect 4518 1702 4521 1748
rect 4424 1603 4426 1607
rect 4430 1603 4433 1607
rect 4437 1603 4440 1607
rect 4454 1582 4457 1648
rect 4462 1592 4465 1698
rect 4482 1668 4486 1671
rect 4470 1662 4473 1668
rect 4518 1662 4521 1668
rect 4482 1658 4486 1661
rect 4498 1658 4502 1661
rect 4586 1658 4590 1661
rect 4406 1578 4417 1581
rect 4402 1568 4406 1571
rect 4382 1542 4385 1558
rect 4414 1552 4417 1578
rect 4438 1562 4441 1568
rect 4462 1552 4465 1588
rect 4470 1562 4473 1618
rect 4398 1548 4406 1551
rect 4366 1512 4369 1538
rect 4382 1502 4385 1518
rect 4386 1478 4390 1481
rect 4398 1472 4401 1548
rect 4410 1538 4414 1541
rect 4406 1472 4409 1478
rect 4438 1462 4441 1538
rect 4462 1522 4465 1538
rect 4470 1512 4473 1518
rect 4478 1472 4481 1478
rect 4486 1472 4489 1658
rect 4494 1552 4497 1578
rect 4494 1512 4497 1538
rect 4502 1532 4505 1618
rect 4526 1552 4529 1658
rect 4554 1558 4561 1561
rect 4570 1558 4574 1561
rect 4534 1552 4537 1558
rect 4542 1552 4545 1558
rect 4550 1541 4553 1548
rect 4530 1538 4553 1541
rect 4358 1458 4366 1461
rect 4326 1392 4329 1408
rect 4374 1402 4377 1458
rect 4398 1452 4401 1458
rect 4382 1412 4385 1448
rect 4430 1422 4433 1458
rect 4454 1452 4457 1458
rect 4424 1403 4426 1407
rect 4430 1403 4433 1407
rect 4437 1403 4440 1407
rect 4442 1378 4446 1381
rect 4390 1352 4393 1358
rect 4378 1348 4382 1351
rect 4326 1292 4329 1318
rect 4350 1272 4353 1278
rect 4330 1268 4334 1271
rect 4342 1262 4345 1268
rect 4366 1262 4369 1268
rect 4374 1262 4377 1278
rect 4398 1272 4401 1298
rect 4406 1272 4409 1328
rect 4422 1292 4425 1358
rect 4454 1342 4457 1348
rect 4462 1292 4465 1468
rect 4486 1392 4489 1458
rect 4470 1358 4478 1361
rect 4494 1342 4497 1388
rect 4502 1382 4505 1528
rect 4502 1362 4505 1368
rect 4474 1328 4481 1331
rect 4478 1322 4481 1328
rect 4478 1292 4481 1318
rect 4466 1288 4470 1291
rect 4510 1282 4513 1518
rect 4558 1512 4561 1558
rect 4566 1532 4569 1548
rect 4574 1502 4577 1518
rect 4582 1501 4585 1588
rect 4590 1562 4593 1648
rect 4590 1552 4593 1558
rect 4598 1542 4601 1558
rect 4606 1552 4609 1748
rect 4638 1742 4641 1818
rect 4678 1792 4681 1818
rect 4698 1758 4702 1761
rect 4682 1748 4686 1751
rect 4698 1748 4702 1751
rect 4670 1742 4673 1748
rect 4614 1682 4617 1738
rect 4654 1732 4657 1738
rect 4710 1732 4713 1858
rect 4758 1832 4761 1858
rect 4790 1852 4793 1858
rect 4766 1832 4769 1838
rect 4718 1752 4721 1758
rect 4726 1742 4729 1768
rect 4734 1752 4737 1758
rect 4662 1682 4665 1688
rect 4718 1672 4721 1688
rect 4682 1668 4686 1671
rect 4722 1668 4726 1671
rect 4690 1658 4694 1661
rect 4714 1658 4718 1661
rect 4646 1632 4649 1658
rect 4702 1602 4705 1618
rect 4702 1582 4705 1598
rect 4642 1558 4646 1561
rect 4630 1542 4633 1558
rect 4662 1552 4665 1568
rect 4582 1498 4601 1501
rect 4550 1452 4553 1458
rect 4574 1422 4577 1468
rect 4590 1462 4593 1488
rect 4598 1462 4601 1498
rect 4518 1372 4521 1378
rect 4598 1362 4601 1368
rect 4586 1358 4590 1361
rect 4518 1352 4521 1358
rect 4538 1338 4542 1341
rect 4386 1268 4390 1271
rect 4510 1262 4513 1268
rect 4330 1258 4334 1261
rect 4402 1258 4406 1261
rect 4446 1252 4449 1258
rect 4318 1248 4326 1251
rect 4386 1248 4390 1251
rect 4194 1118 4198 1121
rect 4126 1072 4129 1088
rect 4010 1058 4014 1061
rect 4114 1058 4118 1061
rect 4054 1022 4057 1058
rect 3982 971 3985 1018
rect 3974 968 3985 971
rect 3918 932 3921 938
rect 3950 922 3953 948
rect 3862 858 3870 861
rect 3846 792 3849 858
rect 3854 852 3857 858
rect 3678 752 3681 758
rect 3694 752 3697 758
rect 3646 672 3649 698
rect 3670 692 3673 738
rect 3678 662 3681 748
rect 3686 672 3689 688
rect 3690 658 3694 661
rect 3666 648 3670 651
rect 3690 648 3694 651
rect 3678 642 3681 648
rect 3558 562 3561 578
rect 3566 562 3569 568
rect 3586 548 3590 551
rect 3558 472 3561 518
rect 3590 502 3593 538
rect 3598 532 3601 548
rect 3606 512 3609 568
rect 3662 552 3665 638
rect 3690 558 3694 561
rect 3702 552 3705 778
rect 3798 752 3801 758
rect 3814 752 3817 788
rect 3862 772 3865 858
rect 3870 842 3873 848
rect 3878 812 3881 868
rect 3902 862 3905 908
rect 3920 903 3922 907
rect 3926 903 3929 907
rect 3933 903 3936 907
rect 3886 842 3889 848
rect 3710 662 3713 748
rect 3734 722 3737 748
rect 3766 742 3769 747
rect 3802 738 3806 741
rect 3818 738 3822 741
rect 3862 732 3865 748
rect 3878 742 3881 808
rect 3718 672 3721 678
rect 3758 652 3761 658
rect 3650 548 3654 551
rect 3650 538 3654 541
rect 3634 528 3641 531
rect 3606 472 3609 508
rect 3538 468 3542 471
rect 3526 462 3529 468
rect 3466 458 3470 461
rect 3554 458 3558 461
rect 3378 448 3382 451
rect 3390 392 3393 418
rect 3400 403 3402 407
rect 3406 403 3409 407
rect 3413 403 3416 407
rect 3386 348 3390 351
rect 3470 351 3473 418
rect 3486 402 3489 458
rect 3562 448 3566 451
rect 3582 442 3585 448
rect 3598 442 3601 458
rect 3522 438 3526 441
rect 3534 422 3537 428
rect 3534 392 3537 408
rect 3598 392 3601 438
rect 3554 378 3558 381
rect 3606 352 3609 448
rect 3638 392 3641 528
rect 3650 458 3654 461
rect 3662 422 3665 458
rect 3662 402 3665 418
rect 3670 392 3673 538
rect 3686 402 3689 538
rect 3718 502 3721 538
rect 3726 522 3729 528
rect 3766 472 3769 668
rect 3782 662 3785 698
rect 3814 692 3817 728
rect 3870 702 3873 738
rect 3870 682 3873 698
rect 3886 692 3889 788
rect 3910 672 3913 868
rect 3950 862 3953 888
rect 3958 872 3961 888
rect 3966 882 3969 918
rect 3974 872 3977 968
rect 3990 932 3993 938
rect 4014 932 4017 948
rect 4002 888 4006 891
rect 3922 858 3926 861
rect 3970 858 3974 861
rect 3938 848 3942 851
rect 3918 762 3921 768
rect 3950 752 3953 768
rect 3966 752 3969 758
rect 3974 752 3977 758
rect 3958 742 3961 748
rect 3938 738 3942 741
rect 3974 732 3977 738
rect 3982 732 3985 818
rect 4014 802 4017 878
rect 4038 872 4041 948
rect 4014 761 4017 798
rect 4038 762 4041 788
rect 4054 782 4057 1018
rect 4102 1012 4105 1058
rect 4150 1052 4153 1078
rect 4178 1068 4182 1071
rect 4166 1062 4169 1068
rect 4202 1058 4206 1061
rect 4214 1061 4217 1188
rect 4326 1182 4329 1248
rect 4334 1192 4337 1248
rect 4358 1192 4361 1248
rect 4422 1242 4425 1248
rect 4510 1221 4513 1258
rect 4502 1218 4513 1221
rect 4246 1092 4249 1168
rect 4354 1158 4358 1161
rect 4366 1152 4369 1168
rect 4382 1162 4385 1168
rect 4386 1148 4390 1151
rect 4254 1132 4257 1148
rect 4294 1142 4297 1148
rect 4278 1122 4281 1138
rect 4326 1132 4329 1138
rect 4346 1128 4350 1131
rect 4326 1092 4329 1128
rect 4358 1122 4361 1148
rect 4398 1142 4401 1148
rect 4406 1142 4409 1168
rect 4350 1092 4353 1118
rect 4398 1102 4401 1138
rect 4414 1122 4417 1208
rect 4424 1203 4426 1207
rect 4430 1203 4433 1207
rect 4437 1203 4440 1207
rect 4462 1182 4465 1218
rect 4502 1172 4505 1218
rect 4526 1172 4529 1338
rect 4574 1322 4577 1338
rect 4542 1302 4545 1318
rect 4574 1272 4577 1278
rect 4582 1262 4585 1358
rect 4594 1348 4598 1351
rect 4590 1271 4593 1318
rect 4606 1292 4609 1508
rect 4614 1502 4617 1538
rect 4622 1512 4625 1518
rect 4630 1512 4633 1528
rect 4654 1492 4657 1548
rect 4670 1541 4673 1578
rect 4686 1562 4689 1568
rect 4702 1562 4705 1568
rect 4666 1538 4673 1541
rect 4734 1552 4737 1728
rect 4742 1662 4745 1828
rect 4846 1762 4849 1858
rect 4862 1762 4865 1858
rect 4874 1848 4878 1851
rect 4846 1752 4849 1758
rect 4866 1748 4870 1751
rect 4798 1742 4801 1747
rect 4830 1742 4833 1748
rect 4878 1742 4881 1778
rect 4886 1742 4889 2058
rect 4926 2002 4929 2148
rect 4936 2103 4938 2107
rect 4942 2103 4945 2107
rect 4949 2103 4952 2107
rect 4958 2062 4961 2198
rect 4998 2182 5001 2218
rect 5030 2202 5033 2278
rect 5042 2268 5046 2271
rect 5022 2152 5025 2158
rect 5030 2152 5033 2158
rect 4970 2148 4974 2151
rect 4894 1862 4897 1918
rect 4850 1738 4854 1741
rect 4814 1732 4817 1738
rect 4886 1732 4889 1738
rect 4902 1722 4905 1928
rect 4922 1918 4926 1921
rect 4918 1892 4921 1908
rect 4936 1903 4938 1907
rect 4942 1903 4945 1907
rect 4949 1903 4952 1907
rect 4926 1882 4929 1888
rect 4742 1652 4745 1658
rect 4734 1472 4737 1548
rect 4622 1462 4625 1468
rect 4638 1392 4641 1398
rect 4618 1358 4622 1361
rect 4654 1352 4657 1468
rect 4698 1458 4702 1461
rect 4750 1452 4753 1698
rect 4774 1672 4777 1678
rect 4786 1668 4790 1671
rect 4862 1662 4865 1668
rect 4894 1662 4897 1688
rect 4910 1671 4913 1858
rect 4950 1851 4953 1868
rect 4958 1862 4961 1878
rect 4966 1872 4969 2058
rect 4974 2032 4977 2148
rect 4982 2092 4985 2148
rect 5014 2141 5017 2148
rect 5054 2142 5057 2148
rect 5014 2138 5025 2141
rect 4994 2128 4998 2131
rect 5022 2092 5025 2138
rect 5046 2092 5049 2118
rect 5014 2062 5017 2068
rect 5002 2058 5006 2061
rect 5042 2058 5046 2061
rect 4990 2022 4993 2058
rect 5018 1948 5022 1951
rect 4982 1912 4985 1947
rect 5018 1938 5025 1941
rect 4998 1932 5001 1938
rect 4982 1882 4985 1888
rect 4950 1848 4961 1851
rect 4946 1738 4950 1741
rect 4936 1703 4938 1707
rect 4942 1703 4945 1707
rect 4949 1703 4952 1707
rect 4906 1668 4913 1671
rect 4918 1672 4921 1678
rect 4770 1658 4774 1661
rect 4882 1658 4886 1661
rect 4758 1652 4761 1658
rect 4822 1652 4825 1658
rect 4822 1552 4825 1558
rect 4830 1552 4833 1558
rect 4838 1552 4841 1558
rect 4862 1552 4865 1638
rect 4878 1572 4881 1648
rect 4902 1602 4905 1668
rect 4958 1622 4961 1848
rect 4974 1831 4977 1848
rect 4982 1842 4985 1848
rect 4974 1828 4985 1831
rect 4982 1792 4985 1828
rect 4998 1772 5001 1928
rect 5014 1882 5017 1888
rect 5006 1872 5009 1878
rect 5022 1872 5025 1938
rect 5030 1872 5033 2028
rect 5046 1952 5049 1958
rect 5042 1938 5046 1941
rect 5046 1882 5049 1918
rect 5030 1862 5033 1868
rect 5010 1858 5014 1861
rect 5042 1858 5046 1861
rect 5014 1812 5017 1818
rect 5054 1792 5057 2068
rect 5062 2062 5065 2378
rect 5070 2252 5073 2458
rect 5078 2452 5081 2468
rect 5126 2452 5129 2548
rect 5158 2522 5161 2538
rect 5190 2492 5193 2498
rect 5198 2492 5201 2608
rect 5218 2548 5222 2551
rect 5206 2472 5209 2548
rect 5246 2542 5249 2648
rect 5262 2581 5265 2748
rect 5270 2592 5273 2818
rect 5278 2742 5281 2748
rect 5286 2732 5289 2808
rect 5302 2792 5305 2948
rect 5286 2692 5289 2728
rect 5262 2578 5273 2581
rect 5262 2552 5265 2558
rect 5150 2462 5153 2468
rect 5206 2462 5209 2468
rect 5078 2392 5081 2448
rect 5134 2392 5137 2458
rect 5150 2442 5153 2458
rect 5122 2388 5126 2391
rect 5070 2222 5073 2248
rect 5078 2212 5081 2388
rect 5110 2362 5113 2368
rect 5150 2352 5153 2438
rect 5174 2352 5177 2448
rect 5222 2392 5225 2459
rect 5242 2358 5246 2361
rect 5254 2352 5257 2518
rect 5270 2482 5273 2578
rect 5278 2522 5281 2528
rect 5278 2418 5286 2421
rect 5262 2352 5265 2388
rect 5278 2372 5281 2418
rect 5270 2362 5273 2368
rect 5278 2352 5281 2358
rect 5294 2352 5297 2408
rect 5074 2188 5078 2191
rect 5078 2132 5081 2168
rect 5086 2162 5089 2298
rect 5126 2282 5129 2338
rect 5158 2292 5161 2348
rect 5146 2288 5150 2291
rect 5174 2282 5177 2338
rect 5214 2332 5217 2338
rect 5222 2312 5225 2348
rect 5242 2338 5246 2341
rect 5254 2312 5257 2348
rect 5102 2272 5105 2278
rect 5174 2272 5177 2278
rect 5146 2268 5150 2271
rect 5150 2262 5153 2268
rect 5198 2262 5201 2268
rect 5106 2258 5110 2261
rect 5134 2162 5137 2168
rect 5142 2161 5145 2218
rect 5150 2192 5153 2248
rect 5158 2242 5161 2258
rect 5182 2192 5185 2218
rect 5198 2192 5201 2198
rect 5142 2158 5153 2161
rect 5150 2152 5153 2158
rect 5166 2152 5169 2158
rect 5174 2152 5177 2158
rect 5114 2148 5118 2151
rect 5138 2148 5142 2151
rect 5146 2138 5150 2141
rect 5086 2081 5089 2118
rect 5102 2112 5105 2138
rect 5110 2122 5113 2138
rect 5118 2092 5121 2128
rect 5126 2092 5129 2138
rect 5078 2078 5089 2081
rect 5070 2072 5073 2078
rect 5078 2052 5081 2078
rect 5086 2062 5089 2068
rect 5110 2062 5113 2068
rect 5086 2042 5089 2048
rect 5102 2032 5105 2058
rect 5062 1962 5065 1968
rect 5126 1961 5129 2088
rect 5158 2062 5161 2078
rect 5118 1958 5129 1961
rect 5062 1942 5065 1958
rect 5062 1872 5065 1908
rect 5094 1862 5097 1868
rect 5118 1862 5121 1958
rect 5126 1942 5129 1948
rect 5134 1922 5137 2038
rect 5150 1932 5153 1938
rect 5182 1922 5185 2178
rect 5190 2132 5193 2138
rect 5214 2082 5217 2308
rect 5258 2288 5262 2291
rect 5294 2282 5297 2348
rect 5302 2342 5305 2378
rect 5302 2262 5305 2338
rect 5266 2258 5270 2261
rect 5222 2191 5225 2258
rect 5222 2188 5233 2191
rect 5230 2152 5233 2188
rect 5222 2092 5225 2098
rect 5230 2082 5233 2148
rect 5198 2072 5201 2078
rect 5226 2068 5230 2071
rect 5230 1952 5233 2068
rect 5238 2062 5241 2228
rect 5266 2218 5270 2221
rect 5254 2152 5257 2168
rect 5254 2062 5257 2088
rect 5262 2061 5265 2198
rect 5286 2182 5289 2218
rect 5274 2068 5278 2071
rect 5262 2058 5273 2061
rect 5282 2058 5286 2061
rect 5246 2022 5249 2058
rect 5262 1962 5265 1968
rect 5126 1891 5129 1918
rect 5126 1888 5134 1891
rect 5142 1862 5145 1878
rect 5106 1858 5110 1861
rect 4970 1758 4974 1761
rect 4906 1598 4913 1601
rect 4886 1562 4889 1568
rect 4762 1547 4766 1550
rect 4850 1548 4854 1551
rect 4898 1548 4902 1551
rect 4806 1542 4809 1548
rect 4814 1542 4817 1548
rect 4850 1538 4854 1541
rect 4798 1532 4801 1538
rect 4862 1531 4865 1548
rect 4854 1528 4865 1531
rect 4878 1532 4881 1548
rect 4910 1542 4913 1598
rect 4926 1552 4929 1568
rect 4758 1472 4761 1488
rect 4766 1462 4769 1478
rect 4670 1422 4673 1438
rect 4702 1392 4705 1408
rect 4686 1362 4689 1378
rect 4742 1362 4745 1418
rect 4774 1382 4777 1468
rect 4782 1462 4785 1468
rect 4790 1462 4793 1488
rect 4838 1482 4841 1488
rect 4814 1472 4817 1478
rect 4822 1472 4825 1478
rect 4854 1472 4857 1528
rect 4862 1492 4865 1518
rect 4870 1482 4873 1518
rect 4806 1462 4809 1468
rect 4818 1458 4822 1461
rect 4846 1452 4849 1458
rect 4794 1428 4798 1431
rect 4790 1392 4793 1418
rect 4826 1378 4830 1381
rect 4718 1352 4721 1358
rect 4806 1352 4809 1358
rect 4634 1348 4638 1351
rect 4786 1348 4793 1351
rect 4618 1338 4622 1341
rect 4650 1338 4654 1341
rect 4670 1332 4673 1338
rect 4622 1272 4625 1288
rect 4590 1268 4601 1271
rect 4542 1252 4545 1259
rect 4546 1158 4558 1161
rect 4470 1142 4473 1148
rect 4238 1082 4241 1088
rect 4254 1072 4257 1088
rect 4234 1068 4238 1071
rect 4214 1058 4222 1061
rect 4174 1052 4177 1058
rect 4210 1048 4217 1051
rect 4142 1042 4145 1048
rect 4110 952 4113 1018
rect 4166 992 4169 1048
rect 4190 1002 4193 1018
rect 4198 992 4201 1048
rect 4214 992 4217 1048
rect 4134 952 4137 978
rect 4074 948 4078 951
rect 4070 922 4073 938
rect 4086 902 4089 938
rect 4094 922 4097 928
rect 4110 902 4113 948
rect 4134 932 4137 938
rect 4094 882 4097 888
rect 4062 863 4065 868
rect 4078 842 4081 868
rect 4014 758 4025 761
rect 3998 752 4001 758
rect 4010 748 4014 751
rect 3990 742 3993 748
rect 3920 703 3922 707
rect 3926 703 3929 707
rect 3933 703 3936 707
rect 3982 692 3985 728
rect 3990 682 3993 738
rect 3926 672 3929 678
rect 3998 671 4001 738
rect 3994 668 4001 671
rect 4022 672 4025 758
rect 4050 758 4054 761
rect 4030 752 4033 758
rect 4062 752 4065 768
rect 4074 758 4078 761
rect 4086 752 4089 778
rect 4102 752 4105 878
rect 4114 868 4118 871
rect 4142 862 4145 988
rect 4198 962 4201 968
rect 4206 962 4209 968
rect 4222 952 4225 958
rect 4186 948 4193 951
rect 4202 948 4206 951
rect 4190 942 4193 948
rect 4178 938 4182 941
rect 4222 932 4225 938
rect 4150 902 4153 928
rect 4150 862 4153 868
rect 4110 752 4113 758
rect 4086 738 4094 741
rect 4062 732 4065 738
rect 4030 672 4033 718
rect 4062 702 4065 728
rect 4086 722 4089 738
rect 3782 542 3785 658
rect 3838 652 3841 668
rect 3846 652 3849 668
rect 3862 662 3865 668
rect 3870 662 3873 668
rect 3790 551 3793 578
rect 3782 492 3785 508
rect 3790 482 3793 518
rect 3806 492 3809 628
rect 3858 578 3862 581
rect 3870 552 3873 658
rect 3958 652 3961 659
rect 3878 552 3881 578
rect 3886 562 3889 588
rect 3898 548 3902 551
rect 3822 532 3825 538
rect 3830 482 3833 548
rect 3886 542 3889 548
rect 3918 542 3921 568
rect 3974 562 3977 668
rect 3990 662 3993 668
rect 4002 658 4006 661
rect 4026 658 4030 661
rect 4018 648 4030 651
rect 3998 592 4001 618
rect 4002 568 4006 571
rect 3954 558 3958 561
rect 4030 552 4033 578
rect 3954 548 3958 551
rect 4018 548 4022 551
rect 3962 538 3966 541
rect 3950 532 3953 538
rect 3938 528 3942 531
rect 3854 482 3857 508
rect 3878 502 3881 518
rect 3920 503 3922 507
rect 3926 503 3929 507
rect 3933 503 3936 507
rect 3974 502 3977 548
rect 3982 542 3985 548
rect 3990 542 3993 548
rect 3998 542 4001 548
rect 3982 522 3985 538
rect 4022 532 4025 538
rect 4030 532 4033 538
rect 3714 468 3718 471
rect 3702 442 3705 448
rect 3710 442 3713 458
rect 3622 352 3625 358
rect 3366 342 3369 348
rect 3546 348 3550 351
rect 3570 348 3574 351
rect 3582 342 3585 348
rect 3646 342 3649 348
rect 3566 338 3574 341
rect 3342 272 3345 278
rect 3338 258 3342 261
rect 3374 252 3377 259
rect 3334 242 3337 248
rect 3382 172 3385 268
rect 3390 202 3393 328
rect 3438 292 3441 298
rect 3470 262 3473 318
rect 3482 278 3486 281
rect 3518 272 3521 278
rect 3534 263 3537 268
rect 3498 258 3502 261
rect 3400 203 3402 207
rect 3406 203 3409 207
rect 3413 203 3416 207
rect 3390 191 3393 198
rect 3390 188 3398 191
rect 3318 142 3321 168
rect 3334 151 3337 158
rect 3422 152 3425 168
rect 3430 142 3433 148
rect 3358 92 3361 98
rect 3310 72 3313 78
rect 3314 68 3318 71
rect 3414 62 3417 138
rect 3454 132 3457 228
rect 3462 192 3465 258
rect 3478 172 3481 258
rect 3542 192 3545 338
rect 3470 152 3473 158
rect 3478 152 3481 168
rect 3550 152 3553 218
rect 3566 192 3569 338
rect 3578 328 3582 331
rect 3598 302 3601 328
rect 3614 292 3617 318
rect 3622 272 3625 298
rect 3646 292 3649 328
rect 3654 292 3657 358
rect 3694 352 3697 428
rect 3710 362 3713 408
rect 3718 382 3721 468
rect 3742 462 3745 468
rect 3738 448 3742 451
rect 3758 432 3761 458
rect 3730 388 3734 391
rect 3758 372 3761 428
rect 3766 372 3769 468
rect 3774 452 3777 458
rect 3790 392 3793 468
rect 3826 458 3830 461
rect 3726 352 3729 358
rect 3666 348 3670 351
rect 3678 322 3681 338
rect 3686 332 3689 338
rect 3670 272 3673 278
rect 3678 272 3681 298
rect 3622 212 3625 258
rect 3646 222 3649 248
rect 3670 242 3673 258
rect 3654 232 3657 238
rect 3654 192 3657 198
rect 3678 172 3681 268
rect 3702 252 3705 348
rect 3710 342 3713 348
rect 3718 292 3721 338
rect 3710 282 3713 288
rect 3718 278 3726 281
rect 3718 271 3721 278
rect 3714 268 3721 271
rect 3698 248 3702 251
rect 3582 162 3585 168
rect 3678 162 3681 168
rect 3606 152 3609 158
rect 3654 152 3657 158
rect 3694 152 3697 188
rect 3702 152 3705 238
rect 3726 222 3729 258
rect 3734 182 3737 368
rect 3742 352 3745 358
rect 3766 352 3769 358
rect 3754 348 3758 351
rect 3770 338 3774 341
rect 3742 292 3745 328
rect 3750 322 3753 338
rect 3782 332 3785 348
rect 3766 328 3774 331
rect 3750 242 3753 268
rect 3758 262 3761 298
rect 3766 252 3769 328
rect 3790 282 3793 378
rect 3790 272 3793 278
rect 3798 272 3801 398
rect 3822 392 3825 448
rect 3862 362 3865 468
rect 3878 452 3881 498
rect 4006 482 4009 498
rect 3898 468 3902 471
rect 3930 468 3934 471
rect 3978 468 3982 471
rect 3990 462 3993 478
rect 4030 472 4033 478
rect 4018 458 4022 461
rect 3926 452 3929 458
rect 3810 358 3814 361
rect 3838 352 3841 358
rect 3830 342 3833 348
rect 3818 328 3822 331
rect 3834 328 3838 331
rect 3822 272 3825 308
rect 3830 272 3833 278
rect 3798 262 3801 268
rect 3838 262 3841 268
rect 3810 258 3814 261
rect 3794 248 3798 251
rect 3766 192 3769 248
rect 3782 242 3785 248
rect 3814 242 3817 258
rect 3846 241 3849 338
rect 3854 292 3857 328
rect 3862 302 3865 358
rect 3854 252 3857 288
rect 3846 238 3857 241
rect 3746 188 3750 191
rect 3814 191 3817 218
rect 3806 188 3817 191
rect 3854 192 3857 238
rect 3734 152 3737 178
rect 3466 148 3470 151
rect 3514 148 3518 151
rect 3642 148 3646 151
rect 3806 151 3809 188
rect 3838 162 3841 168
rect 3486 142 3489 148
rect 3526 132 3529 148
rect 3438 92 3441 118
rect 3454 112 3457 128
rect 3466 88 3470 91
rect 3482 88 3486 91
rect 3494 82 3497 118
rect 3534 102 3537 128
rect 3566 122 3569 148
rect 3606 142 3609 148
rect 3702 142 3705 148
rect 3822 142 3825 158
rect 3626 138 3630 141
rect 3650 138 3654 141
rect 3682 138 3686 141
rect 3626 128 3630 131
rect 3682 128 3686 131
rect 3590 102 3593 128
rect 3710 112 3713 118
rect 3426 68 3430 71
rect 3542 63 3545 88
rect 3606 82 3609 98
rect 3854 92 3857 148
rect 3862 142 3865 218
rect 3870 152 3873 408
rect 3926 392 3929 448
rect 3934 402 3937 458
rect 3946 448 3950 451
rect 3982 432 3985 458
rect 3878 322 3881 358
rect 3886 342 3889 368
rect 3922 348 3926 351
rect 3974 351 3977 418
rect 3982 362 3985 428
rect 4022 422 4025 428
rect 3974 348 3982 351
rect 3886 312 3889 338
rect 3894 332 3897 348
rect 4022 342 4025 418
rect 4030 372 4033 468
rect 4038 462 4041 678
rect 4058 668 4062 671
rect 4054 592 4057 658
rect 4070 652 4073 718
rect 4094 692 4097 728
rect 4102 722 4105 748
rect 4102 682 4105 708
rect 4118 692 4121 728
rect 4086 672 4089 678
rect 4110 672 4113 678
rect 4126 662 4129 668
rect 4134 662 4137 768
rect 4142 762 4145 858
rect 4158 831 4161 868
rect 4150 828 4161 831
rect 4142 742 4145 748
rect 4150 712 4153 828
rect 4166 812 4169 858
rect 4182 852 4185 898
rect 4214 872 4217 898
rect 4206 862 4209 868
rect 4222 862 4225 908
rect 4230 862 4233 918
rect 4238 892 4241 1058
rect 4246 952 4249 1028
rect 4254 942 4257 978
rect 4286 972 4289 1088
rect 4302 1072 4305 1078
rect 4350 1072 4353 1088
rect 4414 1072 4417 1118
rect 4462 1092 4465 1138
rect 4526 1092 4529 1118
rect 4462 1082 4465 1088
rect 4366 1062 4369 1068
rect 4334 1052 4337 1059
rect 4382 1052 4385 1058
rect 4390 1052 4393 1068
rect 4486 1062 4489 1088
rect 4542 1072 4545 1148
rect 4550 1142 4553 1148
rect 4558 1142 4561 1148
rect 4550 1082 4553 1138
rect 4410 1058 4414 1061
rect 4266 958 4270 961
rect 4262 942 4265 948
rect 4278 912 4281 948
rect 4286 942 4289 968
rect 4390 962 4393 1028
rect 4406 992 4409 1048
rect 4494 1012 4497 1058
rect 4534 1051 4537 1058
rect 4530 1048 4537 1051
rect 4424 1003 4426 1007
rect 4430 1003 4433 1007
rect 4437 1003 4440 1007
rect 4302 932 4305 938
rect 4302 882 4305 928
rect 4334 892 4337 948
rect 4374 932 4377 938
rect 4374 892 4377 918
rect 4286 862 4289 878
rect 4390 871 4393 958
rect 4406 932 4409 948
rect 4382 868 4393 871
rect 4198 852 4201 858
rect 4182 832 4185 848
rect 4158 762 4161 808
rect 4166 762 4169 778
rect 4158 732 4161 758
rect 4174 752 4177 828
rect 4198 792 4201 828
rect 4182 732 4185 748
rect 4190 732 4193 738
rect 4142 672 4145 698
rect 4150 662 4153 708
rect 4214 692 4217 858
rect 4190 662 4193 688
rect 4222 682 4225 708
rect 4198 672 4201 678
rect 4230 672 4233 838
rect 4238 752 4241 848
rect 4254 832 4257 858
rect 4266 848 4270 851
rect 4286 842 4289 848
rect 4294 762 4297 768
rect 4302 762 4305 868
rect 4342 862 4345 868
rect 4358 862 4361 868
rect 4366 862 4369 868
rect 4314 858 4318 861
rect 4346 748 4350 751
rect 4278 732 4281 738
rect 4334 732 4337 748
rect 4334 692 4337 728
rect 4298 668 4302 671
rect 4202 658 4206 661
rect 4298 658 4302 661
rect 4078 652 4081 658
rect 4086 622 4089 658
rect 4046 511 4049 528
rect 4046 508 4057 511
rect 4046 492 4049 498
rect 4038 412 4041 458
rect 4038 392 4041 408
rect 4054 382 4057 508
rect 4042 378 4046 381
rect 3886 272 3889 308
rect 3878 252 3881 258
rect 3886 231 3889 258
rect 3878 228 3889 231
rect 3870 102 3873 138
rect 3714 88 3718 91
rect 3866 88 3870 91
rect 3622 82 3625 88
rect 3774 82 3777 88
rect 3582 72 3585 78
rect 3306 58 3310 61
rect 3558 62 3561 68
rect 3606 62 3609 78
rect 3622 62 3625 68
rect 3578 58 3582 61
rect 3686 62 3689 78
rect 3738 68 3742 71
rect 3758 62 3761 68
rect 1398 52 1401 58
rect 1494 52 1497 58
rect 2126 52 2129 58
rect 2230 52 2233 58
rect 3598 52 3601 58
rect 3654 52 3657 59
rect 3730 58 3734 61
rect 3838 62 3841 78
rect 3878 62 3881 228
rect 3902 222 3905 318
rect 3920 303 3922 307
rect 3926 303 3929 307
rect 3933 303 3936 307
rect 3910 282 3913 288
rect 3974 282 3977 338
rect 4022 292 4025 328
rect 4022 282 4025 288
rect 4046 272 4049 368
rect 4058 288 4062 291
rect 4046 262 4049 268
rect 3962 258 3966 261
rect 4010 258 4014 261
rect 4038 252 4041 258
rect 4054 242 4057 258
rect 3902 132 3905 208
rect 3926 162 3929 238
rect 4046 192 4049 228
rect 4054 182 4057 238
rect 4078 202 4081 358
rect 3998 152 4001 168
rect 4058 158 4062 161
rect 4078 152 4081 198
rect 3918 142 3921 148
rect 3974 142 3977 148
rect 4074 138 4078 141
rect 3886 122 3889 128
rect 3920 103 3922 107
rect 3926 103 3929 107
rect 3933 103 3936 107
rect 3898 88 3902 91
rect 3942 82 3945 98
rect 3950 92 3953 128
rect 3966 82 3969 128
rect 4030 122 4033 138
rect 4054 132 4057 138
rect 4038 122 4041 128
rect 3890 68 3894 71
rect 3910 62 3913 68
rect 4014 63 4017 88
rect 4030 72 4033 78
rect 3806 52 3809 59
rect 3882 58 3886 61
rect 4046 62 4049 118
rect 4058 88 4062 91
rect 4094 82 4097 618
rect 4134 602 4137 658
rect 4318 652 4321 678
rect 4170 648 4174 651
rect 4194 618 4198 621
rect 4110 552 4113 588
rect 4214 572 4217 618
rect 4302 592 4305 648
rect 4314 638 4318 641
rect 4202 568 4206 571
rect 4134 542 4137 558
rect 4150 542 4153 568
rect 4222 562 4225 568
rect 4334 552 4337 618
rect 4342 552 4345 618
rect 4358 582 4361 858
rect 4382 782 4385 868
rect 4430 862 4433 988
rect 4442 958 4446 961
rect 4454 952 4457 968
rect 4474 948 4478 951
rect 4466 938 4470 941
rect 4486 932 4489 988
rect 4510 942 4513 948
rect 4526 942 4529 1008
rect 4494 932 4497 938
rect 4506 928 4510 931
rect 4542 922 4545 947
rect 4402 858 4406 861
rect 4390 842 4393 858
rect 4430 852 4433 858
rect 4390 792 4393 808
rect 4414 782 4417 818
rect 4424 803 4426 807
rect 4430 803 4433 807
rect 4437 803 4440 807
rect 4418 758 4422 761
rect 4430 752 4433 778
rect 4446 772 4449 908
rect 4454 872 4457 878
rect 4470 862 4473 868
rect 4478 862 4481 918
rect 4510 892 4513 918
rect 4550 892 4553 1058
rect 4558 1002 4561 1068
rect 4566 1062 4569 1138
rect 4574 1082 4577 1148
rect 4582 1142 4585 1258
rect 4590 1252 4593 1258
rect 4598 1252 4601 1268
rect 4606 1252 4609 1258
rect 4630 1192 4633 1258
rect 4646 1202 4649 1218
rect 4654 1192 4657 1238
rect 4662 1212 4665 1218
rect 4670 1192 4673 1328
rect 4638 1182 4641 1188
rect 4662 1172 4665 1178
rect 4670 1162 4673 1168
rect 4678 1162 4681 1348
rect 4702 1342 4705 1348
rect 4734 1342 4737 1348
rect 4758 1342 4761 1348
rect 4766 1342 4769 1348
rect 4738 1328 4742 1331
rect 4774 1312 4777 1348
rect 4762 1288 4766 1291
rect 4694 1262 4697 1268
rect 4622 1152 4625 1158
rect 4594 1148 4598 1151
rect 4674 1148 4678 1151
rect 4594 1138 4598 1141
rect 4586 1128 4590 1131
rect 4586 1088 4590 1091
rect 4586 1048 4590 1051
rect 4502 872 4505 888
rect 4458 858 4462 861
rect 4454 772 4457 838
rect 4390 742 4393 748
rect 4410 728 4414 731
rect 4390 672 4393 678
rect 4398 672 4401 688
rect 4410 658 4414 661
rect 4398 622 4401 658
rect 4422 652 4425 738
rect 4438 692 4441 758
rect 4446 742 4449 768
rect 4462 752 4465 818
rect 4454 712 4457 748
rect 4478 722 4481 738
rect 4424 603 4426 607
rect 4430 603 4433 607
rect 4437 603 4440 607
rect 4194 548 4198 551
rect 4166 542 4169 548
rect 4186 538 4190 541
rect 4150 532 4153 538
rect 4142 472 4145 518
rect 4166 482 4169 538
rect 4246 532 4249 548
rect 4286 542 4289 548
rect 4334 542 4337 548
rect 4446 532 4449 538
rect 4186 528 4190 531
rect 4174 472 4177 478
rect 4230 472 4233 508
rect 4438 492 4441 508
rect 4334 472 4337 478
rect 4146 468 4150 471
rect 4250 468 4254 471
rect 4102 462 4105 468
rect 4126 432 4129 468
rect 4166 422 4169 458
rect 4182 452 4185 458
rect 4190 412 4193 468
rect 4198 462 4201 468
rect 4210 458 4214 461
rect 4298 459 4302 462
rect 4350 462 4353 478
rect 4202 448 4206 451
rect 4270 432 4273 458
rect 4102 351 4105 358
rect 4142 352 4145 388
rect 4166 372 4169 378
rect 4182 352 4185 398
rect 4206 352 4209 358
rect 4238 352 4241 388
rect 4246 362 4249 368
rect 4154 348 4158 351
rect 4186 338 4190 341
rect 4134 332 4137 338
rect 4102 272 4105 328
rect 4102 252 4105 258
rect 4110 162 4113 308
rect 4142 272 4145 288
rect 4182 272 4185 328
rect 4190 272 4193 338
rect 4198 312 4201 348
rect 4230 342 4233 348
rect 4254 332 4257 368
rect 4270 342 4273 428
rect 4346 368 4350 371
rect 4286 351 4289 358
rect 4358 352 4361 478
rect 4374 472 4377 478
rect 4366 462 4369 468
rect 4382 462 4385 468
rect 4394 458 4398 461
rect 4406 452 4409 478
rect 4454 472 4457 708
rect 4478 672 4481 718
rect 4470 542 4473 548
rect 4478 542 4481 658
rect 4486 612 4489 868
rect 4526 862 4529 888
rect 4558 881 4561 918
rect 4554 878 4561 881
rect 4542 872 4545 878
rect 4494 812 4497 858
rect 4502 792 4505 848
rect 4494 782 4497 788
rect 4510 712 4513 728
rect 4510 682 4513 698
rect 4526 662 4529 858
rect 4574 762 4577 948
rect 4590 922 4593 928
rect 4598 902 4601 1138
rect 4606 1102 4609 1138
rect 4614 1122 4617 1148
rect 4614 1071 4617 1118
rect 4638 1102 4641 1148
rect 4650 1138 4654 1141
rect 4686 1132 4689 1218
rect 4654 1092 4657 1118
rect 4610 1068 4617 1071
rect 4622 1072 4625 1088
rect 4630 1062 4633 1068
rect 4638 1062 4641 1068
rect 4614 1042 4617 1048
rect 4646 1042 4649 1068
rect 4662 1061 4665 1098
rect 4658 1058 4665 1061
rect 4670 1062 4673 1088
rect 4630 952 4633 1038
rect 4678 1032 4681 1068
rect 4638 962 4641 1008
rect 4646 972 4649 978
rect 4618 948 4622 951
rect 4614 892 4617 938
rect 4654 932 4657 978
rect 4670 892 4673 948
rect 4686 912 4689 1068
rect 4694 1062 4697 1118
rect 4710 1072 4713 1088
rect 4694 952 4697 1058
rect 4710 1052 4713 1068
rect 4582 882 4585 888
rect 4694 882 4697 938
rect 4702 892 4705 948
rect 4594 878 4601 881
rect 4598 862 4601 878
rect 4718 872 4721 1258
rect 4726 1192 4729 1259
rect 4734 1152 4737 1198
rect 4742 1152 4745 1158
rect 4750 1152 4753 1228
rect 4778 1168 4782 1171
rect 4742 1072 4745 1128
rect 4750 1112 4753 1148
rect 4758 1102 4761 1118
rect 4754 1088 4758 1091
rect 4726 1062 4729 1068
rect 4734 1062 4737 1068
rect 4742 932 4745 1068
rect 4790 1012 4793 1348
rect 4838 1272 4841 1368
rect 4854 1362 4857 1468
rect 4878 1442 4881 1468
rect 4886 1462 4889 1538
rect 4894 1482 4897 1538
rect 4886 1452 4889 1458
rect 4902 1452 4905 1488
rect 4886 1351 4889 1368
rect 4902 1342 4905 1428
rect 4910 1412 4913 1538
rect 4936 1503 4938 1507
rect 4942 1503 4945 1507
rect 4949 1503 4952 1507
rect 4954 1488 4958 1491
rect 4930 1468 4934 1471
rect 4922 1458 4926 1461
rect 4934 1451 4937 1458
rect 4930 1448 4937 1451
rect 4918 1342 4921 1388
rect 4930 1368 4934 1371
rect 4926 1342 4929 1348
rect 4942 1342 4945 1458
rect 4966 1432 4969 1678
rect 4974 1662 4977 1708
rect 4982 1662 4985 1768
rect 5046 1752 5049 1778
rect 5070 1752 5073 1768
rect 5078 1752 5081 1758
rect 5018 1748 5022 1751
rect 5038 1742 5041 1748
rect 4998 1682 5001 1728
rect 5030 1712 5033 1718
rect 5022 1582 5025 1668
rect 5030 1652 5033 1658
rect 5038 1642 5041 1738
rect 5046 1672 5049 1748
rect 5058 1728 5062 1731
rect 5078 1672 5081 1678
rect 5070 1662 5073 1668
rect 5086 1662 5089 1728
rect 5082 1658 5086 1661
rect 5046 1652 5049 1658
rect 5062 1652 5065 1658
rect 5030 1592 5033 1618
rect 4974 1522 4977 1548
rect 4990 1452 4993 1578
rect 5054 1552 5057 1568
rect 5042 1548 5046 1551
rect 5014 1542 5017 1548
rect 5014 1472 5017 1538
rect 5010 1458 5014 1461
rect 4950 1372 4953 1378
rect 4990 1352 4993 1448
rect 5038 1412 5041 1528
rect 5054 1492 5057 1548
rect 5054 1472 5057 1478
rect 5062 1462 5065 1628
rect 5094 1622 5097 1858
rect 5118 1782 5121 1858
rect 5106 1738 5110 1741
rect 5126 1692 5129 1728
rect 5126 1652 5129 1658
rect 5094 1592 5097 1608
rect 5074 1548 5078 1551
rect 5086 1542 5089 1548
rect 5078 1492 5081 1528
rect 5078 1432 5081 1448
rect 4998 1342 5001 1408
rect 5062 1382 5065 1388
rect 5022 1352 5025 1358
rect 5046 1352 5049 1358
rect 5034 1348 5038 1351
rect 5006 1342 5009 1348
rect 5046 1342 5049 1348
rect 5054 1342 5057 1368
rect 5062 1352 5065 1358
rect 4854 1282 4857 1288
rect 4902 1272 4905 1338
rect 4926 1292 4929 1318
rect 4936 1303 4938 1307
rect 4942 1303 4945 1307
rect 4949 1303 4952 1307
rect 4954 1288 4958 1291
rect 4982 1272 4985 1328
rect 4990 1282 4993 1338
rect 5006 1292 5009 1338
rect 5030 1332 5033 1338
rect 5042 1318 5046 1321
rect 4874 1268 4878 1271
rect 4822 1263 4825 1268
rect 4830 1152 4833 1158
rect 4838 1142 4841 1268
rect 4894 1262 4897 1268
rect 4866 1258 4870 1261
rect 4902 1202 4905 1258
rect 4886 1172 4889 1178
rect 4870 1162 4873 1168
rect 4902 1162 4905 1168
rect 4894 1152 4897 1158
rect 4910 1151 4913 1268
rect 4982 1262 4985 1268
rect 5014 1263 5017 1308
rect 5070 1292 5073 1408
rect 5078 1311 5081 1358
rect 5086 1352 5089 1418
rect 5094 1362 5097 1478
rect 5102 1462 5105 1468
rect 5102 1372 5105 1418
rect 5110 1352 5113 1618
rect 5142 1572 5145 1858
rect 5150 1682 5153 1918
rect 5166 1902 5169 1918
rect 5190 1892 5193 1908
rect 5158 1882 5161 1888
rect 5166 1872 5169 1878
rect 5182 1862 5185 1868
rect 5166 1772 5169 1858
rect 5206 1832 5209 1858
rect 5150 1552 5153 1678
rect 5166 1662 5169 1768
rect 5214 1752 5217 1938
rect 5222 1912 5225 1948
rect 5262 1932 5265 1938
rect 5238 1892 5241 1908
rect 5230 1862 5233 1868
rect 5222 1852 5225 1858
rect 5174 1742 5177 1748
rect 5214 1742 5217 1748
rect 5230 1742 5233 1748
rect 5270 1692 5273 2058
rect 5286 1952 5289 1978
rect 5278 1942 5281 1948
rect 5278 1882 5281 1898
rect 5202 1688 5206 1691
rect 5254 1682 5257 1688
rect 5278 1682 5281 1868
rect 5238 1672 5241 1678
rect 5190 1662 5193 1668
rect 5262 1662 5265 1668
rect 5218 1658 5222 1661
rect 5182 1652 5185 1658
rect 5238 1652 5241 1658
rect 5230 1591 5233 1618
rect 5222 1588 5233 1591
rect 5138 1548 5142 1551
rect 5150 1542 5153 1548
rect 5118 1462 5121 1478
rect 5126 1442 5129 1468
rect 5150 1462 5153 1508
rect 5190 1482 5193 1518
rect 5198 1501 5201 1528
rect 5206 1512 5209 1518
rect 5198 1498 5209 1501
rect 5198 1472 5201 1478
rect 5170 1458 5174 1461
rect 5194 1458 5198 1461
rect 5134 1452 5137 1458
rect 5098 1338 5102 1341
rect 5086 1322 5089 1328
rect 5094 1312 5097 1318
rect 5110 1312 5113 1348
rect 5078 1308 5089 1311
rect 5078 1292 5081 1298
rect 5050 1268 5054 1271
rect 4922 1248 4926 1251
rect 4902 1148 4913 1151
rect 4918 1152 4921 1158
rect 4966 1152 4969 1238
rect 4998 1192 5001 1258
rect 5054 1252 5057 1258
rect 5070 1252 5073 1288
rect 4978 1158 4982 1161
rect 4998 1152 5001 1188
rect 5046 1152 5049 1158
rect 5054 1152 5057 1248
rect 4814 1082 4817 1138
rect 4886 1122 4889 1148
rect 4894 1132 4897 1138
rect 4846 1082 4849 1088
rect 4886 1062 4889 1068
rect 4894 1062 4897 1078
rect 4802 1058 4806 1061
rect 4866 1058 4870 1061
rect 4878 1052 4881 1058
rect 4806 962 4809 968
rect 4754 958 4758 961
rect 4830 952 4833 1048
rect 4838 992 4841 1028
rect 4862 992 4865 1038
rect 4746 918 4750 921
rect 4734 882 4737 918
rect 4766 891 4769 938
rect 4766 888 4777 891
rect 4766 872 4769 878
rect 4686 868 4694 871
rect 4698 868 4702 871
rect 4606 862 4609 868
rect 4678 862 4681 868
rect 4614 852 4617 858
rect 4638 842 4641 858
rect 4634 818 4638 821
rect 4654 802 4657 858
rect 4602 758 4606 761
rect 4554 748 4558 751
rect 4558 712 4561 728
rect 4542 682 4545 708
rect 4574 692 4577 748
rect 4498 658 4502 661
rect 4554 658 4558 661
rect 4510 552 4513 578
rect 4566 552 4569 668
rect 4582 662 4585 668
rect 4590 662 4593 678
rect 4614 662 4617 798
rect 4662 792 4665 838
rect 4602 658 4606 661
rect 4598 592 4601 648
rect 4622 592 4625 748
rect 4650 738 4654 741
rect 4654 692 4657 718
rect 4634 668 4649 671
rect 4630 642 4633 658
rect 4638 652 4641 658
rect 4646 602 4649 668
rect 4654 662 4657 678
rect 4670 672 4673 678
rect 4686 672 4689 868
rect 4718 862 4721 868
rect 4718 752 4721 818
rect 4694 692 4697 728
rect 4598 552 4601 568
rect 4586 548 4590 551
rect 4478 512 4481 538
rect 4510 522 4513 548
rect 4518 542 4521 548
rect 4530 538 4534 541
rect 4538 528 4542 531
rect 4470 462 4473 498
rect 4510 462 4513 488
rect 4518 472 4521 478
rect 4574 472 4577 518
rect 4590 482 4593 508
rect 4606 492 4609 518
rect 4630 492 4633 548
rect 4622 482 4625 488
rect 4638 472 4641 568
rect 4498 458 4502 461
rect 4570 458 4574 461
rect 4390 352 4393 358
rect 4406 352 4409 388
rect 4398 342 4401 348
rect 4230 272 4233 288
rect 4126 172 4129 268
rect 4174 262 4177 268
rect 4206 262 4209 268
rect 4194 258 4198 261
rect 4158 252 4161 258
rect 4214 252 4217 258
rect 4246 252 4249 259
rect 4278 252 4281 258
rect 4174 242 4177 248
rect 4294 242 4297 338
rect 4350 292 4353 338
rect 4374 322 4377 328
rect 4334 262 4337 288
rect 4354 278 4358 281
rect 4366 272 4369 288
rect 4374 262 4377 318
rect 4382 272 4385 278
rect 4398 272 4401 288
rect 4414 272 4417 458
rect 4490 448 4494 451
rect 4522 448 4526 451
rect 4438 432 4441 448
rect 4424 403 4426 407
rect 4430 403 4433 407
rect 4437 403 4440 407
rect 4454 351 4457 358
rect 4314 258 4318 261
rect 4394 248 4398 251
rect 4206 192 4209 208
rect 4222 192 4225 238
rect 4102 152 4105 158
rect 4110 152 4113 158
rect 4126 142 4129 168
rect 4114 88 4118 91
rect 4142 82 4145 188
rect 4366 172 4369 248
rect 4382 192 4385 218
rect 4406 212 4409 258
rect 4422 252 4425 258
rect 4430 222 4433 278
rect 4424 203 4426 207
rect 4430 203 4433 207
rect 4437 203 4440 207
rect 4370 168 4374 171
rect 4414 152 4417 168
rect 4446 151 4449 168
rect 4150 112 4153 148
rect 4174 102 4177 128
rect 4094 72 4097 78
rect 4126 62 4129 78
rect 4182 62 4185 98
rect 4254 92 4257 98
rect 4242 88 4246 91
rect 4206 62 4209 68
rect 4246 62 4249 78
rect 4262 72 4265 78
rect 4270 62 4273 148
rect 4282 138 4286 141
rect 4286 92 4289 128
rect 4294 112 4297 118
rect 4302 82 4305 148
rect 4462 142 4465 338
rect 4494 262 4497 268
rect 4502 262 4505 328
rect 4514 318 4518 321
rect 4526 292 4529 358
rect 4518 272 4521 288
rect 4534 282 4537 448
rect 4542 392 4545 428
rect 4542 322 4545 348
rect 4542 292 4545 318
rect 4566 282 4569 338
rect 4510 232 4513 258
rect 4534 252 4537 278
rect 4542 272 4545 278
rect 4562 258 4566 261
rect 4562 248 4566 251
rect 4478 172 4481 218
rect 4518 151 4521 158
rect 4314 138 4318 141
rect 4286 62 4289 68
rect 4326 62 4329 118
rect 4334 62 4337 98
rect 4366 92 4369 128
rect 4406 92 4409 108
rect 4486 102 4489 138
rect 4394 78 4398 81
rect 4414 72 4417 88
rect 4542 82 4545 238
rect 4550 152 4553 158
rect 4566 92 4569 248
rect 4582 192 4585 308
rect 4590 262 4593 348
rect 4606 292 4609 348
rect 4590 252 4593 258
rect 4606 252 4609 258
rect 4590 152 4593 178
rect 4598 142 4601 168
rect 4622 132 4625 428
rect 4638 372 4641 468
rect 4646 462 4649 508
rect 4654 492 4657 608
rect 4646 392 4649 458
rect 4654 442 4657 448
rect 4662 392 4665 668
rect 4742 662 4745 828
rect 4766 821 4769 868
rect 4774 862 4777 888
rect 4758 818 4769 821
rect 4758 742 4761 818
rect 4774 752 4777 758
rect 4758 712 4761 738
rect 4758 672 4761 708
rect 4674 658 4678 661
rect 4714 658 4718 661
rect 4686 648 4694 651
rect 4674 548 4678 551
rect 4686 492 4689 648
rect 4702 632 4705 658
rect 4742 641 4745 658
rect 4742 638 4753 641
rect 4730 618 4734 621
rect 4750 592 4753 638
rect 4718 552 4721 578
rect 4702 532 4705 538
rect 4682 468 4686 471
rect 4714 468 4718 471
rect 4638 352 4641 368
rect 4638 321 4641 338
rect 4654 322 4657 338
rect 4638 318 4649 321
rect 4646 302 4649 318
rect 4662 312 4665 348
rect 4630 272 4633 278
rect 4646 272 4649 298
rect 4670 282 4673 458
rect 4678 362 4681 448
rect 4686 442 4689 448
rect 4702 352 4705 468
rect 4734 452 4737 518
rect 4750 472 4753 528
rect 4766 492 4769 608
rect 4774 492 4777 728
rect 4746 468 4750 471
rect 4718 352 4721 398
rect 4742 352 4745 458
rect 4750 432 4753 458
rect 4762 448 4766 451
rect 4782 372 4785 948
rect 4838 942 4841 948
rect 4830 931 4833 938
rect 4854 932 4857 968
rect 4886 952 4889 1058
rect 4882 948 4886 951
rect 4862 942 4865 948
rect 4902 932 4905 1148
rect 4934 1142 4937 1148
rect 4922 1138 4926 1141
rect 4950 1122 4953 1128
rect 4936 1103 4938 1107
rect 4942 1103 4945 1107
rect 4949 1103 4952 1107
rect 4914 1088 4918 1091
rect 4966 1072 4969 1148
rect 4986 1138 4990 1141
rect 4914 958 4918 961
rect 4934 952 4937 958
rect 4926 942 4929 948
rect 4966 942 4969 1068
rect 4974 1052 4977 1058
rect 4998 962 5001 1148
rect 5038 1142 5041 1148
rect 5006 1112 5009 1118
rect 5014 1092 5017 1098
rect 5070 1072 5073 1128
rect 5086 1112 5089 1308
rect 5110 1282 5113 1288
rect 5094 1252 5097 1258
rect 5102 1222 5105 1268
rect 5118 1212 5121 1348
rect 5126 1272 5129 1438
rect 5134 1392 5137 1448
rect 5142 1352 5145 1458
rect 5150 1452 5153 1458
rect 5158 1422 5161 1458
rect 5206 1442 5209 1498
rect 5222 1462 5225 1588
rect 5238 1542 5241 1548
rect 5238 1482 5241 1518
rect 5246 1462 5249 1468
rect 5178 1358 5182 1361
rect 5186 1348 5190 1351
rect 5198 1342 5201 1348
rect 5206 1342 5209 1398
rect 5242 1348 5246 1351
rect 5146 1338 5150 1341
rect 5222 1332 5225 1338
rect 5118 1162 5121 1168
rect 5102 1102 5105 1158
rect 5114 1148 5118 1151
rect 5126 1142 5129 1268
rect 5150 1262 5153 1298
rect 5206 1292 5209 1318
rect 5190 1262 5193 1268
rect 5134 1162 5137 1168
rect 5150 1152 5153 1198
rect 5158 1142 5161 1218
rect 5166 1152 5169 1158
rect 5174 1152 5177 1228
rect 5214 1192 5217 1308
rect 5246 1262 5249 1268
rect 5194 1148 5198 1151
rect 5110 1082 5113 1138
rect 5118 1092 5121 1138
rect 5126 1132 5129 1138
rect 5078 1063 5081 1068
rect 5014 982 5017 1018
rect 5002 948 5006 951
rect 5038 942 5041 948
rect 4830 928 4841 931
rect 4906 928 4910 931
rect 4798 892 4801 928
rect 4806 901 4809 918
rect 4806 898 4817 901
rect 4814 781 4817 898
rect 4838 892 4841 928
rect 4878 922 4881 928
rect 4826 888 4830 891
rect 4838 882 4841 888
rect 4918 872 4921 938
rect 4946 928 4950 931
rect 4936 903 4938 907
rect 4942 903 4945 907
rect 4949 903 4952 907
rect 4958 892 4961 918
rect 4934 882 4937 888
rect 4970 868 4974 871
rect 4902 863 4905 868
rect 4998 862 5001 878
rect 5014 872 5017 918
rect 5038 892 5041 928
rect 5054 922 5057 968
rect 5054 912 5057 918
rect 5062 892 5065 948
rect 5078 882 5081 908
rect 5094 881 5097 1078
rect 5126 1072 5129 1128
rect 5134 1072 5137 1118
rect 5150 1092 5153 1128
rect 5158 1092 5161 1138
rect 5158 1062 5161 1068
rect 5166 1062 5169 1068
rect 5134 1052 5137 1058
rect 5150 992 5153 1048
rect 5106 948 5110 951
rect 5134 942 5137 948
rect 5150 882 5153 888
rect 5094 878 5105 881
rect 5006 862 5009 868
rect 5054 862 5057 868
rect 5102 862 5105 878
rect 5158 872 5161 1058
rect 5174 991 5177 1148
rect 5202 1138 5206 1141
rect 5194 1068 5198 1071
rect 5166 988 5177 991
rect 5190 1022 5193 1058
rect 5166 882 5169 988
rect 5190 972 5193 1018
rect 5198 952 5201 1038
rect 5206 952 5209 1018
rect 5166 862 5169 878
rect 5206 872 5209 938
rect 5198 862 5201 868
rect 4902 858 4905 859
rect 5090 858 5094 861
rect 5130 858 5134 861
rect 5186 858 5190 861
rect 4998 852 5001 858
rect 5022 842 5025 858
rect 5034 848 5038 851
rect 4830 782 4833 818
rect 4814 778 4825 781
rect 4810 768 4814 771
rect 4822 752 4825 778
rect 4802 748 4806 751
rect 4874 748 4878 751
rect 4790 742 4793 748
rect 4790 722 4793 728
rect 4790 662 4793 698
rect 4798 612 4801 738
rect 4806 662 4809 668
rect 4830 652 4833 738
rect 4854 682 4857 688
rect 4870 662 4873 738
rect 4878 692 4881 698
rect 4894 662 4897 768
rect 4910 672 4913 678
rect 4902 662 4905 668
rect 4918 662 4921 838
rect 5046 832 5049 858
rect 4966 792 4969 808
rect 4926 732 4929 768
rect 4950 722 4953 758
rect 4936 703 4938 707
rect 4942 703 4945 707
rect 4949 703 4952 707
rect 4938 688 4942 691
rect 4958 672 4961 778
rect 5014 752 5017 828
rect 4978 748 4982 751
rect 5026 748 5030 751
rect 4966 742 4969 748
rect 5002 738 5006 741
rect 5002 728 5006 731
rect 4982 692 4985 718
rect 4990 682 4993 688
rect 4998 682 5001 698
rect 5006 672 5009 678
rect 5014 672 5017 748
rect 5038 732 5041 758
rect 5050 748 5054 751
rect 5074 748 5078 751
rect 5094 742 5097 758
rect 5062 722 5065 738
rect 5090 718 5094 721
rect 4962 658 4966 661
rect 5022 661 5025 718
rect 5062 672 5065 678
rect 5018 658 5025 661
rect 5042 658 5046 661
rect 5058 658 5062 661
rect 4806 552 4809 618
rect 4798 532 4801 538
rect 4790 452 4793 458
rect 4682 348 4686 351
rect 4746 348 4750 351
rect 4678 263 4681 308
rect 4694 262 4697 338
rect 4714 328 4721 331
rect 4702 312 4705 318
rect 4718 292 4721 328
rect 4714 278 4718 281
rect 4734 272 4737 318
rect 4750 292 4753 338
rect 4806 332 4809 458
rect 4814 342 4817 348
rect 4758 282 4761 288
rect 4766 272 4769 318
rect 4782 272 4785 278
rect 4678 258 4681 259
rect 4638 152 4641 168
rect 4642 138 4646 141
rect 4618 128 4622 131
rect 4602 118 4606 121
rect 4414 62 4417 68
rect 4422 62 4425 68
rect 4446 62 4449 68
rect 4454 62 4457 78
rect 4590 72 4593 78
rect 4482 68 4486 71
rect 4550 62 4553 68
rect 4622 62 4625 88
rect 4638 72 4641 138
rect 4654 92 4657 208
rect 4694 152 4697 258
rect 4710 162 4713 268
rect 4722 258 4726 261
rect 4742 261 4745 268
rect 4790 262 4793 328
rect 4806 302 4809 328
rect 4738 258 4745 261
rect 4774 242 4777 258
rect 4786 248 4790 251
rect 4806 232 4809 258
rect 4770 168 4774 171
rect 4710 152 4713 158
rect 4718 132 4721 168
rect 4750 152 4753 158
rect 4762 148 4766 151
rect 4734 142 4737 148
rect 4762 138 4766 141
rect 4766 92 4769 128
rect 4782 92 4785 168
rect 4750 72 4753 78
rect 4646 62 4649 68
rect 4782 62 4785 88
rect 4790 82 4793 168
rect 4798 82 4801 98
rect 4806 92 4809 218
rect 4814 152 4817 158
rect 4822 141 4825 618
rect 4870 592 4873 658
rect 4830 472 4833 528
rect 4894 512 4897 658
rect 5086 652 5089 718
rect 4946 648 4950 651
rect 4934 592 4937 648
rect 4982 632 4985 648
rect 5006 592 5009 648
rect 5030 642 5033 648
rect 5038 592 5041 648
rect 4982 552 4985 558
rect 4926 542 4929 548
rect 4934 532 4937 548
rect 4998 542 5001 558
rect 5030 552 5033 558
rect 4974 531 4977 538
rect 4974 528 4985 531
rect 4958 512 4961 528
rect 4936 503 4938 507
rect 4942 503 4945 507
rect 4949 503 4952 507
rect 4918 492 4921 498
rect 4890 478 4894 481
rect 4870 472 4873 478
rect 4834 459 4838 461
rect 4870 462 4873 468
rect 4918 462 4921 488
rect 4926 472 4929 478
rect 4958 472 4961 478
rect 4834 458 4841 459
rect 4878 422 4881 458
rect 4898 448 4902 451
rect 4958 392 4961 448
rect 4878 352 4881 358
rect 4870 322 4873 328
rect 4842 268 4846 271
rect 4830 262 4833 268
rect 4878 152 4881 348
rect 4886 342 4889 378
rect 4910 352 4913 378
rect 4974 362 4977 448
rect 4982 422 4985 528
rect 4998 462 5001 518
rect 5006 452 5009 528
rect 5022 522 5025 538
rect 5034 528 5038 531
rect 4898 348 4902 351
rect 4942 332 4945 348
rect 4950 322 4953 338
rect 4936 303 4938 307
rect 4942 303 4945 307
rect 4949 303 4952 307
rect 4906 258 4910 261
rect 4926 182 4929 268
rect 4966 192 4969 328
rect 4974 282 4977 358
rect 4982 352 4985 418
rect 4990 342 4993 368
rect 5014 352 5017 368
rect 5030 352 5033 508
rect 5038 492 5041 508
rect 5046 482 5049 648
rect 5070 632 5073 638
rect 5102 592 5105 848
rect 5126 802 5129 818
rect 5126 772 5129 778
rect 5114 748 5118 751
rect 5126 702 5129 768
rect 5114 658 5118 661
rect 5086 552 5089 558
rect 5062 542 5065 548
rect 5082 538 5086 541
rect 5054 522 5057 538
rect 5062 512 5065 538
rect 5094 512 5097 538
rect 5102 522 5105 548
rect 5046 472 5049 478
rect 5074 468 5078 471
rect 5050 458 5054 461
rect 5070 452 5073 458
rect 5078 452 5081 458
rect 5002 348 5006 351
rect 5074 348 5078 351
rect 4982 292 4985 338
rect 5014 292 5017 338
rect 5006 282 5009 288
rect 5038 282 5041 288
rect 5070 282 5073 338
rect 4974 272 4977 278
rect 4990 272 4993 278
rect 4974 252 4977 268
rect 5002 258 5006 261
rect 5018 258 5022 261
rect 4926 152 4929 178
rect 4990 172 4993 218
rect 4998 192 5001 258
rect 5070 252 5073 259
rect 5006 192 5009 248
rect 5086 222 5089 458
rect 4990 152 4993 168
rect 5014 152 5017 168
rect 5022 152 5025 198
rect 5030 172 5033 218
rect 5082 188 5086 191
rect 5030 152 5033 158
rect 5038 152 5041 158
rect 5062 152 5065 188
rect 4814 138 4825 141
rect 4814 92 4817 138
rect 4894 132 4897 147
rect 5022 142 5025 148
rect 5070 142 5073 148
rect 4954 118 4958 121
rect 4936 103 4938 107
rect 4942 103 4945 107
rect 4949 103 4952 107
rect 5094 92 5097 488
rect 5102 462 5105 468
rect 5110 462 5113 568
rect 5122 528 5126 531
rect 5126 462 5129 478
rect 5134 471 5137 858
rect 5158 822 5161 858
rect 5150 762 5153 768
rect 5158 752 5161 808
rect 5166 782 5169 788
rect 5158 732 5161 738
rect 5150 672 5153 678
rect 5166 672 5169 688
rect 5166 652 5169 658
rect 5150 552 5153 568
rect 5162 548 5166 551
rect 5174 542 5177 748
rect 5198 692 5201 738
rect 5182 582 5185 658
rect 5206 562 5209 568
rect 5190 552 5193 558
rect 5206 542 5209 558
rect 5162 538 5166 541
rect 5186 538 5190 541
rect 5142 522 5145 538
rect 5214 532 5217 1178
rect 5222 992 5225 1248
rect 5246 1152 5249 1258
rect 5262 1182 5265 1548
rect 5270 1482 5273 1528
rect 5270 1282 5273 1478
rect 5270 1152 5273 1259
rect 5286 1192 5289 1948
rect 5294 1742 5297 1758
rect 5302 1362 5305 1368
rect 5254 1142 5257 1148
rect 5270 1082 5273 1138
rect 5246 1062 5249 1068
rect 5278 992 5281 1018
rect 5238 882 5241 918
rect 5246 912 5249 948
rect 5262 932 5265 988
rect 5270 962 5273 988
rect 5286 952 5289 958
rect 5286 942 5289 948
rect 5238 862 5241 868
rect 5246 862 5249 868
rect 5238 851 5241 858
rect 5238 848 5249 851
rect 5222 752 5225 758
rect 5246 742 5249 848
rect 5254 772 5257 918
rect 5262 792 5265 898
rect 5278 792 5281 818
rect 5246 672 5249 738
rect 5266 728 5270 731
rect 5282 728 5286 731
rect 5246 552 5249 668
rect 5254 612 5257 658
rect 5158 492 5161 508
rect 5134 468 5145 471
rect 5102 442 5105 448
rect 5134 402 5137 458
rect 5142 422 5145 468
rect 5166 462 5169 488
rect 5158 412 5161 448
rect 5142 392 5145 408
rect 5166 362 5169 378
rect 5118 152 5121 338
rect 5134 332 5137 338
rect 5142 302 5145 348
rect 5130 288 5134 291
rect 5142 282 5145 298
rect 5158 292 5161 358
rect 5166 282 5169 338
rect 5174 282 5177 518
rect 5182 392 5185 528
rect 5198 452 5201 458
rect 5182 352 5185 358
rect 5190 342 5193 388
rect 5198 352 5201 418
rect 5182 292 5185 328
rect 5150 272 5153 278
rect 5166 272 5169 278
rect 5198 272 5201 348
rect 5214 332 5217 488
rect 5246 472 5249 548
rect 5270 542 5273 548
rect 5270 492 5273 528
rect 5262 482 5265 488
rect 5274 468 5278 471
rect 5222 462 5225 468
rect 5282 458 5286 461
rect 5238 392 5241 398
rect 5294 392 5297 598
rect 5282 388 5286 391
rect 5222 342 5225 358
rect 5250 348 5254 351
rect 5238 322 5241 348
rect 5262 342 5265 368
rect 5254 338 5262 341
rect 5206 312 5209 318
rect 5234 308 5241 311
rect 5238 292 5241 308
rect 5246 302 5249 338
rect 5210 288 5214 291
rect 5218 278 5222 281
rect 5234 268 5238 271
rect 5186 258 5190 261
rect 5142 212 5145 258
rect 5198 202 5201 268
rect 5222 222 5225 258
rect 5246 192 5249 278
rect 5254 272 5257 338
rect 5278 332 5281 338
rect 5270 282 5273 318
rect 5278 292 5281 308
rect 5286 302 5289 348
rect 5298 328 5302 331
rect 5282 278 5286 281
rect 5254 262 5257 268
rect 5278 192 5281 268
rect 5230 182 5233 188
rect 5130 148 5134 151
rect 5158 142 5161 178
rect 4834 88 4838 91
rect 4938 88 4942 91
rect 4826 78 4830 81
rect 4910 72 4913 78
rect 5038 72 5041 78
rect 5110 72 5113 138
rect 5174 132 5177 138
rect 5214 72 5217 78
rect 5106 68 5110 71
rect 4790 62 4793 68
rect 4014 58 4017 59
rect 4074 58 4078 61
rect 4378 58 4382 61
rect 4618 58 4622 61
rect 4714 58 4718 61
rect 4890 59 4894 62
rect 5002 59 5006 62
rect 3750 42 3753 48
rect 4086 42 4089 58
rect 4094 52 4097 58
rect 4454 52 4457 58
rect 4606 42 4609 58
rect 5022 52 5025 68
rect 5230 63 5233 158
rect 5246 152 5249 158
rect 5274 148 5278 151
rect 5262 132 5265 138
rect 5286 132 5289 258
rect 5282 68 5286 71
rect 5178 58 5182 61
rect 5230 58 5233 59
rect 4770 48 4774 51
rect 5170 48 5174 51
rect 5198 42 5201 48
rect 328 3 330 7
rect 334 3 337 7
rect 341 3 344 7
rect 1352 3 1354 7
rect 1358 3 1361 7
rect 1365 3 1368 7
rect 2230 -18 2233 8
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2397 3 2400 7
rect 3400 3 3402 7
rect 3406 3 3409 7
rect 3413 3 3416 7
rect 4424 3 4426 7
rect 4430 3 4433 7
rect 4437 3 4440 7
rect 4526 -18 4529 8
rect 2230 -22 2234 -18
rect 4526 -22 4530 -18
<< m3contact >>
rect 310 5098 314 5102
rect 850 5103 854 5107
rect 857 5103 861 5107
rect 510 5088 514 5092
rect 654 5088 658 5092
rect 702 5088 706 5092
rect 750 5088 754 5092
rect 814 5088 818 5092
rect 110 5078 114 5082
rect 150 5078 154 5082
rect 174 5078 178 5082
rect 294 5078 298 5082
rect 302 5078 306 5082
rect 318 5078 322 5082
rect 382 5078 386 5082
rect 38 5068 42 5072
rect 14 4988 18 4992
rect 54 5058 58 5062
rect 70 4938 74 4942
rect 558 5078 562 5082
rect 318 5068 322 5072
rect 118 5058 122 5062
rect 150 5058 154 5062
rect 158 5058 162 5062
rect 166 5058 170 5062
rect 190 5058 194 5062
rect 214 5059 218 5063
rect 126 5048 130 5052
rect 294 5048 298 5052
rect 222 5018 226 5022
rect 222 4968 226 4972
rect 278 4968 282 4972
rect 330 5003 334 5007
rect 337 5003 341 5007
rect 158 4958 162 4962
rect 142 4948 146 4952
rect 118 4938 122 4942
rect 102 4928 106 4932
rect 134 4918 138 4922
rect 126 4908 130 4912
rect 70 4898 74 4902
rect 110 4878 114 4882
rect 118 4868 122 4872
rect 190 4948 194 4952
rect 206 4948 210 4952
rect 262 4958 266 4962
rect 278 4958 282 4962
rect 286 4958 290 4962
rect 294 4958 298 4962
rect 382 5048 386 5052
rect 374 4998 378 5002
rect 446 5058 450 5062
rect 470 5058 474 5062
rect 462 5048 466 5052
rect 438 5038 442 5042
rect 454 5038 458 5042
rect 414 5018 418 5022
rect 406 5008 410 5012
rect 390 4958 394 4962
rect 238 4948 242 4952
rect 246 4938 250 4942
rect 270 4938 274 4942
rect 182 4928 186 4932
rect 166 4918 170 4922
rect 166 4888 170 4892
rect 214 4928 218 4932
rect 190 4918 194 4922
rect 190 4898 194 4902
rect 150 4858 154 4862
rect 38 4848 42 4852
rect 134 4848 138 4852
rect 158 4848 162 4852
rect 174 4848 178 4852
rect 150 4838 154 4842
rect 102 4828 106 4832
rect 118 4828 122 4832
rect 110 4818 114 4822
rect 62 4768 66 4772
rect 86 4758 90 4762
rect 126 4768 130 4772
rect 102 4748 106 4752
rect 126 4748 130 4752
rect 86 4738 90 4742
rect 6 4728 10 4732
rect 30 4718 34 4722
rect 62 4718 66 4722
rect 86 4718 90 4722
rect 54 4708 58 4712
rect 38 4698 42 4702
rect 46 4668 50 4672
rect 14 4568 18 4572
rect 22 4528 26 4532
rect 102 4668 106 4672
rect 94 4658 98 4662
rect 142 4758 146 4762
rect 158 4748 162 4752
rect 150 4738 154 4742
rect 158 4728 162 4732
rect 142 4718 146 4722
rect 134 4688 138 4692
rect 118 4668 122 4672
rect 150 4628 154 4632
rect 214 4818 218 4822
rect 206 4778 210 4782
rect 190 4768 194 4772
rect 230 4928 234 4932
rect 246 4898 250 4902
rect 254 4868 258 4872
rect 326 4948 330 4952
rect 310 4938 314 4942
rect 350 4948 354 4952
rect 366 4948 370 4952
rect 502 5048 506 5052
rect 494 5028 498 5032
rect 470 5018 474 5022
rect 486 5018 490 5022
rect 558 5058 562 5062
rect 582 5058 586 5062
rect 542 5048 546 5052
rect 598 5038 602 5042
rect 622 5038 626 5042
rect 606 5028 610 5032
rect 502 5008 506 5012
rect 534 5008 538 5012
rect 494 4998 498 5002
rect 454 4978 458 4982
rect 486 4968 490 4972
rect 422 4958 426 4962
rect 454 4958 458 4962
rect 470 4958 474 4962
rect 534 4988 538 4992
rect 502 4978 506 4982
rect 534 4978 538 4982
rect 358 4938 362 4942
rect 390 4938 394 4942
rect 446 4938 450 4942
rect 462 4938 466 4942
rect 342 4928 346 4932
rect 358 4928 362 4932
rect 414 4928 418 4932
rect 310 4888 314 4892
rect 350 4918 354 4922
rect 470 4918 474 4922
rect 302 4878 306 4882
rect 342 4878 346 4882
rect 310 4868 314 4872
rect 310 4858 314 4862
rect 254 4848 258 4852
rect 318 4848 322 4852
rect 222 4768 226 4772
rect 230 4768 234 4772
rect 198 4748 202 4752
rect 230 4738 234 4742
rect 262 4738 266 4742
rect 182 4638 186 4642
rect 158 4618 162 4622
rect 110 4598 114 4602
rect 110 4588 114 4592
rect 94 4568 98 4572
rect 214 4728 218 4732
rect 238 4718 242 4722
rect 222 4708 226 4712
rect 246 4698 250 4702
rect 206 4678 210 4682
rect 198 4668 202 4672
rect 206 4668 210 4672
rect 198 4658 202 4662
rect 214 4648 218 4652
rect 254 4648 258 4652
rect 198 4638 202 4642
rect 222 4638 226 4642
rect 230 4638 234 4642
rect 182 4578 186 4582
rect 134 4568 138 4572
rect 158 4568 162 4572
rect 174 4568 178 4572
rect 262 4578 266 4582
rect 230 4568 234 4572
rect 254 4568 258 4572
rect 46 4558 50 4562
rect 70 4558 74 4562
rect 94 4558 98 4562
rect 198 4558 202 4562
rect 54 4548 58 4552
rect 86 4548 90 4552
rect 54 4538 58 4542
rect 30 4508 34 4512
rect 6 4448 10 4452
rect 6 4438 10 4442
rect 22 4348 26 4352
rect 6 4298 10 4302
rect 30 4328 34 4332
rect 14 4288 18 4292
rect 22 4288 26 4292
rect 78 4518 82 4522
rect 54 4478 58 4482
rect 62 4468 66 4472
rect 278 4838 282 4842
rect 334 4838 338 4842
rect 342 4838 346 4842
rect 278 4778 282 4782
rect 330 4803 334 4807
rect 337 4803 341 4807
rect 334 4788 338 4792
rect 318 4768 322 4772
rect 318 4698 322 4702
rect 294 4668 298 4672
rect 278 4648 282 4652
rect 334 4648 338 4652
rect 390 4898 394 4902
rect 430 4908 434 4912
rect 462 4898 466 4902
rect 374 4878 378 4882
rect 390 4878 394 4882
rect 406 4878 410 4882
rect 430 4878 434 4882
rect 454 4878 458 4882
rect 422 4868 426 4872
rect 358 4858 362 4862
rect 518 4948 522 4952
rect 614 4998 618 5002
rect 606 4948 610 4952
rect 622 4968 626 4972
rect 798 5078 802 5082
rect 822 5078 826 5082
rect 910 5078 914 5082
rect 654 5068 658 5072
rect 694 5068 698 5072
rect 718 5068 722 5072
rect 742 5068 746 5072
rect 846 5068 850 5072
rect 662 5058 666 5062
rect 662 5028 666 5032
rect 558 4938 562 4942
rect 574 4938 578 4942
rect 518 4928 522 4932
rect 534 4928 538 4932
rect 542 4928 546 4932
rect 606 4928 610 4932
rect 566 4908 570 4912
rect 582 4898 586 4902
rect 774 5058 778 5062
rect 830 5058 834 5062
rect 734 5028 738 5032
rect 742 5028 746 5032
rect 734 4968 738 4972
rect 638 4938 642 4942
rect 646 4918 650 4922
rect 670 4918 674 4922
rect 542 4878 546 4882
rect 582 4878 586 4882
rect 646 4878 650 4882
rect 478 4868 482 4872
rect 374 4848 378 4852
rect 398 4848 402 4852
rect 406 4848 410 4852
rect 350 4628 354 4632
rect 318 4618 322 4622
rect 342 4618 346 4622
rect 330 4603 334 4607
rect 337 4603 341 4607
rect 294 4568 298 4572
rect 166 4548 170 4552
rect 270 4548 274 4552
rect 318 4558 322 4562
rect 366 4818 370 4822
rect 510 4858 514 4862
rect 526 4858 530 4862
rect 486 4848 490 4852
rect 502 4848 506 4852
rect 446 4838 450 4842
rect 398 4798 402 4802
rect 390 4768 394 4772
rect 438 4818 442 4822
rect 518 4838 522 4842
rect 526 4808 530 4812
rect 606 4858 610 4862
rect 622 4858 626 4862
rect 638 4858 642 4862
rect 574 4838 578 4842
rect 558 4818 562 4822
rect 638 4848 642 4852
rect 654 4828 658 4832
rect 614 4818 618 4822
rect 590 4798 594 4802
rect 606 4798 610 4802
rect 582 4788 586 4792
rect 438 4778 442 4782
rect 462 4778 466 4782
rect 486 4778 490 4782
rect 550 4778 554 4782
rect 566 4778 570 4782
rect 422 4768 426 4772
rect 470 4758 474 4762
rect 550 4758 554 4762
rect 430 4748 434 4752
rect 390 4738 394 4742
rect 438 4718 442 4722
rect 366 4688 370 4692
rect 366 4668 370 4672
rect 422 4658 426 4662
rect 406 4648 410 4652
rect 398 4638 402 4642
rect 390 4618 394 4622
rect 486 4738 490 4742
rect 502 4738 506 4742
rect 518 4738 522 4742
rect 462 4708 466 4712
rect 494 4698 498 4702
rect 542 4748 546 4752
rect 526 4688 530 4692
rect 534 4688 538 4692
rect 502 4678 506 4682
rect 582 4768 586 4772
rect 606 4778 610 4782
rect 670 4818 674 4822
rect 622 4788 626 4792
rect 662 4788 666 4792
rect 646 4778 650 4782
rect 662 4758 666 4762
rect 574 4738 578 4742
rect 598 4738 602 4742
rect 558 4728 562 4732
rect 590 4728 594 4732
rect 622 4728 626 4732
rect 646 4718 650 4722
rect 638 4708 642 4712
rect 606 4698 610 4702
rect 598 4688 602 4692
rect 606 4678 610 4682
rect 614 4668 618 4672
rect 638 4668 642 4672
rect 486 4658 490 4662
rect 542 4658 546 4662
rect 606 4658 610 4662
rect 478 4648 482 4652
rect 598 4648 602 4652
rect 582 4608 586 4612
rect 446 4598 450 4602
rect 526 4598 530 4602
rect 534 4598 538 4602
rect 358 4578 362 4582
rect 470 4568 474 4572
rect 446 4558 450 4562
rect 158 4538 162 4542
rect 126 4528 130 4532
rect 142 4518 146 4522
rect 110 4508 114 4512
rect 142 4488 146 4492
rect 166 4478 170 4482
rect 182 4468 186 4472
rect 102 4458 106 4462
rect 86 4448 90 4452
rect 118 4448 122 4452
rect 78 4388 82 4392
rect 110 4428 114 4432
rect 166 4458 170 4462
rect 206 4528 210 4532
rect 230 4538 234 4542
rect 270 4538 274 4542
rect 246 4528 250 4532
rect 230 4518 234 4522
rect 214 4508 218 4512
rect 246 4508 250 4512
rect 214 4478 218 4482
rect 190 4418 194 4422
rect 126 4408 130 4412
rect 190 4408 194 4412
rect 230 4458 234 4462
rect 278 4528 282 4532
rect 374 4538 378 4542
rect 382 4538 386 4542
rect 406 4538 410 4542
rect 366 4498 370 4502
rect 358 4478 362 4482
rect 262 4468 266 4472
rect 294 4468 298 4472
rect 326 4458 330 4462
rect 270 4448 274 4452
rect 142 4388 146 4392
rect 214 4388 218 4392
rect 230 4388 234 4392
rect 102 4368 106 4372
rect 174 4378 178 4382
rect 198 4378 202 4382
rect 214 4378 218 4382
rect 78 4358 82 4362
rect 102 4358 106 4362
rect 126 4358 130 4362
rect 142 4358 146 4362
rect 94 4338 98 4342
rect 118 4298 122 4302
rect 134 4298 138 4302
rect 158 4348 162 4352
rect 198 4348 202 4352
rect 150 4328 154 4332
rect 102 4278 106 4282
rect 62 4268 66 4272
rect 14 4248 18 4252
rect 102 4258 106 4262
rect 118 4248 122 4252
rect 78 4198 82 4202
rect 22 4168 26 4172
rect 102 4238 106 4242
rect 166 4298 170 4302
rect 246 4368 250 4372
rect 310 4448 314 4452
rect 278 4428 282 4432
rect 278 4418 282 4422
rect 430 4538 434 4542
rect 462 4538 466 4542
rect 510 4538 514 4542
rect 406 4528 410 4532
rect 446 4528 450 4532
rect 462 4518 466 4522
rect 390 4498 394 4502
rect 358 4458 362 4462
rect 342 4428 346 4432
rect 330 4403 334 4407
rect 337 4403 341 4407
rect 374 4418 378 4422
rect 366 4378 370 4382
rect 278 4368 282 4372
rect 302 4368 306 4372
rect 318 4368 322 4372
rect 214 4308 218 4312
rect 182 4278 186 4282
rect 214 4278 218 4282
rect 222 4278 226 4282
rect 230 4258 234 4262
rect 222 4248 226 4252
rect 150 4238 154 4242
rect 142 4198 146 4202
rect 254 4348 258 4352
rect 270 4348 274 4352
rect 302 4348 306 4352
rect 310 4278 314 4282
rect 246 4268 250 4272
rect 246 4258 250 4262
rect 302 4248 306 4252
rect 318 4248 322 4252
rect 230 4228 234 4232
rect 214 4188 218 4192
rect 142 4178 146 4182
rect 174 4178 178 4182
rect 110 4148 114 4152
rect 134 4148 138 4152
rect 94 4138 98 4142
rect 70 4108 74 4112
rect 86 4108 90 4112
rect 150 4168 154 4172
rect 238 4218 242 4222
rect 166 4148 170 4152
rect 214 4148 218 4152
rect 118 4128 122 4132
rect 166 4118 170 4122
rect 134 4108 138 4112
rect 134 4098 138 4102
rect 206 4128 210 4132
rect 206 4088 210 4092
rect 206 4078 210 4082
rect 230 4078 234 4082
rect 158 4068 162 4072
rect 182 4068 186 4072
rect 70 4058 74 4062
rect 46 4028 50 4032
rect 22 3988 26 3992
rect 6 3968 10 3972
rect 38 3958 42 3962
rect 6 3928 10 3932
rect 14 3868 18 3872
rect 62 4008 66 4012
rect 62 3948 66 3952
rect 198 4058 202 4062
rect 102 4048 106 4052
rect 150 4048 154 4052
rect 94 4038 98 4042
rect 102 4038 106 4042
rect 190 4038 194 4042
rect 86 3998 90 4002
rect 86 3978 90 3982
rect 54 3938 58 3942
rect 70 3938 74 3942
rect 62 3918 66 3922
rect 62 3908 66 3912
rect 54 3898 58 3902
rect 134 3998 138 4002
rect 174 3998 178 4002
rect 126 3958 130 3962
rect 174 3978 178 3982
rect 150 3958 154 3962
rect 110 3928 114 3932
rect 86 3868 90 3872
rect 22 3838 26 3842
rect 38 3838 42 3842
rect 126 3878 130 3882
rect 126 3858 130 3862
rect 110 3848 114 3852
rect 78 3838 82 3842
rect 70 3828 74 3832
rect 102 3828 106 3832
rect 126 3838 130 3842
rect 134 3838 138 3842
rect 70 3808 74 3812
rect 30 3778 34 3782
rect 38 3768 42 3772
rect 62 3768 66 3772
rect 54 3748 58 3752
rect 38 3698 42 3702
rect 62 3698 66 3702
rect 14 3678 18 3682
rect 118 3778 122 3782
rect 78 3768 82 3772
rect 102 3768 106 3772
rect 86 3758 90 3762
rect 86 3748 90 3752
rect 102 3748 106 3752
rect 110 3738 114 3742
rect 6 3668 10 3672
rect 102 3668 106 3672
rect 38 3658 42 3662
rect 62 3658 66 3662
rect 86 3658 90 3662
rect 14 3648 18 3652
rect 54 3648 58 3652
rect 78 3648 82 3652
rect 14 3518 18 3522
rect 126 3768 130 3772
rect 158 3938 162 3942
rect 182 3898 186 3902
rect 150 3888 154 3892
rect 166 3888 170 3892
rect 174 3888 178 3892
rect 158 3878 162 3882
rect 206 3988 210 3992
rect 198 3958 202 3962
rect 198 3938 202 3942
rect 230 4018 234 4022
rect 494 4488 498 4492
rect 518 4528 522 4532
rect 438 4478 442 4482
rect 446 4468 450 4472
rect 494 4468 498 4472
rect 406 4458 410 4462
rect 438 4458 442 4462
rect 486 4458 490 4462
rect 398 4448 402 4452
rect 470 4448 474 4452
rect 406 4428 410 4432
rect 414 4398 418 4402
rect 390 4368 394 4372
rect 342 4358 346 4362
rect 358 4358 362 4362
rect 374 4358 378 4362
rect 334 4348 338 4352
rect 366 4348 370 4352
rect 390 4348 394 4352
rect 406 4348 410 4352
rect 494 4398 498 4402
rect 494 4378 498 4382
rect 462 4348 466 4352
rect 366 4328 370 4332
rect 470 4328 474 4332
rect 494 4328 498 4332
rect 598 4578 602 4582
rect 582 4568 586 4572
rect 566 4558 570 4562
rect 542 4548 546 4552
rect 550 4538 554 4542
rect 582 4538 586 4542
rect 542 4528 546 4532
rect 526 4508 530 4512
rect 518 4458 522 4462
rect 526 4448 530 4452
rect 534 4448 538 4452
rect 534 4428 538 4432
rect 526 4368 530 4372
rect 462 4318 466 4322
rect 510 4318 514 4322
rect 494 4308 498 4312
rect 486 4298 490 4302
rect 374 4278 378 4282
rect 382 4278 386 4282
rect 414 4278 418 4282
rect 462 4278 466 4282
rect 366 4268 370 4272
rect 390 4268 394 4272
rect 414 4268 418 4272
rect 374 4258 378 4262
rect 358 4248 362 4252
rect 294 4228 298 4232
rect 326 4228 330 4232
rect 262 4178 266 4182
rect 246 4148 250 4152
rect 286 4158 290 4162
rect 330 4203 334 4207
rect 337 4203 341 4207
rect 382 4238 386 4242
rect 406 4228 410 4232
rect 390 4208 394 4212
rect 366 4188 370 4192
rect 326 4168 330 4172
rect 310 4148 314 4152
rect 270 4128 274 4132
rect 278 4128 282 4132
rect 318 4098 322 4102
rect 254 4068 258 4072
rect 286 4058 290 4062
rect 302 4058 306 4062
rect 254 4048 258 4052
rect 270 4038 274 4042
rect 254 4008 258 4012
rect 238 3998 242 4002
rect 222 3978 226 3982
rect 230 3958 234 3962
rect 350 4128 354 4132
rect 390 4178 394 4182
rect 430 4268 434 4272
rect 446 4268 450 4272
rect 422 4258 426 4262
rect 422 4238 426 4242
rect 374 4148 378 4152
rect 390 4148 394 4152
rect 382 4118 386 4122
rect 390 4088 394 4092
rect 414 4078 418 4082
rect 358 4068 362 4072
rect 342 4058 346 4062
rect 374 4048 378 4052
rect 310 4038 314 4042
rect 286 3998 290 4002
rect 630 4658 634 4662
rect 622 4638 626 4642
rect 614 4628 618 4632
rect 622 4608 626 4612
rect 670 4738 674 4742
rect 662 4698 666 4702
rect 654 4658 658 4662
rect 718 4918 722 4922
rect 702 4908 706 4912
rect 694 4878 698 4882
rect 702 4858 706 4862
rect 694 4848 698 4852
rect 702 4838 706 4842
rect 710 4788 714 4792
rect 694 4708 698 4712
rect 734 4928 738 4932
rect 870 5058 874 5062
rect 790 5048 794 5052
rect 758 5038 762 5042
rect 822 5038 826 5042
rect 894 4998 898 5002
rect 774 4978 778 4982
rect 862 4978 866 4982
rect 894 4978 898 4982
rect 838 4968 842 4972
rect 846 4968 850 4972
rect 886 4968 890 4972
rect 902 4968 906 4972
rect 766 4938 770 4942
rect 790 4938 794 4942
rect 782 4928 786 4932
rect 750 4908 754 4912
rect 782 4918 786 4922
rect 766 4908 770 4912
rect 814 4958 818 4962
rect 830 4958 834 4962
rect 934 5048 938 5052
rect 1054 5058 1058 5062
rect 1126 5088 1130 5092
rect 1118 5068 1122 5072
rect 1134 5068 1138 5072
rect 1190 5068 1194 5072
rect 1182 5058 1186 5062
rect 1070 5048 1074 5052
rect 1078 5038 1082 5042
rect 1094 5038 1098 5042
rect 942 5028 946 5032
rect 1038 5028 1042 5032
rect 926 5018 930 5022
rect 942 5008 946 5012
rect 1046 5008 1050 5012
rect 942 4998 946 5002
rect 934 4958 938 4962
rect 918 4948 922 4952
rect 830 4938 834 4942
rect 838 4928 842 4932
rect 798 4888 802 4892
rect 822 4878 826 4882
rect 734 4838 738 4842
rect 774 4858 778 4862
rect 790 4858 794 4862
rect 806 4858 810 4862
rect 766 4828 770 4832
rect 774 4828 778 4832
rect 750 4758 754 4762
rect 742 4738 746 4742
rect 734 4728 738 4732
rect 750 4728 754 4732
rect 726 4718 730 4722
rect 774 4708 778 4712
rect 806 4848 810 4852
rect 850 4903 854 4907
rect 857 4903 861 4907
rect 934 4928 938 4932
rect 926 4918 930 4922
rect 958 4988 962 4992
rect 950 4968 954 4972
rect 974 4968 978 4972
rect 1006 4968 1010 4972
rect 966 4958 970 4962
rect 950 4898 954 4902
rect 926 4878 930 4882
rect 846 4848 850 4852
rect 838 4828 842 4832
rect 814 4808 818 4812
rect 806 4778 810 4782
rect 830 4768 834 4772
rect 814 4758 818 4762
rect 862 4858 866 4862
rect 870 4858 874 4862
rect 894 4858 898 4862
rect 950 4858 954 4862
rect 886 4838 890 4842
rect 862 4828 866 4832
rect 878 4818 882 4822
rect 958 4798 962 4802
rect 926 4788 930 4792
rect 950 4788 954 4792
rect 918 4768 922 4772
rect 854 4758 858 4762
rect 958 4778 962 4782
rect 846 4748 850 4752
rect 798 4738 802 4742
rect 814 4738 818 4742
rect 830 4738 834 4742
rect 854 4738 858 4742
rect 902 4738 906 4742
rect 918 4738 922 4742
rect 886 4728 890 4732
rect 902 4728 906 4732
rect 790 4718 794 4722
rect 822 4718 826 4722
rect 862 4718 866 4722
rect 902 4708 906 4712
rect 734 4678 738 4682
rect 734 4668 738 4672
rect 758 4668 762 4672
rect 850 4703 854 4707
rect 857 4703 861 4707
rect 822 4688 826 4692
rect 886 4688 890 4692
rect 870 4678 874 4682
rect 822 4668 826 4672
rect 694 4658 698 4662
rect 718 4658 722 4662
rect 750 4658 754 4662
rect 686 4638 690 4642
rect 662 4628 666 4632
rect 654 4578 658 4582
rect 614 4558 618 4562
rect 678 4568 682 4572
rect 694 4628 698 4632
rect 702 4628 706 4632
rect 758 4628 762 4632
rect 742 4568 746 4572
rect 702 4558 706 4562
rect 670 4548 674 4552
rect 590 4518 594 4522
rect 598 4508 602 4512
rect 566 4498 570 4502
rect 590 4498 594 4502
rect 574 4488 578 4492
rect 582 4478 586 4482
rect 598 4478 602 4482
rect 550 4468 554 4472
rect 566 4448 570 4452
rect 582 4448 586 4452
rect 550 4418 554 4422
rect 550 4398 554 4402
rect 574 4358 578 4362
rect 534 4288 538 4292
rect 478 4268 482 4272
rect 526 4268 530 4272
rect 542 4268 546 4272
rect 486 4258 490 4262
rect 614 4458 618 4462
rect 606 4398 610 4402
rect 662 4538 666 4542
rect 638 4518 642 4522
rect 638 4508 642 4512
rect 630 4498 634 4502
rect 630 4488 634 4492
rect 678 4498 682 4502
rect 670 4488 674 4492
rect 654 4458 658 4462
rect 638 4448 642 4452
rect 710 4548 714 4552
rect 766 4618 770 4622
rect 694 4528 698 4532
rect 830 4658 834 4662
rect 870 4658 874 4662
rect 822 4638 826 4642
rect 798 4558 802 4562
rect 806 4558 810 4562
rect 782 4548 786 4552
rect 790 4548 794 4552
rect 782 4518 786 4522
rect 702 4468 706 4472
rect 718 4468 722 4472
rect 766 4468 770 4472
rect 846 4638 850 4642
rect 854 4628 858 4632
rect 814 4538 818 4542
rect 854 4538 858 4542
rect 798 4488 802 4492
rect 806 4478 810 4482
rect 798 4468 802 4472
rect 702 4458 706 4462
rect 774 4458 778 4462
rect 710 4448 714 4452
rect 838 4528 842 4532
rect 822 4518 826 4522
rect 830 4508 834 4512
rect 830 4468 834 4472
rect 822 4458 826 4462
rect 766 4448 770 4452
rect 814 4448 818 4452
rect 686 4438 690 4442
rect 718 4438 722 4442
rect 646 4428 650 4432
rect 662 4418 666 4422
rect 622 4378 626 4382
rect 750 4428 754 4432
rect 702 4398 706 4402
rect 726 4398 730 4402
rect 702 4368 706 4372
rect 606 4358 610 4362
rect 622 4358 626 4362
rect 638 4358 642 4362
rect 662 4358 666 4362
rect 606 4348 610 4352
rect 582 4338 586 4342
rect 598 4338 602 4342
rect 566 4328 570 4332
rect 646 4348 650 4352
rect 598 4318 602 4322
rect 558 4308 562 4312
rect 590 4308 594 4312
rect 438 4248 442 4252
rect 534 4248 538 4252
rect 478 4218 482 4222
rect 494 4208 498 4212
rect 470 4198 474 4202
rect 550 4208 554 4212
rect 566 4278 570 4282
rect 590 4278 594 4282
rect 606 4278 610 4282
rect 566 4238 570 4242
rect 566 4228 570 4232
rect 590 4268 594 4272
rect 742 4358 746 4362
rect 686 4338 690 4342
rect 694 4328 698 4332
rect 710 4328 714 4332
rect 662 4298 666 4302
rect 662 4288 666 4292
rect 670 4268 674 4272
rect 830 4438 834 4442
rect 822 4408 826 4412
rect 806 4358 810 4362
rect 774 4348 778 4352
rect 734 4318 738 4322
rect 758 4318 762 4322
rect 686 4298 690 4302
rect 694 4278 698 4282
rect 702 4278 706 4282
rect 766 4308 770 4312
rect 726 4288 730 4292
rect 734 4288 738 4292
rect 710 4268 714 4272
rect 726 4268 730 4272
rect 606 4258 610 4262
rect 686 4258 690 4262
rect 622 4238 626 4242
rect 582 4208 586 4212
rect 558 4188 562 4192
rect 718 4258 722 4262
rect 742 4278 746 4282
rect 758 4268 762 4272
rect 734 4258 738 4262
rect 710 4218 714 4222
rect 718 4208 722 4212
rect 702 4178 706 4182
rect 430 4168 434 4172
rect 478 4168 482 4172
rect 598 4168 602 4172
rect 646 4168 650 4172
rect 502 4158 506 4162
rect 494 4148 498 4152
rect 478 4138 482 4142
rect 438 4098 442 4102
rect 462 4088 466 4092
rect 422 4058 426 4062
rect 430 4058 434 4062
rect 414 4048 418 4052
rect 454 4058 458 4062
rect 478 4058 482 4062
rect 438 4038 442 4042
rect 470 4038 474 4042
rect 486 4038 490 4042
rect 398 4018 402 4022
rect 406 4018 410 4022
rect 330 4003 334 4007
rect 337 4003 341 4007
rect 318 3998 322 4002
rect 454 4028 458 4032
rect 438 4008 442 4012
rect 326 3988 330 3992
rect 406 3988 410 3992
rect 278 3958 282 3962
rect 222 3948 226 3952
rect 254 3938 258 3942
rect 222 3918 226 3922
rect 294 3958 298 3962
rect 318 3958 322 3962
rect 302 3948 306 3952
rect 286 3938 290 3942
rect 230 3878 234 3882
rect 190 3868 194 3872
rect 286 3868 290 3872
rect 374 3978 378 3982
rect 366 3968 370 3972
rect 414 3968 418 3972
rect 510 4138 514 4142
rect 518 4138 522 4142
rect 574 4158 578 4162
rect 534 4148 538 4152
rect 582 4138 586 4142
rect 502 4128 506 4132
rect 526 4128 530 4132
rect 550 4128 554 4132
rect 542 4118 546 4122
rect 518 4108 522 4112
rect 630 4158 634 4162
rect 678 4168 682 4172
rect 702 4168 706 4172
rect 614 4148 618 4152
rect 654 4148 658 4152
rect 670 4148 674 4152
rect 622 4138 626 4142
rect 686 4138 690 4142
rect 574 4088 578 4092
rect 542 4078 546 4082
rect 518 4058 522 4062
rect 534 4058 538 4062
rect 550 4058 554 4062
rect 558 4058 562 4062
rect 574 4058 578 4062
rect 542 4038 546 4042
rect 510 4018 514 4022
rect 502 4008 506 4012
rect 494 3978 498 3982
rect 462 3968 466 3972
rect 630 4128 634 4132
rect 646 4128 650 4132
rect 606 4088 610 4092
rect 694 4108 698 4112
rect 710 4098 714 4102
rect 726 4158 730 4162
rect 798 4348 802 4352
rect 850 4503 854 4507
rect 857 4503 861 4507
rect 894 4588 898 4592
rect 902 4518 906 4522
rect 854 4488 858 4492
rect 894 4468 898 4472
rect 862 4458 866 4462
rect 870 4448 874 4452
rect 886 4438 890 4442
rect 894 4438 898 4442
rect 862 4418 866 4422
rect 878 4348 882 4352
rect 830 4338 834 4342
rect 798 4328 802 4332
rect 814 4328 818 4332
rect 782 4288 786 4292
rect 774 4258 778 4262
rect 782 4258 786 4262
rect 806 4258 810 4262
rect 814 4228 818 4232
rect 814 4208 818 4212
rect 814 4198 818 4202
rect 758 4148 762 4152
rect 766 4148 770 4152
rect 750 4138 754 4142
rect 850 4303 854 4307
rect 857 4303 861 4307
rect 870 4288 874 4292
rect 838 4268 842 4272
rect 862 4268 866 4272
rect 870 4258 874 4262
rect 870 4238 874 4242
rect 854 4218 858 4222
rect 878 4208 882 4212
rect 942 4718 946 4722
rect 990 4948 994 4952
rect 1062 4948 1066 4952
rect 1014 4938 1018 4942
rect 982 4928 986 4932
rect 1006 4888 1010 4892
rect 982 4878 986 4882
rect 1022 4868 1026 4872
rect 1006 4858 1010 4862
rect 974 4838 978 4842
rect 1030 4838 1034 4842
rect 1166 4948 1170 4952
rect 1134 4938 1138 4942
rect 1174 4938 1178 4942
rect 1054 4928 1058 4932
rect 1078 4918 1082 4922
rect 1230 5088 1234 5092
rect 1238 5068 1242 5072
rect 1270 5068 1274 5072
rect 1406 5068 1410 5072
rect 1270 5058 1274 5062
rect 1230 5048 1234 5052
rect 1246 5048 1250 5052
rect 1150 4888 1154 4892
rect 1182 4888 1186 4892
rect 1054 4878 1058 4882
rect 1086 4868 1090 4872
rect 1182 4868 1186 4872
rect 1086 4858 1090 4862
rect 1078 4848 1082 4852
rect 1102 4848 1106 4852
rect 1038 4828 1042 4832
rect 1094 4828 1098 4832
rect 982 4778 986 4782
rect 1014 4768 1018 4772
rect 1038 4768 1042 4772
rect 990 4748 994 4752
rect 1038 4748 1042 4752
rect 974 4728 978 4732
rect 926 4698 930 4702
rect 934 4698 938 4702
rect 990 4698 994 4702
rect 942 4688 946 4692
rect 966 4688 970 4692
rect 950 4678 954 4682
rect 918 4668 922 4672
rect 934 4658 938 4662
rect 934 4618 938 4622
rect 926 4558 930 4562
rect 950 4558 954 4562
rect 1022 4718 1026 4722
rect 1134 4848 1138 4852
rect 1158 4848 1162 4852
rect 1174 4858 1178 4862
rect 1222 4958 1226 4962
rect 1254 4998 1258 5002
rect 1262 4968 1266 4972
rect 1334 5038 1338 5042
rect 1278 4998 1282 5002
rect 1270 4958 1274 4962
rect 1294 4968 1298 4972
rect 1354 5003 1358 5007
rect 1361 5003 1365 5007
rect 1350 4958 1354 4962
rect 1222 4948 1226 4952
rect 1302 4948 1306 4952
rect 1342 4948 1346 4952
rect 1222 4928 1226 4932
rect 1254 4928 1258 4932
rect 1270 4928 1274 4932
rect 1198 4918 1202 4922
rect 1214 4878 1218 4882
rect 1230 4878 1234 4882
rect 1238 4868 1242 4872
rect 1254 4868 1258 4872
rect 1230 4858 1234 4862
rect 1182 4838 1186 4842
rect 1126 4828 1130 4832
rect 1166 4828 1170 4832
rect 1118 4808 1122 4812
rect 1126 4788 1130 4792
rect 1158 4778 1162 4782
rect 1182 4778 1186 4782
rect 1158 4768 1162 4772
rect 1102 4758 1106 4762
rect 1094 4748 1098 4752
rect 1110 4748 1114 4752
rect 1142 4748 1146 4752
rect 1054 4728 1058 4732
rect 1070 4728 1074 4732
rect 1046 4708 1050 4712
rect 1054 4708 1058 4712
rect 1006 4698 1010 4702
rect 998 4678 1002 4682
rect 1006 4668 1010 4672
rect 982 4648 986 4652
rect 1046 4658 1050 4662
rect 1038 4648 1042 4652
rect 1014 4618 1018 4622
rect 1022 4618 1026 4622
rect 1110 4738 1114 4742
rect 1142 4738 1146 4742
rect 1102 4728 1106 4732
rect 1134 4728 1138 4732
rect 1158 4738 1162 4742
rect 1150 4718 1154 4722
rect 1086 4698 1090 4702
rect 1102 4698 1106 4702
rect 1078 4688 1082 4692
rect 1078 4658 1082 4662
rect 1094 4658 1098 4662
rect 1102 4648 1106 4652
rect 1062 4638 1066 4642
rect 1054 4628 1058 4632
rect 1078 4628 1082 4632
rect 1030 4608 1034 4612
rect 982 4578 986 4582
rect 974 4538 978 4542
rect 918 4528 922 4532
rect 910 4498 914 4502
rect 934 4498 938 4502
rect 934 4458 938 4462
rect 918 4398 922 4402
rect 1046 4578 1050 4582
rect 1038 4558 1042 4562
rect 1126 4698 1130 4702
rect 1134 4698 1138 4702
rect 1158 4688 1162 4692
rect 1134 4678 1138 4682
rect 1142 4678 1146 4682
rect 1246 4828 1250 4832
rect 1238 4768 1242 4772
rect 1198 4758 1202 4762
rect 1246 4748 1250 4752
rect 1174 4738 1178 4742
rect 1182 4728 1186 4732
rect 1190 4728 1194 4732
rect 1206 4738 1210 4742
rect 1182 4678 1186 4682
rect 1190 4678 1194 4682
rect 1198 4678 1202 4682
rect 1126 4648 1130 4652
rect 1158 4648 1162 4652
rect 1118 4588 1122 4592
rect 1110 4578 1114 4582
rect 1118 4578 1122 4582
rect 1078 4568 1082 4572
rect 1102 4568 1106 4572
rect 1014 4538 1018 4542
rect 1134 4588 1138 4592
rect 1118 4558 1122 4562
rect 1038 4538 1042 4542
rect 1070 4538 1074 4542
rect 1078 4528 1082 4532
rect 990 4518 994 4522
rect 1014 4508 1018 4512
rect 982 4478 986 4482
rect 950 4468 954 4472
rect 966 4468 970 4472
rect 982 4468 986 4472
rect 958 4448 962 4452
rect 998 4448 1002 4452
rect 950 4428 954 4432
rect 1006 4398 1010 4402
rect 950 4388 954 4392
rect 982 4388 986 4392
rect 918 4368 922 4372
rect 974 4368 978 4372
rect 934 4338 938 4342
rect 966 4348 970 4352
rect 958 4338 962 4342
rect 974 4338 978 4342
rect 1070 4468 1074 4472
rect 1030 4458 1034 4462
rect 1046 4458 1050 4462
rect 1014 4368 1018 4372
rect 1030 4368 1034 4372
rect 1006 4348 1010 4352
rect 1142 4558 1146 4562
rect 1166 4558 1170 4562
rect 1182 4568 1186 4572
rect 1230 4728 1234 4732
rect 1222 4718 1226 4722
rect 1222 4668 1226 4672
rect 1198 4658 1202 4662
rect 1190 4558 1194 4562
rect 1134 4538 1138 4542
rect 1190 4538 1194 4542
rect 1246 4708 1250 4712
rect 1238 4698 1242 4702
rect 1246 4678 1250 4682
rect 1246 4648 1250 4652
rect 1230 4638 1234 4642
rect 1278 4818 1282 4822
rect 1382 5028 1386 5032
rect 1874 5103 1878 5107
rect 1881 5103 1885 5107
rect 1662 5098 1666 5102
rect 1734 5078 1738 5082
rect 1822 5078 1826 5082
rect 1542 5068 1546 5072
rect 1590 5068 1594 5072
rect 1662 5068 1666 5072
rect 1734 5068 1738 5072
rect 1478 5058 1482 5062
rect 1454 4968 1458 4972
rect 1390 4958 1394 4962
rect 1374 4928 1378 4932
rect 1342 4898 1346 4902
rect 1350 4888 1354 4892
rect 1406 4948 1410 4952
rect 1438 4948 1442 4952
rect 1470 4948 1474 4952
rect 1398 4938 1402 4942
rect 1406 4898 1410 4902
rect 1430 4928 1434 4932
rect 1422 4898 1426 4902
rect 1574 5058 1578 5062
rect 1654 5008 1658 5012
rect 1654 4998 1658 5002
rect 1542 4968 1546 4972
rect 1590 4958 1594 4962
rect 1710 4958 1714 4962
rect 1518 4948 1522 4952
rect 1726 4948 1730 4952
rect 1494 4938 1498 4942
rect 1486 4888 1490 4892
rect 1654 4938 1658 4942
rect 1614 4928 1618 4932
rect 1414 4878 1418 4882
rect 1470 4878 1474 4882
rect 1798 5058 1802 5062
rect 1846 4998 1850 5002
rect 2890 5103 2894 5107
rect 2897 5103 2901 5107
rect 3922 5103 3926 5107
rect 3929 5103 3933 5107
rect 4938 5103 4942 5107
rect 4945 5103 4949 5107
rect 2310 5088 2314 5092
rect 2454 5088 2458 5092
rect 2526 5088 2530 5092
rect 2614 5088 2618 5092
rect 4150 5088 4154 5092
rect 4238 5088 4242 5092
rect 4486 5088 4490 5092
rect 1934 5078 1938 5082
rect 2126 5078 2130 5082
rect 2430 5078 2434 5082
rect 2462 5078 2466 5082
rect 4502 5078 4506 5082
rect 5014 5078 5018 5082
rect 5022 5078 5026 5082
rect 1982 5068 1986 5072
rect 2246 5068 2250 5072
rect 2406 5068 2410 5072
rect 2446 5068 2450 5072
rect 2062 5058 2066 5062
rect 1910 5018 1914 5022
rect 1958 5018 1962 5022
rect 1942 4998 1946 5002
rect 1926 4958 1930 4962
rect 1934 4958 1938 4962
rect 1894 4938 1898 4942
rect 1862 4928 1866 4932
rect 1902 4928 1906 4932
rect 1854 4918 1858 4922
rect 1870 4918 1874 4922
rect 1806 4908 1810 4912
rect 1726 4888 1730 4892
rect 1742 4888 1746 4892
rect 1382 4868 1386 4872
rect 1438 4866 1442 4870
rect 1494 4868 1498 4872
rect 1662 4868 1666 4872
rect 1454 4858 1458 4862
rect 1502 4858 1506 4862
rect 1574 4858 1578 4862
rect 1354 4803 1358 4807
rect 1361 4803 1365 4807
rect 1430 4818 1434 4822
rect 1358 4788 1362 4792
rect 1406 4788 1410 4792
rect 1334 4768 1338 4772
rect 1278 4758 1282 4762
rect 1310 4758 1314 4762
rect 1270 4748 1274 4752
rect 1302 4748 1306 4752
rect 1270 4728 1274 4732
rect 1270 4688 1274 4692
rect 1302 4728 1306 4732
rect 1286 4698 1290 4702
rect 1310 4698 1314 4702
rect 1318 4668 1322 4672
rect 1270 4628 1274 4632
rect 1254 4608 1258 4612
rect 1310 4658 1314 4662
rect 1326 4648 1330 4652
rect 1302 4638 1306 4642
rect 1310 4618 1314 4622
rect 1318 4618 1322 4622
rect 1294 4608 1298 4612
rect 1230 4588 1234 4592
rect 1238 4568 1242 4572
rect 1302 4578 1306 4582
rect 1302 4568 1306 4572
rect 1206 4558 1210 4562
rect 1214 4558 1218 4562
rect 1310 4558 1314 4562
rect 1214 4548 1218 4552
rect 1254 4548 1258 4552
rect 1270 4548 1274 4552
rect 1206 4538 1210 4542
rect 1238 4538 1242 4542
rect 1174 4528 1178 4532
rect 1166 4518 1170 4522
rect 1126 4488 1130 4492
rect 1142 4478 1146 4482
rect 1102 4458 1106 4462
rect 1118 4458 1122 4462
rect 1094 4448 1098 4452
rect 1086 4438 1090 4442
rect 1102 4438 1106 4442
rect 1102 4428 1106 4432
rect 1094 4388 1098 4392
rect 1046 4348 1050 4352
rect 1158 4508 1162 4512
rect 1182 4518 1186 4522
rect 1174 4508 1178 4512
rect 1158 4468 1162 4472
rect 1174 4468 1178 4472
rect 1030 4338 1034 4342
rect 1134 4378 1138 4382
rect 1238 4528 1242 4532
rect 1262 4538 1266 4542
rect 1214 4518 1218 4522
rect 1222 4478 1226 4482
rect 1222 4458 1226 4462
rect 1182 4448 1186 4452
rect 1214 4448 1218 4452
rect 1270 4518 1274 4522
rect 1278 4518 1282 4522
rect 1262 4488 1266 4492
rect 1246 4468 1250 4472
rect 1254 4458 1258 4462
rect 1342 4728 1346 4732
rect 1366 4778 1370 4782
rect 1390 4768 1394 4772
rect 1382 4738 1386 4742
rect 1342 4688 1346 4692
rect 1366 4688 1370 4692
rect 1406 4668 1410 4672
rect 1422 4668 1426 4672
rect 1398 4658 1402 4662
rect 1406 4658 1410 4662
rect 1334 4638 1338 4642
rect 1366 4638 1370 4642
rect 1366 4618 1370 4622
rect 1354 4603 1358 4607
rect 1361 4603 1365 4607
rect 1382 4588 1386 4592
rect 1350 4548 1354 4552
rect 1366 4548 1370 4552
rect 1334 4528 1338 4532
rect 1342 4518 1346 4522
rect 1326 4498 1330 4502
rect 1326 4488 1330 4492
rect 1382 4538 1386 4542
rect 1358 4528 1362 4532
rect 1406 4638 1410 4642
rect 1414 4628 1418 4632
rect 1862 4908 1866 4912
rect 1874 4903 1878 4907
rect 1881 4903 1885 4907
rect 1910 4888 1914 4892
rect 1742 4858 1746 4862
rect 1774 4858 1778 4862
rect 1862 4858 1866 4862
rect 1886 4858 1890 4862
rect 1654 4818 1658 4822
rect 1518 4778 1522 4782
rect 1574 4758 1578 4762
rect 1486 4748 1490 4752
rect 1526 4748 1530 4752
rect 1582 4748 1586 4752
rect 1614 4748 1618 4752
rect 1446 4738 1450 4742
rect 1462 4728 1466 4732
rect 1438 4698 1442 4702
rect 1462 4688 1466 4692
rect 1470 4688 1474 4692
rect 1438 4638 1442 4642
rect 1382 4518 1386 4522
rect 1398 4518 1402 4522
rect 1406 4518 1410 4522
rect 1358 4488 1362 4492
rect 1390 4488 1394 4492
rect 1286 4478 1290 4482
rect 1294 4478 1298 4482
rect 1310 4478 1314 4482
rect 1350 4478 1354 4482
rect 1374 4478 1378 4482
rect 1286 4468 1290 4472
rect 1294 4468 1298 4472
rect 1286 4448 1290 4452
rect 1254 4438 1258 4442
rect 1246 4408 1250 4412
rect 1302 4408 1306 4412
rect 1230 4398 1234 4402
rect 1150 4348 1154 4352
rect 1158 4348 1162 4352
rect 974 4328 978 4332
rect 1030 4328 1034 4332
rect 1110 4328 1114 4332
rect 1134 4328 1138 4332
rect 942 4318 946 4322
rect 958 4318 962 4322
rect 982 4278 986 4282
rect 990 4268 994 4272
rect 926 4258 930 4262
rect 958 4258 962 4262
rect 1054 4308 1058 4312
rect 1046 4288 1050 4292
rect 1022 4268 1026 4272
rect 950 4248 954 4252
rect 1014 4248 1018 4252
rect 1022 4248 1026 4252
rect 950 4238 954 4242
rect 918 4188 922 4192
rect 894 4168 898 4172
rect 910 4168 914 4172
rect 974 4168 978 4172
rect 830 4148 834 4152
rect 838 4148 842 4152
rect 822 4128 826 4132
rect 790 4118 794 4122
rect 798 4118 802 4122
rect 678 4088 682 4092
rect 766 4088 770 4092
rect 678 4068 682 4072
rect 702 4068 706 4072
rect 614 4058 618 4062
rect 646 4058 650 4062
rect 670 4058 674 4062
rect 518 3988 522 3992
rect 614 3988 618 3992
rect 526 3978 530 3982
rect 598 3978 602 3982
rect 622 3978 626 3982
rect 358 3958 362 3962
rect 462 3958 466 3962
rect 558 3968 562 3972
rect 582 3968 586 3972
rect 638 3998 642 4002
rect 662 4038 666 4042
rect 662 4018 666 4022
rect 646 3988 650 3992
rect 694 4058 698 4062
rect 686 4038 690 4042
rect 678 3968 682 3972
rect 726 4078 730 4082
rect 718 4048 722 4052
rect 694 4008 698 4012
rect 702 3978 706 3982
rect 726 3978 730 3982
rect 702 3968 706 3972
rect 374 3948 378 3952
rect 550 3948 554 3952
rect 582 3948 586 3952
rect 302 3908 306 3912
rect 326 3908 330 3912
rect 206 3848 210 3852
rect 214 3848 218 3852
rect 222 3818 226 3822
rect 206 3798 210 3802
rect 158 3778 162 3782
rect 134 3758 138 3762
rect 126 3678 130 3682
rect 150 3738 154 3742
rect 142 3698 146 3702
rect 110 3648 114 3652
rect 102 3578 106 3582
rect 110 3558 114 3562
rect 118 3548 122 3552
rect 134 3548 138 3552
rect 70 3538 74 3542
rect 86 3528 90 3532
rect 6 3468 10 3472
rect 54 3468 58 3472
rect 14 3338 18 3342
rect 22 3338 26 3342
rect 14 3288 18 3292
rect 62 3298 66 3302
rect 102 3518 106 3522
rect 134 3468 138 3472
rect 78 3368 82 3372
rect 118 3368 122 3372
rect 102 3348 106 3352
rect 110 3348 114 3352
rect 198 3728 202 3732
rect 190 3718 194 3722
rect 198 3708 202 3712
rect 214 3728 218 3732
rect 206 3698 210 3702
rect 262 3858 266 3862
rect 350 3878 354 3882
rect 374 3938 378 3942
rect 390 3938 394 3942
rect 406 3938 410 3942
rect 430 3938 434 3942
rect 406 3928 410 3932
rect 374 3888 378 3892
rect 366 3868 370 3872
rect 358 3858 362 3862
rect 262 3848 266 3852
rect 262 3838 266 3842
rect 238 3828 242 3832
rect 246 3788 250 3792
rect 254 3768 258 3772
rect 230 3748 234 3752
rect 190 3678 194 3682
rect 174 3668 178 3672
rect 206 3668 210 3672
rect 246 3668 250 3672
rect 310 3838 314 3842
rect 278 3828 282 3832
rect 278 3808 282 3812
rect 310 3798 314 3802
rect 350 3828 354 3832
rect 330 3803 334 3807
rect 337 3803 341 3807
rect 278 3778 282 3782
rect 278 3758 282 3762
rect 310 3758 314 3762
rect 262 3738 266 3742
rect 294 3738 298 3742
rect 318 3738 322 3742
rect 294 3728 298 3732
rect 374 3848 378 3852
rect 374 3838 378 3842
rect 366 3818 370 3822
rect 358 3748 362 3752
rect 382 3828 386 3832
rect 470 3938 474 3942
rect 454 3928 458 3932
rect 446 3918 450 3922
rect 430 3908 434 3912
rect 574 3938 578 3942
rect 486 3928 490 3932
rect 510 3928 514 3932
rect 478 3918 482 3922
rect 438 3878 442 3882
rect 486 3878 490 3882
rect 526 3918 530 3922
rect 566 3908 570 3912
rect 534 3878 538 3882
rect 502 3868 506 3872
rect 414 3848 418 3852
rect 390 3818 394 3822
rect 406 3768 410 3772
rect 446 3848 450 3852
rect 606 3938 610 3942
rect 646 3928 650 3932
rect 638 3918 642 3922
rect 654 3918 658 3922
rect 630 3888 634 3892
rect 574 3878 578 3882
rect 598 3878 602 3882
rect 686 3908 690 3912
rect 734 3968 738 3972
rect 734 3938 738 3942
rect 750 3938 754 3942
rect 750 3928 754 3932
rect 710 3878 714 3882
rect 494 3848 498 3852
rect 518 3848 522 3852
rect 478 3838 482 3842
rect 422 3788 426 3792
rect 446 3768 450 3772
rect 398 3748 402 3752
rect 414 3748 418 3752
rect 390 3738 394 3742
rect 326 3708 330 3712
rect 270 3668 274 3672
rect 166 3658 170 3662
rect 198 3658 202 3662
rect 254 3658 258 3662
rect 150 3648 154 3652
rect 262 3618 266 3622
rect 150 3558 154 3562
rect 158 3558 162 3562
rect 158 3538 162 3542
rect 174 3528 178 3532
rect 206 3528 210 3532
rect 222 3508 226 3512
rect 166 3468 170 3472
rect 206 3468 210 3472
rect 118 3338 122 3342
rect 142 3338 146 3342
rect 70 3268 74 3272
rect 102 3288 106 3292
rect 86 3258 90 3262
rect 110 3188 114 3192
rect 70 3148 74 3152
rect 86 3148 90 3152
rect 14 3138 18 3142
rect 22 3138 26 3142
rect 126 3118 130 3122
rect 78 3078 82 3082
rect 6 3068 10 3072
rect 166 3378 170 3382
rect 294 3608 298 3612
rect 330 3603 334 3607
rect 337 3603 341 3607
rect 398 3728 402 3732
rect 430 3728 434 3732
rect 406 3698 410 3702
rect 446 3698 450 3702
rect 462 3828 466 3832
rect 470 3818 474 3822
rect 550 3748 554 3752
rect 566 3748 570 3752
rect 462 3718 466 3722
rect 590 3728 594 3732
rect 774 3938 778 3942
rect 758 3918 762 3922
rect 766 3888 770 3892
rect 758 3868 762 3872
rect 702 3828 706 3832
rect 638 3768 642 3772
rect 662 3748 666 3752
rect 758 3748 762 3752
rect 646 3728 650 3732
rect 678 3728 682 3732
rect 486 3708 490 3712
rect 598 3708 602 3712
rect 686 3708 690 3712
rect 478 3688 482 3692
rect 566 3688 570 3692
rect 398 3678 402 3682
rect 454 3678 458 3682
rect 526 3678 530 3682
rect 590 3678 594 3682
rect 670 3678 674 3682
rect 430 3668 434 3672
rect 446 3668 450 3672
rect 390 3658 394 3662
rect 374 3598 378 3602
rect 366 3568 370 3572
rect 302 3558 306 3562
rect 262 3538 266 3542
rect 310 3538 314 3542
rect 326 3538 330 3542
rect 262 3518 266 3522
rect 246 3498 250 3502
rect 318 3528 322 3532
rect 718 3678 722 3682
rect 742 3678 746 3682
rect 758 3678 762 3682
rect 850 4103 854 4107
rect 857 4103 861 4107
rect 902 4138 906 4142
rect 870 4088 874 4092
rect 1182 4358 1186 4362
rect 1190 4348 1194 4352
rect 1478 4568 1482 4572
rect 1470 4558 1474 4562
rect 1502 4558 1506 4562
rect 1470 4538 1474 4542
rect 1454 4508 1458 4512
rect 1438 4498 1442 4502
rect 1470 4468 1474 4472
rect 1414 4458 1418 4462
rect 1446 4458 1450 4462
rect 1462 4458 1466 4462
rect 1350 4448 1354 4452
rect 1382 4448 1386 4452
rect 1430 4438 1434 4442
rect 1310 4388 1314 4392
rect 1354 4403 1358 4407
rect 1361 4403 1365 4407
rect 1390 4398 1394 4402
rect 1414 4398 1418 4402
rect 1326 4368 1330 4372
rect 1254 4358 1258 4362
rect 1326 4358 1330 4362
rect 1182 4338 1186 4342
rect 1222 4338 1226 4342
rect 1246 4328 1250 4332
rect 1198 4288 1202 4292
rect 1086 4278 1090 4282
rect 1094 4278 1098 4282
rect 1190 4278 1194 4282
rect 1078 4268 1082 4272
rect 1102 4268 1106 4272
rect 1118 4268 1122 4272
rect 1062 4258 1066 4262
rect 1142 4258 1146 4262
rect 1166 4258 1170 4262
rect 1086 4228 1090 4232
rect 1126 4228 1130 4232
rect 1150 4228 1154 4232
rect 1262 4338 1266 4342
rect 1406 4348 1410 4352
rect 1382 4338 1386 4342
rect 1326 4328 1330 4332
rect 1350 4278 1354 4282
rect 1358 4278 1362 4282
rect 1294 4268 1298 4272
rect 1326 4268 1330 4272
rect 1294 4258 1298 4262
rect 1382 4258 1386 4262
rect 1182 4218 1186 4222
rect 1246 4178 1250 4182
rect 1078 4168 1082 4172
rect 1174 4168 1178 4172
rect 1206 4158 1210 4162
rect 1222 4158 1226 4162
rect 1118 4148 1122 4152
rect 1166 4148 1170 4152
rect 1174 4148 1178 4152
rect 918 4138 922 4142
rect 950 4118 954 4122
rect 1006 4108 1010 4112
rect 982 4078 986 4082
rect 942 4068 946 4072
rect 998 4068 1002 4072
rect 814 4058 818 4062
rect 838 4058 842 4062
rect 878 4058 882 4062
rect 910 4058 914 4062
rect 950 4058 954 4062
rect 878 4048 882 4052
rect 934 4048 938 4052
rect 902 4038 906 4042
rect 934 4038 938 4042
rect 990 4038 994 4042
rect 838 4008 842 4012
rect 854 3978 858 3982
rect 998 3988 1002 3992
rect 958 3958 962 3962
rect 798 3948 802 3952
rect 902 3948 906 3952
rect 982 3948 986 3952
rect 838 3938 842 3942
rect 966 3938 970 3942
rect 806 3918 810 3922
rect 822 3918 826 3922
rect 790 3898 794 3902
rect 850 3903 854 3907
rect 857 3903 861 3907
rect 870 3878 874 3882
rect 958 3918 962 3922
rect 990 3918 994 3922
rect 918 3908 922 3912
rect 990 3898 994 3902
rect 918 3888 922 3892
rect 934 3888 938 3892
rect 910 3868 914 3872
rect 846 3858 850 3862
rect 958 3878 962 3882
rect 974 3878 978 3882
rect 934 3868 938 3872
rect 982 3868 986 3872
rect 942 3858 946 3862
rect 782 3748 786 3752
rect 846 3748 850 3752
rect 886 3748 890 3752
rect 734 3668 738 3672
rect 774 3668 778 3672
rect 790 3738 794 3742
rect 878 3738 882 3742
rect 910 3738 914 3742
rect 934 3738 938 3742
rect 918 3728 922 3732
rect 846 3718 850 3722
rect 894 3718 898 3722
rect 510 3658 514 3662
rect 582 3658 586 3662
rect 606 3658 610 3662
rect 638 3658 642 3662
rect 654 3658 658 3662
rect 758 3658 762 3662
rect 462 3608 466 3612
rect 590 3648 594 3652
rect 622 3648 626 3652
rect 590 3608 594 3612
rect 510 3588 514 3592
rect 494 3568 498 3572
rect 542 3568 546 3572
rect 566 3568 570 3572
rect 382 3558 386 3562
rect 422 3558 426 3562
rect 486 3558 490 3562
rect 438 3548 442 3552
rect 390 3538 394 3542
rect 518 3548 522 3552
rect 542 3548 546 3552
rect 510 3538 514 3542
rect 526 3538 530 3542
rect 342 3518 346 3522
rect 326 3488 330 3492
rect 286 3478 290 3482
rect 278 3468 282 3472
rect 302 3468 306 3472
rect 270 3458 274 3462
rect 294 3458 298 3462
rect 262 3448 266 3452
rect 310 3448 314 3452
rect 318 3428 322 3432
rect 478 3528 482 3532
rect 454 3498 458 3502
rect 446 3488 450 3492
rect 446 3468 450 3472
rect 390 3458 394 3462
rect 390 3428 394 3432
rect 342 3418 346 3422
rect 330 3403 334 3407
rect 337 3403 341 3407
rect 222 3358 226 3362
rect 174 3338 178 3342
rect 190 3318 194 3322
rect 190 3268 194 3272
rect 350 3378 354 3382
rect 262 3368 266 3372
rect 374 3368 378 3372
rect 318 3358 322 3362
rect 398 3418 402 3422
rect 278 3278 282 3282
rect 214 3268 218 3272
rect 198 3248 202 3252
rect 174 3168 178 3172
rect 214 3158 218 3162
rect 182 3148 186 3152
rect 182 3128 186 3132
rect 198 3128 202 3132
rect 166 3108 170 3112
rect 214 3118 218 3122
rect 166 3088 170 3092
rect 286 3258 290 3262
rect 438 3418 442 3422
rect 398 3318 402 3322
rect 382 3308 386 3312
rect 342 3298 346 3302
rect 462 3418 466 3422
rect 454 3408 458 3412
rect 446 3298 450 3302
rect 478 3408 482 3412
rect 478 3328 482 3332
rect 454 3278 458 3282
rect 438 3268 442 3272
rect 478 3258 482 3262
rect 630 3578 634 3582
rect 606 3548 610 3552
rect 630 3548 634 3552
rect 702 3648 706 3652
rect 726 3648 730 3652
rect 774 3638 778 3642
rect 662 3628 666 3632
rect 678 3588 682 3592
rect 662 3548 666 3552
rect 766 3568 770 3572
rect 782 3618 786 3622
rect 822 3659 826 3663
rect 806 3618 810 3622
rect 798 3588 802 3592
rect 790 3558 794 3562
rect 710 3548 714 3552
rect 798 3548 802 3552
rect 822 3588 826 3592
rect 638 3538 642 3542
rect 550 3528 554 3532
rect 566 3528 570 3532
rect 766 3528 770 3532
rect 662 3518 666 3522
rect 766 3518 770 3522
rect 542 3488 546 3492
rect 510 3478 514 3482
rect 502 3458 506 3462
rect 526 3458 530 3462
rect 494 3448 498 3452
rect 550 3448 554 3452
rect 518 3438 522 3442
rect 558 3428 562 3432
rect 502 3378 506 3382
rect 558 3368 562 3372
rect 598 3458 602 3462
rect 574 3448 578 3452
rect 574 3428 578 3432
rect 502 3358 506 3362
rect 566 3358 570 3362
rect 758 3478 762 3482
rect 662 3468 666 3472
rect 694 3468 698 3472
rect 638 3458 642 3462
rect 606 3418 610 3422
rect 622 3408 626 3412
rect 598 3398 602 3402
rect 614 3398 618 3402
rect 590 3358 594 3362
rect 518 3338 522 3342
rect 550 3338 554 3342
rect 558 3328 562 3332
rect 582 3328 586 3332
rect 598 3318 602 3322
rect 518 3308 522 3312
rect 534 3308 538 3312
rect 590 3298 594 3302
rect 558 3288 562 3292
rect 534 3268 538 3272
rect 494 3228 498 3232
rect 558 3228 562 3232
rect 334 3218 338 3222
rect 414 3218 418 3222
rect 486 3218 490 3222
rect 330 3203 334 3207
rect 337 3203 341 3207
rect 326 3168 330 3172
rect 302 3148 306 3152
rect 310 3148 314 3152
rect 254 3118 258 3122
rect 230 3108 234 3112
rect 222 3098 226 3102
rect 270 3078 274 3082
rect 214 3068 218 3072
rect 86 3058 90 3062
rect 102 3058 106 3062
rect 174 3058 178 3062
rect 62 2938 66 2942
rect 70 2928 74 2932
rect 14 2918 18 2922
rect 46 2858 50 2862
rect 158 3048 162 3052
rect 198 3048 202 3052
rect 166 2968 170 2972
rect 142 2958 146 2962
rect 126 2948 130 2952
rect 102 2918 106 2922
rect 102 2888 106 2892
rect 110 2878 114 2882
rect 222 2948 226 2952
rect 166 2928 170 2932
rect 150 2918 154 2922
rect 214 2918 218 2922
rect 206 2898 210 2902
rect 182 2878 186 2882
rect 110 2868 114 2872
rect 142 2868 146 2872
rect 158 2868 162 2872
rect 206 2868 210 2872
rect 150 2858 154 2862
rect 86 2848 90 2852
rect 102 2838 106 2842
rect 46 2748 50 2752
rect 62 2738 66 2742
rect 94 2678 98 2682
rect 110 2828 114 2832
rect 134 2828 138 2832
rect 190 2848 194 2852
rect 206 2848 210 2852
rect 198 2838 202 2842
rect 182 2818 186 2822
rect 118 2748 122 2752
rect 126 2748 130 2752
rect 110 2668 114 2672
rect 46 2658 50 2662
rect 38 2558 42 2562
rect 86 2578 90 2582
rect 158 2728 162 2732
rect 150 2688 154 2692
rect 134 2668 138 2672
rect 126 2658 130 2662
rect 166 2658 170 2662
rect 118 2618 122 2622
rect 134 2618 138 2622
rect 142 2618 146 2622
rect 134 2578 138 2582
rect 110 2568 114 2572
rect 126 2568 130 2572
rect 118 2548 122 2552
rect 102 2528 106 2532
rect 134 2508 138 2512
rect 94 2468 98 2472
rect 118 2458 122 2462
rect 38 2448 42 2452
rect 118 2448 122 2452
rect 158 2588 162 2592
rect 150 2568 154 2572
rect 182 2708 186 2712
rect 198 2678 202 2682
rect 246 2928 250 2932
rect 230 2898 234 2902
rect 566 3168 570 3172
rect 510 3158 514 3162
rect 582 3158 586 3162
rect 422 3148 426 3152
rect 342 3138 346 3142
rect 398 3128 402 3132
rect 390 3108 394 3112
rect 374 3098 378 3102
rect 374 3088 378 3092
rect 358 3068 362 3072
rect 278 2988 282 2992
rect 278 2868 282 2872
rect 246 2848 250 2852
rect 254 2838 258 2842
rect 278 2848 282 2852
rect 222 2738 226 2742
rect 230 2678 234 2682
rect 238 2678 242 2682
rect 182 2588 186 2592
rect 302 3018 306 3022
rect 326 3018 330 3022
rect 330 3003 334 3007
rect 337 3003 341 3007
rect 294 2978 298 2982
rect 310 2958 314 2962
rect 446 3138 450 3142
rect 502 3138 506 3142
rect 438 3128 442 3132
rect 414 3078 418 3082
rect 406 3068 410 3072
rect 478 3108 482 3112
rect 494 3088 498 3092
rect 566 3118 570 3122
rect 574 3108 578 3112
rect 510 3068 514 3072
rect 446 3058 450 3062
rect 558 3048 562 3052
rect 406 2988 410 2992
rect 454 2978 458 2982
rect 318 2948 322 2952
rect 350 2938 354 2942
rect 326 2918 330 2922
rect 302 2908 306 2912
rect 342 2898 346 2902
rect 294 2878 298 2882
rect 318 2878 322 2882
rect 310 2838 314 2842
rect 286 2768 290 2772
rect 270 2748 274 2752
rect 286 2748 290 2752
rect 374 2908 378 2912
rect 358 2868 362 2872
rect 366 2868 370 2872
rect 350 2858 354 2862
rect 366 2848 370 2852
rect 358 2838 362 2842
rect 330 2803 334 2807
rect 337 2803 341 2807
rect 342 2778 346 2782
rect 382 2828 386 2832
rect 398 2928 402 2932
rect 558 3028 562 3032
rect 574 3028 578 3032
rect 446 2898 450 2902
rect 542 2928 546 2932
rect 534 2908 538 2912
rect 534 2888 538 2892
rect 566 2888 570 2892
rect 494 2878 498 2882
rect 502 2878 506 2882
rect 574 2878 578 2882
rect 446 2868 450 2872
rect 502 2868 506 2872
rect 534 2868 538 2872
rect 398 2838 402 2842
rect 390 2808 394 2812
rect 382 2778 386 2782
rect 302 2718 306 2722
rect 318 2718 322 2722
rect 270 2698 274 2702
rect 270 2678 274 2682
rect 318 2708 322 2712
rect 214 2658 218 2662
rect 230 2658 234 2662
rect 246 2658 250 2662
rect 254 2658 258 2662
rect 286 2658 290 2662
rect 198 2558 202 2562
rect 214 2548 218 2552
rect 158 2538 162 2542
rect 190 2538 194 2542
rect 150 2498 154 2502
rect 166 2518 170 2522
rect 158 2478 162 2482
rect 150 2468 154 2472
rect 158 2448 162 2452
rect 110 2438 114 2442
rect 118 2348 122 2352
rect 38 2328 42 2332
rect 38 2278 42 2282
rect 150 2438 154 2442
rect 158 2358 162 2362
rect 126 2338 130 2342
rect 134 2338 138 2342
rect 142 2338 146 2342
rect 174 2498 178 2502
rect 270 2638 274 2642
rect 262 2568 266 2572
rect 278 2558 282 2562
rect 278 2548 282 2552
rect 262 2528 266 2532
rect 222 2518 226 2522
rect 262 2498 266 2502
rect 182 2478 186 2482
rect 302 2568 306 2572
rect 294 2558 298 2562
rect 294 2528 298 2532
rect 350 2698 354 2702
rect 350 2668 354 2672
rect 330 2603 334 2607
rect 337 2603 341 2607
rect 390 2748 394 2752
rect 710 3438 714 3442
rect 694 3408 698 3412
rect 718 3398 722 3402
rect 742 3378 746 3382
rect 750 3368 754 3372
rect 742 3358 746 3362
rect 638 3328 642 3332
rect 654 3328 658 3332
rect 670 3328 674 3332
rect 630 3308 634 3312
rect 622 3298 626 3302
rect 750 3338 754 3342
rect 774 3478 778 3482
rect 830 3558 834 3562
rect 830 3538 834 3542
rect 886 3708 890 3712
rect 850 3703 854 3707
rect 857 3703 861 3707
rect 846 3688 850 3692
rect 878 3678 882 3682
rect 926 3698 930 3702
rect 974 3738 978 3742
rect 958 3688 962 3692
rect 958 3678 962 3682
rect 1094 4088 1098 4092
rect 1046 4078 1050 4082
rect 1030 4038 1034 4042
rect 1078 3998 1082 4002
rect 1062 3978 1066 3982
rect 1046 3968 1050 3972
rect 1222 4138 1226 4142
rect 1230 4128 1234 4132
rect 1174 4118 1178 4122
rect 1238 4118 1242 4122
rect 1174 4098 1178 4102
rect 1110 4048 1114 4052
rect 1094 3958 1098 3962
rect 1006 3948 1010 3952
rect 1054 3948 1058 3952
rect 1030 3938 1034 3942
rect 1014 3928 1018 3932
rect 1006 3858 1010 3862
rect 1006 3848 1010 3852
rect 1054 3928 1058 3932
rect 1078 3918 1082 3922
rect 1022 3908 1026 3912
rect 1054 3878 1058 3882
rect 1190 4068 1194 4072
rect 1150 4058 1154 4062
rect 1166 4058 1170 4062
rect 1126 3948 1130 3952
rect 1110 3918 1114 3922
rect 1134 3918 1138 3922
rect 1046 3858 1050 3862
rect 1070 3858 1074 3862
rect 1054 3848 1058 3852
rect 1078 3848 1082 3852
rect 1086 3848 1090 3852
rect 1094 3848 1098 3852
rect 1038 3838 1042 3842
rect 1014 3828 1018 3832
rect 1022 3798 1026 3802
rect 1102 3798 1106 3802
rect 1094 3738 1098 3742
rect 966 3668 970 3672
rect 998 3668 1002 3672
rect 918 3658 922 3662
rect 974 3658 978 3662
rect 910 3648 914 3652
rect 942 3648 946 3652
rect 1030 3688 1034 3692
rect 1014 3678 1018 3682
rect 1158 4048 1162 4052
rect 1222 4038 1226 4042
rect 1150 3988 1154 3992
rect 1222 3968 1226 3972
rect 1230 3948 1234 3952
rect 1278 4238 1282 4242
rect 1366 4248 1370 4252
rect 1354 4203 1358 4207
rect 1361 4203 1365 4207
rect 1294 4178 1298 4182
rect 1286 4158 1290 4162
rect 1254 4138 1258 4142
rect 1246 4088 1250 4092
rect 1382 4148 1386 4152
rect 1294 4128 1298 4132
rect 1310 4128 1314 4132
rect 1470 4448 1474 4452
rect 1470 4358 1474 4362
rect 1446 4328 1450 4332
rect 1446 4318 1450 4322
rect 1454 4318 1458 4322
rect 1438 4288 1442 4292
rect 1398 4278 1402 4282
rect 1422 4278 1426 4282
rect 1430 4268 1434 4272
rect 1406 4258 1410 4262
rect 1422 4238 1426 4242
rect 1398 4178 1402 4182
rect 1334 4128 1338 4132
rect 1390 4128 1394 4132
rect 1310 4118 1314 4122
rect 1326 4118 1330 4122
rect 1286 4108 1290 4112
rect 1294 4088 1298 4092
rect 1302 4058 1306 4062
rect 1326 4058 1330 4062
rect 1358 4118 1362 4122
rect 1382 4118 1386 4122
rect 1390 4088 1394 4092
rect 1342 4078 1346 4082
rect 1358 4078 1362 4082
rect 1374 4068 1378 4072
rect 1414 4168 1418 4172
rect 1446 4258 1450 4262
rect 1494 4538 1498 4542
rect 1534 4678 1538 4682
rect 1566 4738 1570 4742
rect 1598 4738 1602 4742
rect 1566 4728 1570 4732
rect 1558 4698 1562 4702
rect 1606 4718 1610 4722
rect 1550 4658 1554 4662
rect 1574 4659 1578 4663
rect 1654 4798 1658 4802
rect 1646 4748 1650 4752
rect 1638 4718 1642 4722
rect 1646 4718 1650 4722
rect 1630 4708 1634 4712
rect 1646 4698 1650 4702
rect 1838 4788 1842 4792
rect 1870 4788 1874 4792
rect 1846 4778 1850 4782
rect 1854 4778 1858 4782
rect 1686 4748 1690 4752
rect 1726 4748 1730 4752
rect 1798 4748 1802 4752
rect 1830 4748 1834 4752
rect 1670 4738 1674 4742
rect 1678 4698 1682 4702
rect 1686 4688 1690 4692
rect 1598 4668 1602 4672
rect 1662 4668 1666 4672
rect 1590 4658 1594 4662
rect 1606 4608 1610 4612
rect 1574 4558 1578 4562
rect 1542 4538 1546 4542
rect 1510 4508 1514 4512
rect 1486 4488 1490 4492
rect 1590 4518 1594 4522
rect 1574 4488 1578 4492
rect 1686 4659 1690 4663
rect 1758 4718 1762 4722
rect 1726 4708 1730 4712
rect 1710 4648 1714 4652
rect 1694 4588 1698 4592
rect 1662 4558 1666 4562
rect 1614 4548 1618 4552
rect 1742 4698 1746 4702
rect 1798 4688 1802 4692
rect 1782 4678 1786 4682
rect 1758 4668 1762 4672
rect 1782 4668 1786 4672
rect 1774 4658 1778 4662
rect 1854 4758 1858 4762
rect 1878 4758 1882 4762
rect 1886 4748 1890 4752
rect 1894 4738 1898 4742
rect 1886 4728 1890 4732
rect 1874 4703 1878 4707
rect 1881 4703 1885 4707
rect 1886 4688 1890 4692
rect 1846 4658 1850 4662
rect 1814 4648 1818 4652
rect 1830 4648 1834 4652
rect 1774 4638 1778 4642
rect 1750 4628 1754 4632
rect 1742 4598 1746 4602
rect 1742 4578 1746 4582
rect 1638 4538 1642 4542
rect 1654 4538 1658 4542
rect 1686 4508 1690 4512
rect 1686 4498 1690 4502
rect 1614 4478 1618 4482
rect 1670 4478 1674 4482
rect 1710 4478 1714 4482
rect 1718 4478 1722 4482
rect 1622 4468 1626 4472
rect 1654 4468 1658 4472
rect 1518 4448 1522 4452
rect 1566 4448 1570 4452
rect 1582 4448 1586 4452
rect 1598 4378 1602 4382
rect 1630 4458 1634 4462
rect 1702 4438 1706 4442
rect 1702 4428 1706 4432
rect 1622 4368 1626 4372
rect 1598 4358 1602 4362
rect 1614 4358 1618 4362
rect 1486 4348 1490 4352
rect 1542 4348 1546 4352
rect 1566 4348 1570 4352
rect 1542 4328 1546 4332
rect 1558 4318 1562 4322
rect 1510 4278 1514 4282
rect 1486 4268 1490 4272
rect 1542 4268 1546 4272
rect 1550 4268 1554 4272
rect 1510 4258 1514 4262
rect 1502 4238 1506 4242
rect 1494 4218 1498 4222
rect 1478 4208 1482 4212
rect 1502 4208 1506 4212
rect 1470 4188 1474 4192
rect 1446 4178 1450 4182
rect 1486 4168 1490 4172
rect 1462 4158 1466 4162
rect 1438 4138 1442 4142
rect 1422 4118 1426 4122
rect 1398 4068 1402 4072
rect 1294 4038 1298 4042
rect 1302 4008 1306 4012
rect 1354 4003 1358 4007
rect 1361 4003 1365 4007
rect 1286 3998 1290 4002
rect 1278 3988 1282 3992
rect 1310 3988 1314 3992
rect 1286 3978 1290 3982
rect 1350 3968 1354 3972
rect 1374 3958 1378 3962
rect 1582 4328 1586 4332
rect 1614 4348 1618 4352
rect 1678 4348 1682 4352
rect 1606 4338 1610 4342
rect 1654 4338 1658 4342
rect 1598 4328 1602 4332
rect 1590 4308 1594 4312
rect 1574 4298 1578 4302
rect 1606 4298 1610 4302
rect 1622 4298 1626 4302
rect 1662 4298 1666 4302
rect 1526 4188 1530 4192
rect 1566 4188 1570 4192
rect 1502 4148 1506 4152
rect 1430 4078 1434 4082
rect 1462 4108 1466 4112
rect 1398 4048 1402 4052
rect 1446 4038 1450 4042
rect 1478 4078 1482 4082
rect 1502 4068 1506 4072
rect 1550 4178 1554 4182
rect 1606 4268 1610 4272
rect 1654 4278 1658 4282
rect 1678 4278 1682 4282
rect 1686 4278 1690 4282
rect 1574 4158 1578 4162
rect 1582 4138 1586 4142
rect 1534 4128 1538 4132
rect 1566 4128 1570 4132
rect 1534 4108 1538 4112
rect 1534 4068 1538 4072
rect 1550 4068 1554 4072
rect 1502 4038 1506 4042
rect 1518 4038 1522 4042
rect 1510 4018 1514 4022
rect 1462 3978 1466 3982
rect 1502 3978 1506 3982
rect 1502 3958 1506 3962
rect 1294 3948 1298 3952
rect 1334 3948 1338 3952
rect 1414 3948 1418 3952
rect 1486 3948 1490 3952
rect 1510 3948 1514 3952
rect 1398 3938 1402 3942
rect 1238 3928 1242 3932
rect 1278 3928 1282 3932
rect 1142 3908 1146 3912
rect 1150 3908 1154 3912
rect 1174 3908 1178 3912
rect 1214 3908 1218 3912
rect 1246 3908 1250 3912
rect 1174 3888 1178 3892
rect 1182 3878 1186 3882
rect 1198 3878 1202 3882
rect 1238 3878 1242 3882
rect 1334 3898 1338 3902
rect 1334 3878 1338 3882
rect 1382 3878 1386 3882
rect 1318 3868 1322 3872
rect 1182 3858 1186 3862
rect 1174 3798 1178 3802
rect 1142 3778 1146 3782
rect 1158 3768 1162 3772
rect 1158 3748 1162 3752
rect 1222 3858 1226 3862
rect 1262 3858 1266 3862
rect 1422 3878 1426 3882
rect 1366 3858 1370 3862
rect 1382 3858 1386 3862
rect 1398 3858 1402 3862
rect 1206 3848 1210 3852
rect 1254 3848 1258 3852
rect 1230 3818 1234 3822
rect 1214 3788 1218 3792
rect 1206 3768 1210 3772
rect 1238 3768 1242 3772
rect 1222 3748 1226 3752
rect 1166 3738 1170 3742
rect 1190 3738 1194 3742
rect 1254 3738 1258 3742
rect 1118 3728 1122 3732
rect 1182 3718 1186 3722
rect 1110 3708 1114 3712
rect 1190 3708 1194 3712
rect 1254 3698 1258 3702
rect 1398 3848 1402 3852
rect 1354 3803 1358 3807
rect 1361 3803 1365 3807
rect 1374 3778 1378 3782
rect 1438 3898 1442 3902
rect 1422 3828 1426 3832
rect 1470 3928 1474 3932
rect 1486 3928 1490 3932
rect 1510 3928 1514 3932
rect 1454 3898 1458 3902
rect 1534 4028 1538 4032
rect 1606 4128 1610 4132
rect 1622 4118 1626 4122
rect 1630 4108 1634 4112
rect 1606 4078 1610 4082
rect 1598 4058 1602 4062
rect 1574 4038 1578 4042
rect 1590 4008 1594 4012
rect 1542 3938 1546 3942
rect 1598 3938 1602 3942
rect 1550 3928 1554 3932
rect 1526 3918 1530 3922
rect 1486 3878 1490 3882
rect 1446 3828 1450 3832
rect 1550 3868 1554 3872
rect 1598 3878 1602 3882
rect 1630 3878 1634 3882
rect 1462 3858 1466 3862
rect 1550 3858 1554 3862
rect 1630 3858 1634 3862
rect 1454 3818 1458 3822
rect 1470 3808 1474 3812
rect 1446 3798 1450 3802
rect 1454 3788 1458 3792
rect 1414 3768 1418 3772
rect 1438 3768 1442 3772
rect 1486 3768 1490 3772
rect 1310 3738 1314 3742
rect 1390 3738 1394 3742
rect 1302 3728 1306 3732
rect 1286 3698 1290 3702
rect 1150 3688 1154 3692
rect 1110 3678 1114 3682
rect 1158 3678 1162 3682
rect 1246 3678 1250 3682
rect 1110 3668 1114 3672
rect 1006 3648 1010 3652
rect 950 3638 954 3642
rect 966 3638 970 3642
rect 926 3598 930 3602
rect 894 3548 898 3552
rect 854 3538 858 3542
rect 886 3538 890 3542
rect 902 3538 906 3542
rect 910 3528 914 3532
rect 870 3518 874 3522
rect 850 3503 854 3507
rect 857 3503 861 3507
rect 902 3508 906 3512
rect 878 3498 882 3502
rect 822 3488 826 3492
rect 870 3488 874 3492
rect 958 3588 962 3592
rect 998 3618 1002 3622
rect 1046 3618 1050 3622
rect 1054 3598 1058 3602
rect 1014 3568 1018 3572
rect 974 3558 978 3562
rect 998 3558 1002 3562
rect 1046 3548 1050 3552
rect 814 3478 818 3482
rect 886 3478 890 3482
rect 918 3478 922 3482
rect 910 3468 914 3472
rect 918 3458 922 3462
rect 806 3398 810 3402
rect 774 3368 778 3372
rect 862 3448 866 3452
rect 870 3438 874 3442
rect 926 3438 930 3442
rect 862 3418 866 3422
rect 798 3338 802 3342
rect 838 3338 842 3342
rect 854 3338 858 3342
rect 742 3328 746 3332
rect 742 3308 746 3312
rect 702 3298 706 3302
rect 678 3288 682 3292
rect 638 3278 642 3282
rect 694 3278 698 3282
rect 670 3268 674 3272
rect 638 3238 642 3242
rect 614 3208 618 3212
rect 654 3238 658 3242
rect 678 3238 682 3242
rect 862 3328 866 3332
rect 850 3303 854 3307
rect 857 3303 861 3307
rect 774 3288 778 3292
rect 758 3278 762 3282
rect 846 3278 850 3282
rect 734 3268 738 3272
rect 710 3238 714 3242
rect 734 3228 738 3232
rect 646 3198 650 3202
rect 686 3198 690 3202
rect 606 3178 610 3182
rect 638 3178 642 3182
rect 630 3168 634 3172
rect 710 3158 714 3162
rect 606 3148 610 3152
rect 622 3148 626 3152
rect 670 3148 674 3152
rect 694 3148 698 3152
rect 614 3138 618 3142
rect 590 3128 594 3132
rect 606 3128 610 3132
rect 598 3088 602 3092
rect 614 3068 618 3072
rect 838 3248 842 3252
rect 886 3358 890 3362
rect 886 3338 890 3342
rect 926 3338 930 3342
rect 902 3328 906 3332
rect 886 3278 890 3282
rect 910 3278 914 3282
rect 910 3248 914 3252
rect 918 3248 922 3252
rect 774 3238 778 3242
rect 870 3238 874 3242
rect 1126 3638 1130 3642
rect 1206 3668 1210 3672
rect 1246 3668 1250 3672
rect 1270 3668 1274 3672
rect 1182 3648 1186 3652
rect 1150 3638 1154 3642
rect 1142 3628 1146 3632
rect 1182 3628 1186 3632
rect 1166 3608 1170 3612
rect 1158 3588 1162 3592
rect 1094 3568 1098 3572
rect 1102 3568 1106 3572
rect 1094 3548 1098 3552
rect 1158 3548 1162 3552
rect 1246 3648 1250 3652
rect 1222 3638 1226 3642
rect 1358 3688 1362 3692
rect 1310 3678 1314 3682
rect 1302 3668 1306 3672
rect 1310 3668 1314 3672
rect 1310 3648 1314 3652
rect 1414 3738 1418 3742
rect 1606 3848 1610 3852
rect 1646 4188 1650 4192
rect 1758 4598 1762 4602
rect 1766 4558 1770 4562
rect 1774 4538 1778 4542
rect 1750 4508 1754 4512
rect 1742 4478 1746 4482
rect 1742 4458 1746 4462
rect 1726 4408 1730 4412
rect 1750 4368 1754 4372
rect 1782 4518 1786 4522
rect 1782 4488 1786 4492
rect 1806 4528 1810 4532
rect 1838 4508 1842 4512
rect 1862 4508 1866 4512
rect 1874 4503 1878 4507
rect 1881 4503 1885 4507
rect 1918 4538 1922 4542
rect 1894 4498 1898 4502
rect 1854 4478 1858 4482
rect 1918 4478 1922 4482
rect 1790 4458 1794 4462
rect 1806 4458 1810 4462
rect 1830 4458 1834 4462
rect 1846 4458 1850 4462
rect 1790 4448 1794 4452
rect 1798 4428 1802 4432
rect 1726 4358 1730 4362
rect 1766 4358 1770 4362
rect 1718 4348 1722 4352
rect 1766 4348 1770 4352
rect 1734 4328 1738 4332
rect 1694 4268 1698 4272
rect 1726 4308 1730 4312
rect 1742 4298 1746 4302
rect 1758 4318 1762 4322
rect 1782 4318 1786 4322
rect 1774 4298 1778 4302
rect 1750 4278 1754 4282
rect 1766 4278 1770 4282
rect 1742 4268 1746 4272
rect 1750 4258 1754 4262
rect 1694 4248 1698 4252
rect 1734 4248 1738 4252
rect 1758 4238 1762 4242
rect 1742 4208 1746 4212
rect 1694 4188 1698 4192
rect 1726 4188 1730 4192
rect 1678 4168 1682 4172
rect 1654 4158 1658 4162
rect 1662 4048 1666 4052
rect 1670 4038 1674 4042
rect 1734 4158 1738 4162
rect 1694 4128 1698 4132
rect 1734 4098 1738 4102
rect 1710 4078 1714 4082
rect 1726 4078 1730 4082
rect 1782 4248 1786 4252
rect 1774 4238 1778 4242
rect 1766 4198 1770 4202
rect 1782 4188 1786 4192
rect 1758 4138 1762 4142
rect 1758 4088 1762 4092
rect 1742 4078 1746 4082
rect 1774 4078 1778 4082
rect 1798 4178 1802 4182
rect 1814 4318 1818 4322
rect 1814 4308 1818 4312
rect 1846 4308 1850 4312
rect 1942 4738 1946 4742
rect 1966 4998 1970 5002
rect 2222 5058 2226 5062
rect 2318 5058 2322 5062
rect 2150 5048 2154 5052
rect 2350 5048 2354 5052
rect 2342 5038 2346 5042
rect 2086 5028 2090 5032
rect 2030 5018 2034 5022
rect 2134 4998 2138 5002
rect 2014 4948 2018 4952
rect 2030 4918 2034 4922
rect 1982 4878 1986 4882
rect 2078 4958 2082 4962
rect 2150 4958 2154 4962
rect 2262 5018 2266 5022
rect 2206 4988 2210 4992
rect 2198 4958 2202 4962
rect 2214 4958 2218 4962
rect 2070 4948 2074 4952
rect 2134 4948 2138 4952
rect 2182 4948 2186 4952
rect 2190 4948 2194 4952
rect 2238 4948 2242 4952
rect 2158 4928 2162 4932
rect 2054 4918 2058 4922
rect 2086 4918 2090 4922
rect 2094 4918 2098 4922
rect 2102 4908 2106 4912
rect 2070 4868 2074 4872
rect 1982 4858 1986 4862
rect 1990 4858 1994 4862
rect 2022 4858 2026 4862
rect 1966 4768 1970 4772
rect 2166 4868 2170 4872
rect 2142 4858 2146 4862
rect 2142 4848 2146 4852
rect 2158 4848 2162 4852
rect 2126 4788 2130 4792
rect 2118 4778 2122 4782
rect 1966 4758 1970 4762
rect 2046 4758 2050 4762
rect 2102 4758 2106 4762
rect 2110 4758 2114 4762
rect 2134 4758 2138 4762
rect 2190 4938 2194 4942
rect 2222 4938 2226 4942
rect 2206 4928 2210 4932
rect 2190 4858 2194 4862
rect 2174 4798 2178 4802
rect 2182 4798 2186 4802
rect 2158 4778 2162 4782
rect 2158 4748 2162 4752
rect 2022 4738 2026 4742
rect 2070 4738 2074 4742
rect 2150 4738 2154 4742
rect 1950 4698 1954 4702
rect 2006 4708 2010 4712
rect 2078 4698 2082 4702
rect 2086 4678 2090 4682
rect 1998 4668 2002 4672
rect 2014 4668 2018 4672
rect 2054 4668 2058 4672
rect 2006 4648 2010 4652
rect 1974 4608 1978 4612
rect 1950 4548 1954 4552
rect 1942 4538 1946 4542
rect 1958 4538 1962 4542
rect 1926 4378 1930 4382
rect 1894 4368 1898 4372
rect 1942 4368 1946 4372
rect 1934 4358 1938 4362
rect 1862 4338 1866 4342
rect 1878 4328 1882 4332
rect 1902 4318 1906 4322
rect 1874 4303 1878 4307
rect 1881 4303 1885 4307
rect 1918 4298 1922 4302
rect 1822 4278 1826 4282
rect 1814 4248 1818 4252
rect 1814 4228 1818 4232
rect 1814 4198 1818 4202
rect 1830 4258 1834 4262
rect 1958 4328 1962 4332
rect 1934 4258 1938 4262
rect 1838 4248 1842 4252
rect 1926 4248 1930 4252
rect 1862 4238 1866 4242
rect 1838 4188 1842 4192
rect 1830 4168 1834 4172
rect 1854 4148 1858 4152
rect 1822 4128 1826 4132
rect 1822 4118 1826 4122
rect 1830 4108 1834 4112
rect 1846 4088 1850 4092
rect 1838 4078 1842 4082
rect 1718 4058 1722 4062
rect 1750 4058 1754 4062
rect 1798 4058 1802 4062
rect 1830 4058 1834 4062
rect 1686 4028 1690 4032
rect 1702 3988 1706 3992
rect 1790 4048 1794 4052
rect 1830 4048 1834 4052
rect 1806 4038 1810 4042
rect 1750 3978 1754 3982
rect 1662 3968 1666 3972
rect 1694 3968 1698 3972
rect 1702 3968 1706 3972
rect 1654 3958 1658 3962
rect 1662 3948 1666 3952
rect 1686 3938 1690 3942
rect 1662 3928 1666 3932
rect 1670 3928 1674 3932
rect 1662 3878 1666 3882
rect 1646 3848 1650 3852
rect 1678 3828 1682 3832
rect 1638 3818 1642 3822
rect 1646 3808 1650 3812
rect 1542 3798 1546 3802
rect 1518 3768 1522 3772
rect 1470 3748 1474 3752
rect 1502 3748 1506 3752
rect 1486 3728 1490 3732
rect 1398 3698 1402 3702
rect 1486 3698 1490 3702
rect 1430 3678 1434 3682
rect 1478 3678 1482 3682
rect 1454 3668 1458 3672
rect 1406 3658 1410 3662
rect 1422 3658 1426 3662
rect 1374 3648 1378 3652
rect 1366 3628 1370 3632
rect 1278 3618 1282 3622
rect 1354 3603 1358 3607
rect 1361 3603 1365 3607
rect 1190 3598 1194 3602
rect 1214 3588 1218 3592
rect 1342 3588 1346 3592
rect 1342 3578 1346 3582
rect 1190 3558 1194 3562
rect 1214 3558 1218 3562
rect 1230 3558 1234 3562
rect 1022 3538 1026 3542
rect 1038 3538 1042 3542
rect 1174 3528 1178 3532
rect 1038 3518 1042 3522
rect 1006 3508 1010 3512
rect 966 3498 970 3502
rect 1070 3498 1074 3502
rect 942 3488 946 3492
rect 1062 3488 1066 3492
rect 1190 3488 1194 3492
rect 966 3478 970 3482
rect 1094 3478 1098 3482
rect 990 3468 994 3472
rect 1198 3468 1202 3472
rect 950 3458 954 3462
rect 942 3438 946 3442
rect 974 3398 978 3402
rect 982 3368 986 3372
rect 1006 3448 1010 3452
rect 1078 3438 1082 3442
rect 1094 3398 1098 3402
rect 1238 3548 1242 3552
rect 1270 3538 1274 3542
rect 1254 3478 1258 3482
rect 1350 3538 1354 3542
rect 1294 3528 1298 3532
rect 1390 3528 1394 3532
rect 1286 3518 1290 3522
rect 1278 3508 1282 3512
rect 1310 3508 1314 3512
rect 1334 3508 1338 3512
rect 1366 3508 1370 3512
rect 1278 3468 1282 3472
rect 1150 3458 1154 3462
rect 1238 3458 1242 3462
rect 1286 3458 1290 3462
rect 1198 3448 1202 3452
rect 1238 3448 1242 3452
rect 1286 3448 1290 3452
rect 1254 3418 1258 3422
rect 1414 3618 1418 3622
rect 1422 3558 1426 3562
rect 1478 3658 1482 3662
rect 1438 3648 1442 3652
rect 1502 3688 1506 3692
rect 1502 3668 1506 3672
rect 1574 3788 1578 3792
rect 1606 3748 1610 3752
rect 1614 3748 1618 3752
rect 1670 3748 1674 3752
rect 1646 3738 1650 3742
rect 1550 3728 1554 3732
rect 1638 3728 1642 3732
rect 1646 3728 1650 3732
rect 1550 3718 1554 3722
rect 1598 3688 1602 3692
rect 1566 3678 1570 3682
rect 1582 3668 1586 3672
rect 1510 3658 1514 3662
rect 1574 3658 1578 3662
rect 1614 3658 1618 3662
rect 1494 3638 1498 3642
rect 1550 3638 1554 3642
rect 1582 3638 1586 3642
rect 1606 3638 1610 3642
rect 1622 3638 1626 3642
rect 1462 3608 1466 3612
rect 1486 3598 1490 3602
rect 1470 3588 1474 3592
rect 1446 3568 1450 3572
rect 1414 3488 1418 3492
rect 1406 3468 1410 3472
rect 1354 3403 1358 3407
rect 1361 3403 1365 3407
rect 1478 3558 1482 3562
rect 1662 3688 1666 3692
rect 1638 3638 1642 3642
rect 1830 4008 1834 4012
rect 1806 3998 1810 4002
rect 1774 3968 1778 3972
rect 1758 3948 1762 3952
rect 1790 3948 1794 3952
rect 1798 3948 1802 3952
rect 1750 3938 1754 3942
rect 1806 3938 1810 3942
rect 1790 3928 1794 3932
rect 1718 3918 1722 3922
rect 1734 3908 1738 3912
rect 1718 3898 1722 3902
rect 1750 3898 1754 3902
rect 1710 3878 1714 3882
rect 1814 3928 1818 3932
rect 1806 3908 1810 3912
rect 1822 3898 1826 3902
rect 2046 4648 2050 4652
rect 2094 4638 2098 4642
rect 2038 4628 2042 4632
rect 2070 4628 2074 4632
rect 2094 4588 2098 4592
rect 2038 4558 2042 4562
rect 2118 4708 2122 4712
rect 2110 4668 2114 4672
rect 2110 4558 2114 4562
rect 2134 4558 2138 4562
rect 2118 4548 2122 4552
rect 2110 4528 2114 4532
rect 2022 4498 2026 4502
rect 2102 4498 2106 4502
rect 2014 4488 2018 4492
rect 2070 4488 2074 4492
rect 2078 4468 2082 4472
rect 2102 4468 2106 4472
rect 1998 4448 2002 4452
rect 2022 4448 2026 4452
rect 2030 4448 2034 4452
rect 1990 4358 1994 4362
rect 1990 4318 1994 4322
rect 2302 5008 2306 5012
rect 2254 4928 2258 4932
rect 2262 4928 2266 4932
rect 2486 5068 2490 5072
rect 2510 5068 2514 5072
rect 2558 5068 2562 5072
rect 2662 5068 2666 5072
rect 2742 5068 2746 5072
rect 3022 5068 3026 5072
rect 3078 5068 3082 5072
rect 3118 5068 3122 5072
rect 3150 5068 3154 5072
rect 3182 5068 3186 5072
rect 3262 5068 3266 5072
rect 3366 5068 3370 5072
rect 3470 5068 3474 5072
rect 3566 5068 3570 5072
rect 3766 5068 3770 5072
rect 3926 5068 3930 5072
rect 3958 5068 3962 5072
rect 4030 5068 4034 5072
rect 4390 5068 4394 5072
rect 4854 5068 4858 5072
rect 5046 5068 5050 5072
rect 5238 5068 5242 5072
rect 2454 5048 2458 5052
rect 2454 5038 2458 5042
rect 2406 5018 2410 5022
rect 2430 5018 2434 5022
rect 2446 5018 2450 5022
rect 2386 5003 2390 5007
rect 2393 5003 2397 5007
rect 2390 4988 2394 4992
rect 2406 4978 2410 4982
rect 2318 4948 2322 4952
rect 2334 4948 2338 4952
rect 2350 4948 2354 4952
rect 2326 4938 2330 4942
rect 2326 4878 2330 4882
rect 2222 4848 2226 4852
rect 2326 4848 2330 4852
rect 2206 4808 2210 4812
rect 2222 4798 2226 4802
rect 2214 4778 2218 4782
rect 2190 4768 2194 4772
rect 2182 4738 2186 4742
rect 2254 4768 2258 4772
rect 2206 4748 2210 4752
rect 2270 4748 2274 4752
rect 2278 4738 2282 4742
rect 2414 4958 2418 4962
rect 2502 5058 2506 5062
rect 2542 5058 2546 5062
rect 2638 5058 2642 5062
rect 2486 5038 2490 5042
rect 2478 4998 2482 5002
rect 2438 4948 2442 4952
rect 2470 4948 2474 4952
rect 2494 4948 2498 4952
rect 2406 4918 2410 4922
rect 2422 4918 2426 4922
rect 2414 4888 2418 4892
rect 2334 4808 2338 4812
rect 2294 4758 2298 4762
rect 2414 4808 2418 4812
rect 2386 4803 2390 4807
rect 2393 4803 2397 4807
rect 2454 4878 2458 4882
rect 2430 4868 2434 4872
rect 2486 4928 2490 4932
rect 2614 5048 2618 5052
rect 2510 5038 2514 5042
rect 2518 5028 2522 5032
rect 2558 4978 2562 4982
rect 2582 4968 2586 4972
rect 2566 4958 2570 4962
rect 2790 5058 2794 5062
rect 2822 5058 2826 5062
rect 2894 5058 2898 5062
rect 2774 5048 2778 5052
rect 2742 5038 2746 5042
rect 2766 5038 2770 5042
rect 2638 5018 2642 5022
rect 2726 5018 2730 5022
rect 2622 4958 2626 4962
rect 2790 4978 2794 4982
rect 2662 4968 2666 4972
rect 2694 4958 2698 4962
rect 2526 4948 2530 4952
rect 2550 4948 2554 4952
rect 2566 4948 2570 4952
rect 2646 4948 2650 4952
rect 2862 4968 2866 4972
rect 2894 4968 2898 4972
rect 2870 4948 2874 4952
rect 2510 4938 2514 4942
rect 2542 4938 2546 4942
rect 2638 4938 2642 4942
rect 2502 4868 2506 4872
rect 2438 4858 2442 4862
rect 2478 4858 2482 4862
rect 2438 4838 2442 4842
rect 2598 4918 2602 4922
rect 2574 4888 2578 4892
rect 2558 4878 2562 4882
rect 2574 4878 2578 4882
rect 2630 4898 2634 4902
rect 2590 4868 2594 4872
rect 2582 4858 2586 4862
rect 2590 4858 2594 4862
rect 2606 4858 2610 4862
rect 2670 4918 2674 4922
rect 2646 4878 2650 4882
rect 2518 4848 2522 4852
rect 2542 4848 2546 4852
rect 2510 4808 2514 4812
rect 2462 4788 2466 4792
rect 2430 4778 2434 4782
rect 2422 4758 2426 4762
rect 2454 4748 2458 4752
rect 2166 4638 2170 4642
rect 2174 4618 2178 4622
rect 2358 4738 2362 4742
rect 2334 4718 2338 4722
rect 2214 4668 2218 4672
rect 2206 4658 2210 4662
rect 2286 4698 2290 4702
rect 2310 4688 2314 4692
rect 2390 4708 2394 4712
rect 2270 4678 2274 4682
rect 2294 4678 2298 4682
rect 2286 4648 2290 4652
rect 2326 4648 2330 4652
rect 2278 4638 2282 4642
rect 2230 4578 2234 4582
rect 2190 4558 2194 4562
rect 2190 4538 2194 4542
rect 2158 4488 2162 4492
rect 2070 4458 2074 4462
rect 2094 4458 2098 4462
rect 2126 4458 2130 4462
rect 2110 4398 2114 4402
rect 2070 4368 2074 4372
rect 2054 4328 2058 4332
rect 2046 4318 2050 4322
rect 1974 4308 1978 4312
rect 1990 4308 1994 4312
rect 1998 4308 2002 4312
rect 2022 4298 2026 4302
rect 2038 4298 2042 4302
rect 2062 4298 2066 4302
rect 2014 4268 2018 4272
rect 1966 4248 1970 4252
rect 1958 4238 1962 4242
rect 1998 4238 2002 4242
rect 1926 4218 1930 4222
rect 1878 4188 1882 4192
rect 1934 4168 1938 4172
rect 1886 4158 1890 4162
rect 1902 4158 1906 4162
rect 1870 4138 1874 4142
rect 1874 4103 1878 4107
rect 1881 4103 1885 4107
rect 1926 4148 1930 4152
rect 1902 4138 1906 4142
rect 1902 4118 1906 4122
rect 1974 4228 1978 4232
rect 1990 4208 1994 4212
rect 2086 4358 2090 4362
rect 2102 4348 2106 4352
rect 2158 4398 2162 4402
rect 2150 4358 2154 4362
rect 2214 4548 2218 4552
rect 2222 4538 2226 4542
rect 2206 4518 2210 4522
rect 2190 4468 2194 4472
rect 2262 4528 2266 4532
rect 2238 4478 2242 4482
rect 2222 4458 2226 4462
rect 2198 4418 2202 4422
rect 2182 4368 2186 4372
rect 2366 4638 2370 4642
rect 2386 4603 2390 4607
rect 2393 4603 2397 4607
rect 2326 4568 2330 4572
rect 2358 4558 2362 4562
rect 2398 4558 2402 4562
rect 2286 4538 2290 4542
rect 2302 4448 2306 4452
rect 2278 4418 2282 4422
rect 2262 4398 2266 4402
rect 2222 4358 2226 4362
rect 2190 4348 2194 4352
rect 2238 4348 2242 4352
rect 2150 4328 2154 4332
rect 2166 4328 2170 4332
rect 2150 4308 2154 4312
rect 2086 4278 2090 4282
rect 2142 4278 2146 4282
rect 2054 4228 2058 4232
rect 2054 4218 2058 4222
rect 1998 4198 2002 4202
rect 2046 4198 2050 4202
rect 2030 4158 2034 4162
rect 2142 4268 2146 4272
rect 2126 4258 2130 4262
rect 2102 4248 2106 4252
rect 2086 4188 2090 4192
rect 2094 4188 2098 4192
rect 2142 4188 2146 4192
rect 2078 4168 2082 4172
rect 2070 4158 2074 4162
rect 1966 4138 1970 4142
rect 2046 4138 2050 4142
rect 1918 4108 1922 4112
rect 1974 4108 1978 4112
rect 1934 4078 1938 4082
rect 1950 4078 1954 4082
rect 1950 4058 1954 4062
rect 1958 4058 1962 4062
rect 1862 4048 1866 4052
rect 1918 4048 1922 4052
rect 1918 4028 1922 4032
rect 1854 4008 1858 4012
rect 1846 3998 1850 4002
rect 1870 3948 1874 3952
rect 1902 3948 1906 3952
rect 1830 3888 1834 3892
rect 1782 3878 1786 3882
rect 1814 3878 1818 3882
rect 1758 3868 1762 3872
rect 1830 3868 1834 3872
rect 1694 3858 1698 3862
rect 1726 3858 1730 3862
rect 1806 3858 1810 3862
rect 1798 3848 1802 3852
rect 1830 3848 1834 3852
rect 1694 3798 1698 3802
rect 1702 3778 1706 3782
rect 1766 3808 1770 3812
rect 1790 3788 1794 3792
rect 1734 3748 1738 3752
rect 1750 3748 1754 3752
rect 1742 3738 1746 3742
rect 1710 3708 1714 3712
rect 1686 3698 1690 3702
rect 1734 3728 1738 3732
rect 1718 3678 1722 3682
rect 1750 3678 1754 3682
rect 1630 3628 1634 3632
rect 1654 3628 1658 3632
rect 1662 3628 1666 3632
rect 1630 3598 1634 3602
rect 1662 3588 1666 3592
rect 1502 3568 1506 3572
rect 1622 3568 1626 3572
rect 1502 3548 1506 3552
rect 1526 3548 1530 3552
rect 1534 3548 1538 3552
rect 1574 3548 1578 3552
rect 1686 3598 1690 3602
rect 1670 3558 1674 3562
rect 1590 3548 1594 3552
rect 1614 3548 1618 3552
rect 1638 3548 1642 3552
rect 1654 3548 1658 3552
rect 1486 3538 1490 3542
rect 1454 3528 1458 3532
rect 1454 3518 1458 3522
rect 1430 3508 1434 3512
rect 1470 3488 1474 3492
rect 1470 3468 1474 3472
rect 1422 3398 1426 3402
rect 1118 3388 1122 3392
rect 1206 3388 1210 3392
rect 1310 3388 1314 3392
rect 1382 3388 1386 3392
rect 1134 3378 1138 3382
rect 966 3308 970 3312
rect 838 3228 842 3232
rect 934 3228 938 3232
rect 750 3218 754 3222
rect 774 3178 778 3182
rect 758 3158 762 3162
rect 790 3158 794 3162
rect 878 3218 882 3222
rect 918 3218 922 3222
rect 870 3208 874 3212
rect 870 3178 874 3182
rect 870 3158 874 3162
rect 902 3198 906 3202
rect 886 3178 890 3182
rect 934 3208 938 3212
rect 950 3198 954 3202
rect 934 3158 938 3162
rect 790 3148 794 3152
rect 822 3148 826 3152
rect 830 3148 834 3152
rect 894 3148 898 3152
rect 910 3148 914 3152
rect 678 3138 682 3142
rect 718 3138 722 3142
rect 646 3118 650 3122
rect 726 3118 730 3122
rect 630 3088 634 3092
rect 678 3098 682 3102
rect 662 3078 666 3082
rect 678 3078 682 3082
rect 662 3068 666 3072
rect 598 3058 602 3062
rect 622 3058 626 3062
rect 662 3058 666 3062
rect 646 3048 650 3052
rect 614 3018 618 3022
rect 606 2968 610 2972
rect 606 2958 610 2962
rect 694 3048 698 3052
rect 766 3108 770 3112
rect 750 3088 754 3092
rect 814 3128 818 3132
rect 782 3118 786 3122
rect 798 3118 802 3122
rect 774 3088 778 3092
rect 774 3058 778 3062
rect 750 3018 754 3022
rect 662 2998 666 3002
rect 766 3008 770 3012
rect 790 3058 794 3062
rect 806 3058 810 3062
rect 814 3038 818 3042
rect 742 2988 746 2992
rect 750 2988 754 2992
rect 774 2988 778 2992
rect 734 2978 738 2982
rect 654 2968 658 2972
rect 622 2938 626 2942
rect 638 2938 642 2942
rect 630 2928 634 2932
rect 590 2888 594 2892
rect 710 2958 714 2962
rect 678 2938 682 2942
rect 686 2928 690 2932
rect 718 2938 722 2942
rect 686 2918 690 2922
rect 694 2918 698 2922
rect 646 2898 650 2902
rect 670 2898 674 2902
rect 662 2888 666 2892
rect 622 2878 626 2882
rect 638 2878 642 2882
rect 678 2878 682 2882
rect 582 2868 586 2872
rect 662 2868 666 2872
rect 526 2858 530 2862
rect 494 2788 498 2792
rect 502 2778 506 2782
rect 510 2758 514 2762
rect 534 2848 538 2852
rect 542 2838 546 2842
rect 630 2848 634 2852
rect 598 2838 602 2842
rect 614 2838 618 2842
rect 566 2828 570 2832
rect 558 2798 562 2802
rect 574 2788 578 2792
rect 638 2808 642 2812
rect 630 2798 634 2802
rect 582 2778 586 2782
rect 614 2778 618 2782
rect 550 2758 554 2762
rect 566 2758 570 2762
rect 526 2748 530 2752
rect 406 2738 410 2742
rect 382 2718 386 2722
rect 366 2708 370 2712
rect 518 2738 522 2742
rect 454 2728 458 2732
rect 430 2698 434 2702
rect 654 2758 658 2762
rect 686 2818 690 2822
rect 718 2898 722 2902
rect 702 2888 706 2892
rect 758 2968 762 2972
rect 806 2948 810 2952
rect 750 2918 754 2922
rect 766 2918 770 2922
rect 782 2908 786 2912
rect 814 2908 818 2912
rect 734 2868 738 2872
rect 806 2888 810 2892
rect 742 2848 746 2852
rect 710 2838 714 2842
rect 694 2808 698 2812
rect 702 2808 706 2812
rect 694 2788 698 2792
rect 718 2788 722 2792
rect 726 2758 730 2762
rect 766 2808 770 2812
rect 598 2748 602 2752
rect 622 2748 626 2752
rect 638 2748 642 2752
rect 710 2748 714 2752
rect 742 2748 746 2752
rect 542 2728 546 2732
rect 550 2728 554 2732
rect 630 2728 634 2732
rect 718 2728 722 2732
rect 742 2728 746 2732
rect 598 2708 602 2712
rect 590 2698 594 2702
rect 606 2698 610 2702
rect 614 2698 618 2702
rect 478 2688 482 2692
rect 558 2688 562 2692
rect 582 2688 586 2692
rect 638 2688 642 2692
rect 422 2678 426 2682
rect 430 2678 434 2682
rect 590 2668 594 2672
rect 646 2668 650 2672
rect 438 2658 442 2662
rect 574 2658 578 2662
rect 662 2658 666 2662
rect 430 2648 434 2652
rect 478 2648 482 2652
rect 558 2648 562 2652
rect 382 2638 386 2642
rect 406 2638 410 2642
rect 358 2578 362 2582
rect 326 2568 330 2572
rect 358 2568 362 2572
rect 366 2558 370 2562
rect 390 2618 394 2622
rect 374 2548 378 2552
rect 606 2648 610 2652
rect 446 2638 450 2642
rect 486 2638 490 2642
rect 502 2638 506 2642
rect 550 2638 554 2642
rect 566 2638 570 2642
rect 422 2608 426 2612
rect 406 2548 410 2552
rect 350 2538 354 2542
rect 318 2528 322 2532
rect 318 2518 322 2522
rect 310 2488 314 2492
rect 222 2468 226 2472
rect 310 2468 314 2472
rect 414 2528 418 2532
rect 398 2508 402 2512
rect 350 2488 354 2492
rect 334 2478 338 2482
rect 182 2458 186 2462
rect 286 2458 290 2462
rect 318 2458 322 2462
rect 246 2428 250 2432
rect 230 2418 234 2422
rect 222 2358 226 2362
rect 150 2288 154 2292
rect 126 2278 130 2282
rect 118 2268 122 2272
rect 150 2268 154 2272
rect 174 2328 178 2332
rect 182 2318 186 2322
rect 166 2288 170 2292
rect 174 2268 178 2272
rect 134 2258 138 2262
rect 206 2348 210 2352
rect 206 2288 210 2292
rect 214 2268 218 2272
rect 190 2258 194 2262
rect 182 2178 186 2182
rect 174 2168 178 2172
rect 150 2158 154 2162
rect 118 2148 122 2152
rect 190 2138 194 2142
rect 174 2128 178 2132
rect 166 2078 170 2082
rect 70 2058 74 2062
rect 86 2058 90 2062
rect 118 2058 122 2062
rect 62 1988 66 1992
rect 14 1938 18 1942
rect 6 1898 10 1902
rect 238 2328 242 2332
rect 222 2258 226 2262
rect 230 2258 234 2262
rect 206 2178 210 2182
rect 222 2178 226 2182
rect 206 2168 210 2172
rect 486 2578 490 2582
rect 446 2568 450 2572
rect 438 2548 442 2552
rect 462 2558 466 2562
rect 614 2608 618 2612
rect 566 2598 570 2602
rect 486 2538 490 2542
rect 470 2528 474 2532
rect 462 2518 466 2522
rect 422 2498 426 2502
rect 438 2498 442 2502
rect 414 2448 418 2452
rect 390 2438 394 2442
rect 278 2408 282 2412
rect 318 2408 322 2412
rect 330 2403 334 2407
rect 337 2403 341 2407
rect 374 2378 378 2382
rect 318 2358 322 2362
rect 302 2338 306 2342
rect 350 2328 354 2332
rect 278 2318 282 2322
rect 270 2308 274 2312
rect 294 2308 298 2312
rect 286 2298 290 2302
rect 262 2278 266 2282
rect 286 2278 290 2282
rect 302 2278 306 2282
rect 294 2268 298 2272
rect 414 2358 418 2362
rect 446 2448 450 2452
rect 454 2428 458 2432
rect 470 2498 474 2502
rect 486 2518 490 2522
rect 478 2488 482 2492
rect 462 2418 466 2422
rect 446 2408 450 2412
rect 478 2438 482 2442
rect 470 2378 474 2382
rect 462 2358 466 2362
rect 438 2348 442 2352
rect 454 2338 458 2342
rect 422 2308 426 2312
rect 390 2288 394 2292
rect 406 2288 410 2292
rect 446 2288 450 2292
rect 398 2268 402 2272
rect 430 2268 434 2272
rect 446 2268 450 2272
rect 246 2258 250 2262
rect 294 2258 298 2262
rect 302 2258 306 2262
rect 358 2258 362 2262
rect 422 2258 426 2262
rect 566 2538 570 2542
rect 550 2528 554 2532
rect 542 2508 546 2512
rect 494 2468 498 2472
rect 558 2478 562 2482
rect 606 2488 610 2492
rect 590 2478 594 2482
rect 630 2528 634 2532
rect 574 2468 578 2472
rect 518 2458 522 2462
rect 542 2458 546 2462
rect 606 2458 610 2462
rect 510 2448 514 2452
rect 526 2448 530 2452
rect 502 2368 506 2372
rect 542 2368 546 2372
rect 590 2388 594 2392
rect 646 2468 650 2472
rect 822 2798 826 2802
rect 814 2748 818 2752
rect 790 2728 794 2732
rect 798 2718 802 2722
rect 790 2708 794 2712
rect 774 2698 778 2702
rect 718 2668 722 2672
rect 726 2668 730 2672
rect 734 2668 738 2672
rect 710 2638 714 2642
rect 758 2668 762 2672
rect 766 2658 770 2662
rect 766 2648 770 2652
rect 742 2638 746 2642
rect 718 2628 722 2632
rect 670 2618 674 2622
rect 854 3138 858 3142
rect 950 3138 954 3142
rect 894 3128 898 3132
rect 838 3108 842 3112
rect 850 3103 854 3107
rect 857 3103 861 3107
rect 990 3358 994 3362
rect 1038 3368 1042 3372
rect 1014 3358 1018 3362
rect 990 3338 994 3342
rect 998 3258 1002 3262
rect 1022 3338 1026 3342
rect 1118 3338 1122 3342
rect 1062 3328 1066 3332
rect 1078 3328 1082 3332
rect 1126 3328 1130 3332
rect 1102 3268 1106 3272
rect 1086 3258 1090 3262
rect 1174 3368 1178 3372
rect 1142 3358 1146 3362
rect 1198 3358 1202 3362
rect 1158 3338 1162 3342
rect 1142 3328 1146 3332
rect 1150 3308 1154 3312
rect 1142 3278 1146 3282
rect 1254 3378 1258 3382
rect 1262 3378 1266 3382
rect 1318 3368 1322 3372
rect 1278 3358 1282 3362
rect 1294 3358 1298 3362
rect 1326 3358 1330 3362
rect 1166 3268 1170 3272
rect 1174 3268 1178 3272
rect 1078 3248 1082 3252
rect 1102 3248 1106 3252
rect 1126 3248 1130 3252
rect 1158 3248 1162 3252
rect 1206 3248 1210 3252
rect 1022 3218 1026 3222
rect 1006 3208 1010 3212
rect 1014 3178 1018 3182
rect 1030 3148 1034 3152
rect 1054 3138 1058 3142
rect 966 3128 970 3132
rect 1014 3128 1018 3132
rect 1022 3098 1026 3102
rect 1134 3198 1138 3202
rect 1182 3238 1186 3242
rect 1206 3208 1210 3212
rect 1094 3168 1098 3172
rect 1126 3168 1130 3172
rect 1086 3148 1090 3152
rect 1158 3158 1162 3162
rect 1222 3178 1226 3182
rect 1342 3340 1346 3344
rect 1462 3458 1466 3462
rect 1446 3388 1450 3392
rect 1422 3378 1426 3382
rect 1462 3358 1466 3362
rect 1318 3318 1322 3322
rect 1270 3308 1274 3312
rect 1302 3268 1306 3272
rect 1342 3268 1346 3272
rect 1270 3238 1274 3242
rect 1270 3228 1274 3232
rect 1326 3248 1330 3252
rect 1294 3238 1298 3242
rect 1326 3228 1330 3232
rect 1310 3218 1314 3222
rect 1494 3528 1498 3532
rect 1534 3518 1538 3522
rect 1542 3508 1546 3512
rect 1510 3488 1514 3492
rect 1526 3488 1530 3492
rect 1518 3468 1522 3472
rect 1494 3458 1498 3462
rect 1510 3458 1514 3462
rect 1566 3528 1570 3532
rect 1574 3528 1578 3532
rect 1590 3528 1594 3532
rect 1558 3518 1562 3522
rect 1574 3518 1578 3522
rect 1558 3508 1562 3512
rect 1566 3468 1570 3472
rect 1486 3438 1490 3442
rect 1502 3408 1506 3412
rect 1494 3378 1498 3382
rect 1502 3358 1506 3362
rect 1406 3328 1410 3332
rect 1470 3328 1474 3332
rect 1478 3328 1482 3332
rect 1518 3448 1522 3452
rect 1550 3448 1554 3452
rect 1534 3438 1538 3442
rect 1542 3428 1546 3432
rect 1534 3418 1538 3422
rect 1526 3378 1530 3382
rect 1518 3368 1522 3372
rect 1550 3368 1554 3372
rect 1542 3358 1546 3362
rect 1526 3328 1530 3332
rect 1510 3308 1514 3312
rect 1390 3288 1394 3292
rect 1494 3288 1498 3292
rect 1526 3288 1530 3292
rect 1478 3278 1482 3282
rect 1510 3278 1514 3282
rect 1630 3528 1634 3532
rect 1622 3508 1626 3512
rect 1598 3488 1602 3492
rect 1590 3478 1594 3482
rect 1654 3478 1658 3482
rect 1702 3548 1706 3552
rect 1686 3528 1690 3532
rect 1710 3498 1714 3502
rect 1782 3668 1786 3672
rect 1726 3648 1730 3652
rect 1790 3628 1794 3632
rect 1790 3588 1794 3592
rect 1766 3578 1770 3582
rect 1790 3558 1794 3562
rect 1774 3548 1778 3552
rect 1750 3538 1754 3542
rect 1766 3538 1770 3542
rect 1790 3538 1794 3542
rect 1758 3528 1762 3532
rect 1750 3508 1754 3512
rect 1718 3488 1722 3492
rect 1750 3488 1754 3492
rect 1774 3478 1778 3482
rect 1942 3988 1946 3992
rect 1966 3988 1970 3992
rect 1926 3978 1930 3982
rect 1958 3978 1962 3982
rect 1942 3948 1946 3952
rect 1934 3938 1938 3942
rect 1918 3918 1922 3922
rect 1874 3903 1878 3907
rect 1881 3903 1885 3907
rect 1886 3888 1890 3892
rect 1894 3868 1898 3872
rect 1878 3838 1882 3842
rect 1830 3828 1834 3832
rect 1854 3828 1858 3832
rect 1814 3768 1818 3772
rect 1854 3778 1858 3782
rect 1902 3858 1906 3862
rect 1910 3798 1914 3802
rect 1910 3778 1914 3782
rect 1886 3758 1890 3762
rect 1878 3748 1882 3752
rect 1846 3718 1850 3722
rect 1814 3688 1818 3692
rect 1830 3678 1834 3682
rect 1874 3703 1878 3707
rect 1881 3703 1885 3707
rect 1894 3698 1898 3702
rect 1926 3868 1930 3872
rect 1942 3858 1946 3862
rect 1926 3848 1930 3852
rect 1918 3688 1922 3692
rect 1950 3848 1954 3852
rect 1942 3818 1946 3822
rect 1934 3758 1938 3762
rect 1966 3808 1970 3812
rect 1958 3758 1962 3762
rect 1942 3728 1946 3732
rect 2030 4098 2034 4102
rect 1998 4088 2002 4092
rect 1982 4058 1986 4062
rect 1990 4038 1994 4042
rect 2006 3988 2010 3992
rect 2014 3948 2018 3952
rect 2022 3938 2026 3942
rect 1990 3928 1994 3932
rect 1998 3878 2002 3882
rect 2038 4078 2042 4082
rect 2102 4158 2106 4162
rect 2238 4318 2242 4322
rect 2230 4308 2234 4312
rect 2222 4278 2226 4282
rect 2174 4268 2178 4272
rect 2214 4268 2218 4272
rect 2158 4248 2162 4252
rect 2134 4148 2138 4152
rect 2110 4138 2114 4142
rect 2078 4128 2082 4132
rect 2110 4128 2114 4132
rect 2086 4118 2090 4122
rect 2102 4078 2106 4082
rect 2190 4248 2194 4252
rect 2254 4248 2258 4252
rect 2206 4238 2210 4242
rect 2190 4208 2194 4212
rect 2198 4188 2202 4192
rect 2190 4168 2194 4172
rect 2174 4148 2178 4152
rect 2198 4148 2202 4152
rect 2246 4148 2250 4152
rect 2334 4528 2338 4532
rect 2350 4528 2354 4532
rect 2374 4518 2378 4522
rect 2398 4518 2402 4522
rect 2366 4478 2370 4482
rect 2382 4478 2386 4482
rect 2326 4368 2330 4372
rect 2326 4358 2330 4362
rect 2286 4338 2290 4342
rect 2318 4278 2322 4282
rect 2358 4418 2362 4422
rect 2406 4468 2410 4472
rect 2382 4458 2386 4462
rect 2390 4438 2394 4442
rect 2478 4738 2482 4742
rect 2422 4728 2426 4732
rect 2430 4728 2434 4732
rect 2454 4728 2458 4732
rect 2438 4718 2442 4722
rect 2438 4708 2442 4712
rect 2430 4688 2434 4692
rect 2462 4688 2466 4692
rect 2462 4668 2466 4672
rect 2454 4558 2458 4562
rect 2486 4668 2490 4672
rect 2478 4598 2482 4602
rect 2534 4748 2538 4752
rect 2534 4728 2538 4732
rect 2534 4678 2538 4682
rect 2558 4738 2562 4742
rect 2582 4738 2586 4742
rect 2558 4688 2562 4692
rect 2622 4848 2626 4852
rect 2630 4838 2634 4842
rect 2638 4758 2642 4762
rect 2614 4748 2618 4752
rect 2630 4748 2634 4752
rect 2606 4738 2610 4742
rect 2638 4738 2642 4742
rect 2606 4728 2610 4732
rect 2662 4708 2666 4712
rect 2654 4688 2658 4692
rect 2638 4678 2642 4682
rect 2590 4668 2594 4672
rect 2526 4658 2530 4662
rect 2494 4648 2498 4652
rect 2518 4648 2522 4652
rect 2518 4638 2522 4642
rect 2534 4598 2538 4602
rect 2510 4578 2514 4582
rect 2510 4568 2514 4572
rect 2486 4548 2490 4552
rect 2470 4538 2474 4542
rect 2454 4498 2458 4502
rect 2422 4428 2426 4432
rect 2414 4408 2418 4412
rect 2386 4403 2390 4407
rect 2393 4403 2397 4407
rect 2430 4388 2434 4392
rect 2374 4378 2378 4382
rect 2390 4378 2394 4382
rect 2414 4368 2418 4372
rect 2342 4348 2346 4352
rect 2366 4348 2370 4352
rect 2278 4248 2282 4252
rect 2334 4218 2338 4222
rect 2302 4188 2306 4192
rect 2366 4338 2370 4342
rect 2422 4338 2426 4342
rect 2478 4468 2482 4472
rect 2462 4428 2466 4432
rect 2446 4388 2450 4392
rect 2454 4378 2458 4382
rect 2446 4358 2450 4362
rect 2494 4388 2498 4392
rect 2478 4368 2482 4372
rect 2478 4358 2482 4362
rect 2534 4468 2538 4472
rect 2526 4448 2530 4452
rect 2582 4658 2586 4662
rect 2574 4648 2578 4652
rect 2590 4618 2594 4622
rect 2574 4578 2578 4582
rect 2590 4558 2594 4562
rect 2558 4528 2562 4532
rect 2622 4648 2626 4652
rect 2646 4668 2650 4672
rect 2678 4828 2682 4832
rect 2750 4918 2754 4922
rect 2878 4938 2882 4942
rect 2798 4928 2802 4932
rect 2878 4918 2882 4922
rect 2890 4903 2894 4907
rect 2897 4903 2901 4907
rect 2854 4878 2858 4882
rect 2790 4858 2794 4862
rect 2862 4858 2866 4862
rect 2710 4748 2714 4752
rect 2830 4788 2834 4792
rect 2902 4848 2906 4852
rect 2878 4778 2882 4782
rect 2894 4778 2898 4782
rect 2798 4748 2802 4752
rect 2854 4748 2858 4752
rect 2902 4738 2906 4742
rect 2862 4728 2866 4732
rect 2870 4728 2874 4732
rect 2894 4728 2898 4732
rect 2886 4718 2890 4722
rect 2846 4708 2850 4712
rect 2890 4703 2894 4707
rect 2897 4703 2901 4707
rect 2942 5008 2946 5012
rect 2926 4968 2930 4972
rect 2926 4938 2930 4942
rect 2918 4878 2922 4882
rect 2942 4948 2946 4952
rect 2942 4928 2946 4932
rect 2966 5028 2970 5032
rect 2998 5028 3002 5032
rect 2958 5018 2962 5022
rect 2966 4938 2970 4942
rect 2966 4888 2970 4892
rect 2958 4868 2962 4872
rect 2934 4838 2938 4842
rect 2950 4838 2954 4842
rect 2918 4818 2922 4822
rect 2926 4818 2930 4822
rect 2862 4678 2866 4682
rect 2910 4678 2914 4682
rect 2870 4668 2874 4672
rect 2702 4658 2706 4662
rect 2734 4658 2738 4662
rect 2814 4658 2818 4662
rect 2854 4658 2858 4662
rect 2958 4788 2962 4792
rect 2926 4758 2930 4762
rect 2982 4888 2986 4892
rect 2982 4868 2986 4872
rect 3070 5058 3074 5062
rect 3054 5048 3058 5052
rect 3038 5018 3042 5022
rect 3126 5038 3130 5042
rect 3086 5028 3090 5032
rect 3046 4978 3050 4982
rect 3054 4978 3058 4982
rect 3110 4968 3114 4972
rect 3118 4958 3122 4962
rect 3126 4958 3130 4962
rect 3006 4948 3010 4952
rect 3078 4938 3082 4942
rect 3126 4938 3130 4942
rect 3110 4928 3114 4932
rect 3198 5058 3202 5062
rect 3158 5048 3162 5052
rect 3174 5048 3178 5052
rect 3166 5038 3170 5042
rect 3182 5038 3186 5042
rect 3198 5038 3202 5042
rect 3166 5018 3170 5022
rect 3150 4988 3154 4992
rect 3150 4978 3154 4982
rect 3142 4908 3146 4912
rect 3070 4898 3074 4902
rect 3022 4888 3026 4892
rect 3022 4878 3026 4882
rect 3134 4888 3138 4892
rect 3030 4868 3034 4872
rect 3054 4868 3058 4872
rect 3078 4858 3082 4862
rect 3118 4858 3122 4862
rect 2982 4768 2986 4772
rect 2990 4738 2994 4742
rect 2974 4728 2978 4732
rect 2934 4688 2938 4692
rect 3022 4708 3026 4712
rect 2926 4678 2930 4682
rect 2926 4668 2930 4672
rect 2670 4598 2674 4602
rect 2678 4538 2682 4542
rect 2638 4508 2642 4512
rect 2614 4498 2618 4502
rect 2686 4498 2690 4502
rect 2686 4478 2690 4482
rect 2630 4458 2634 4462
rect 2542 4418 2546 4422
rect 2598 4448 2602 4452
rect 2558 4408 2562 4412
rect 2534 4368 2538 4372
rect 2502 4348 2506 4352
rect 2518 4348 2522 4352
rect 2526 4348 2530 4352
rect 2510 4338 2514 4342
rect 2350 4278 2354 4282
rect 2430 4278 2434 4282
rect 2502 4318 2506 4322
rect 2486 4308 2490 4312
rect 2462 4298 2466 4302
rect 2462 4278 2466 4282
rect 2366 4268 2370 4272
rect 2430 4268 2434 4272
rect 2438 4268 2442 4272
rect 2446 4268 2450 4272
rect 2470 4268 2474 4272
rect 2486 4268 2490 4272
rect 2438 4248 2442 4252
rect 2382 4238 2386 4242
rect 2386 4203 2390 4207
rect 2393 4203 2397 4207
rect 2406 4168 2410 4172
rect 2310 4148 2314 4152
rect 2190 4138 2194 4142
rect 2206 4138 2210 4142
rect 2166 4098 2170 4102
rect 2150 4058 2154 4062
rect 2326 4128 2330 4132
rect 2342 4108 2346 4112
rect 2230 4078 2234 4082
rect 2238 4078 2242 4082
rect 2334 4078 2338 4082
rect 2510 4258 2514 4262
rect 2486 4238 2490 4242
rect 2510 4218 2514 4222
rect 2470 4198 2474 4202
rect 2462 4178 2466 4182
rect 2454 4148 2458 4152
rect 2358 4138 2362 4142
rect 2430 4138 2434 4142
rect 2398 4118 2402 4122
rect 2486 4118 2490 4122
rect 2366 4108 2370 4112
rect 2366 4098 2370 4102
rect 2430 4098 2434 4102
rect 2406 4078 2410 4082
rect 2302 4058 2306 4062
rect 2422 4058 2426 4062
rect 2086 4038 2090 4042
rect 2102 4038 2106 4042
rect 2054 4028 2058 4032
rect 2078 3998 2082 4002
rect 2046 3948 2050 3952
rect 2038 3938 2042 3942
rect 2054 3938 2058 3942
rect 2118 4008 2122 4012
rect 2094 3988 2098 3992
rect 2142 4038 2146 4042
rect 2126 3968 2130 3972
rect 2134 3968 2138 3972
rect 2118 3958 2122 3962
rect 2126 3958 2130 3962
rect 2134 3958 2138 3962
rect 2086 3928 2090 3932
rect 2158 3948 2162 3952
rect 2166 3948 2170 3952
rect 2070 3878 2074 3882
rect 2102 3878 2106 3882
rect 2046 3868 2050 3872
rect 2014 3858 2018 3862
rect 2038 3858 2042 3862
rect 2086 3858 2090 3862
rect 2102 3858 2106 3862
rect 1990 3848 1994 3852
rect 2070 3848 2074 3852
rect 2078 3848 2082 3852
rect 2110 3848 2114 3852
rect 2126 3818 2130 3822
rect 2166 3888 2170 3892
rect 2150 3868 2154 3872
rect 2150 3848 2154 3852
rect 2110 3808 2114 3812
rect 2094 3798 2098 3802
rect 2030 3788 2034 3792
rect 1990 3758 1994 3762
rect 2126 3768 2130 3772
rect 2158 3778 2162 3782
rect 1982 3748 1986 3752
rect 2086 3748 2090 3752
rect 2118 3748 2122 3752
rect 2142 3748 2146 3752
rect 2158 3748 2162 3752
rect 1966 3738 1970 3742
rect 1958 3728 1962 3732
rect 1950 3708 1954 3712
rect 1934 3678 1938 3682
rect 1894 3668 1898 3672
rect 1926 3668 1930 3672
rect 1854 3658 1858 3662
rect 1822 3648 1826 3652
rect 1838 3598 1842 3602
rect 1838 3568 1842 3572
rect 1814 3548 1818 3552
rect 1806 3508 1810 3512
rect 1830 3508 1834 3512
rect 1582 3468 1586 3472
rect 1590 3468 1594 3472
rect 1678 3468 1682 3472
rect 1798 3468 1802 3472
rect 1590 3458 1594 3462
rect 1598 3458 1602 3462
rect 1590 3448 1594 3452
rect 1590 3408 1594 3412
rect 1574 3358 1578 3362
rect 1582 3358 1586 3362
rect 1606 3378 1610 3382
rect 1598 3358 1602 3362
rect 1558 3318 1562 3322
rect 1566 3308 1570 3312
rect 1574 3298 1578 3302
rect 1558 3288 1562 3292
rect 1446 3248 1450 3252
rect 1470 3248 1474 3252
rect 1502 3248 1506 3252
rect 1486 3238 1490 3242
rect 1478 3228 1482 3232
rect 1502 3228 1506 3232
rect 1278 3198 1282 3202
rect 1246 3158 1250 3162
rect 1190 3148 1194 3152
rect 1102 3138 1106 3142
rect 1158 3138 1162 3142
rect 1182 3138 1186 3142
rect 1206 3138 1210 3142
rect 1238 3138 1242 3142
rect 1078 3128 1082 3132
rect 1142 3128 1146 3132
rect 1062 3108 1066 3112
rect 1070 3098 1074 3102
rect 846 3078 850 3082
rect 942 3078 946 3082
rect 966 3078 970 3082
rect 1038 3078 1042 3082
rect 870 3059 874 3063
rect 1062 3068 1066 3072
rect 1286 3138 1290 3142
rect 1254 3128 1258 3132
rect 1246 3118 1250 3122
rect 1174 3078 1178 3082
rect 1158 3068 1162 3072
rect 1182 3068 1186 3072
rect 1006 3058 1010 3062
rect 1038 3058 1042 3062
rect 1134 3058 1138 3062
rect 1166 3058 1170 3062
rect 1102 3048 1106 3052
rect 934 3038 938 3042
rect 926 3008 930 3012
rect 942 2958 946 2962
rect 1078 3028 1082 3032
rect 1070 2978 1074 2982
rect 1230 3058 1234 3062
rect 1354 3203 1358 3207
rect 1361 3203 1365 3207
rect 1342 3178 1346 3182
rect 1382 3178 1386 3182
rect 1390 3178 1394 3182
rect 1414 3168 1418 3172
rect 1478 3168 1482 3172
rect 1390 3158 1394 3162
rect 1406 3158 1410 3162
rect 1438 3158 1442 3162
rect 1454 3158 1458 3162
rect 1486 3158 1490 3162
rect 1350 3138 1354 3142
rect 1286 3098 1290 3102
rect 1310 3098 1314 3102
rect 1278 3088 1282 3092
rect 1334 3078 1338 3082
rect 1342 3068 1346 3072
rect 1326 3058 1330 3062
rect 1198 3048 1202 3052
rect 1270 3048 1274 3052
rect 1142 2998 1146 3002
rect 1158 2958 1162 2962
rect 862 2948 866 2952
rect 902 2948 906 2952
rect 1142 2948 1146 2952
rect 878 2928 882 2932
rect 870 2918 874 2922
rect 850 2903 854 2907
rect 857 2903 861 2907
rect 870 2868 874 2872
rect 854 2838 858 2842
rect 830 2788 834 2792
rect 854 2758 858 2762
rect 910 2898 914 2902
rect 894 2848 898 2852
rect 918 2848 922 2852
rect 886 2828 890 2832
rect 862 2718 866 2722
rect 850 2703 854 2707
rect 857 2703 861 2707
rect 854 2688 858 2692
rect 814 2668 818 2672
rect 830 2668 834 2672
rect 782 2628 786 2632
rect 806 2648 810 2652
rect 838 2648 842 2652
rect 790 2618 794 2622
rect 822 2618 826 2622
rect 710 2568 714 2572
rect 766 2538 770 2542
rect 750 2528 754 2532
rect 742 2478 746 2482
rect 670 2458 674 2462
rect 702 2468 706 2472
rect 718 2468 722 2472
rect 726 2468 730 2472
rect 750 2468 754 2472
rect 630 2448 634 2452
rect 654 2438 658 2442
rect 814 2568 818 2572
rect 798 2558 802 2562
rect 830 2578 834 2582
rect 830 2568 834 2572
rect 846 2558 850 2562
rect 830 2538 834 2542
rect 806 2528 810 2532
rect 822 2528 826 2532
rect 790 2508 794 2512
rect 710 2438 714 2442
rect 702 2418 706 2422
rect 670 2408 674 2412
rect 630 2388 634 2392
rect 774 2438 778 2442
rect 758 2428 762 2432
rect 758 2408 762 2412
rect 734 2388 738 2392
rect 694 2378 698 2382
rect 726 2378 730 2382
rect 678 2368 682 2372
rect 574 2358 578 2362
rect 502 2348 506 2352
rect 534 2348 538 2352
rect 542 2348 546 2352
rect 646 2348 650 2352
rect 662 2348 666 2352
rect 718 2358 722 2362
rect 750 2348 754 2352
rect 526 2338 530 2342
rect 574 2338 578 2342
rect 654 2338 658 2342
rect 766 2338 770 2342
rect 782 2338 786 2342
rect 478 2328 482 2332
rect 654 2328 658 2332
rect 702 2328 706 2332
rect 470 2308 474 2312
rect 462 2288 466 2292
rect 550 2288 554 2292
rect 598 2268 602 2272
rect 238 2158 242 2162
rect 254 2098 258 2102
rect 286 2138 290 2142
rect 286 2118 290 2122
rect 294 2078 298 2082
rect 254 2068 258 2072
rect 270 2068 274 2072
rect 190 2058 194 2062
rect 182 2048 186 2052
rect 222 2048 226 2052
rect 198 2038 202 2042
rect 190 1998 194 2002
rect 174 1988 178 1992
rect 126 1948 130 1952
rect 182 1948 186 1952
rect 238 2048 242 2052
rect 230 2018 234 2022
rect 262 2018 266 2022
rect 230 1958 234 1962
rect 254 1958 258 1962
rect 318 2248 322 2252
rect 446 2248 450 2252
rect 494 2248 498 2252
rect 382 2228 386 2232
rect 330 2203 334 2207
rect 337 2203 341 2207
rect 358 2188 362 2192
rect 358 2178 362 2182
rect 334 2158 338 2162
rect 350 2158 354 2162
rect 310 2118 314 2122
rect 342 2098 346 2102
rect 310 2048 314 2052
rect 526 2218 530 2222
rect 542 2218 546 2222
rect 574 2218 578 2222
rect 614 2208 618 2212
rect 726 2298 730 2302
rect 710 2288 714 2292
rect 678 2268 682 2272
rect 758 2278 762 2282
rect 718 2268 722 2272
rect 782 2268 786 2272
rect 798 2458 802 2462
rect 934 2898 938 2902
rect 1310 3048 1314 3052
rect 1366 3048 1370 3052
rect 1302 3038 1306 3042
rect 1294 3018 1298 3022
rect 1286 2998 1290 3002
rect 1354 3003 1358 3007
rect 1361 3003 1365 3007
rect 1318 2968 1322 2972
rect 1342 2968 1346 2972
rect 1270 2958 1274 2962
rect 1262 2948 1266 2952
rect 1054 2938 1058 2942
rect 1102 2938 1106 2942
rect 1142 2938 1146 2942
rect 1190 2938 1194 2942
rect 1254 2938 1258 2942
rect 1118 2928 1122 2932
rect 1254 2928 1258 2932
rect 1310 2928 1314 2932
rect 1334 2938 1338 2942
rect 1358 2938 1362 2942
rect 1350 2928 1354 2932
rect 1318 2918 1322 2922
rect 1014 2908 1018 2912
rect 1038 2908 1042 2912
rect 942 2888 946 2892
rect 1262 2908 1266 2912
rect 1086 2898 1090 2902
rect 1038 2888 1042 2892
rect 1078 2888 1082 2892
rect 1126 2888 1130 2892
rect 1246 2888 1250 2892
rect 974 2878 978 2882
rect 998 2878 1002 2882
rect 966 2868 970 2872
rect 1038 2868 1042 2872
rect 926 2838 930 2842
rect 1078 2848 1082 2852
rect 1094 2848 1098 2852
rect 966 2828 970 2832
rect 958 2808 962 2812
rect 894 2798 898 2802
rect 982 2798 986 2802
rect 942 2758 946 2762
rect 958 2758 962 2762
rect 902 2748 906 2752
rect 934 2748 938 2752
rect 894 2738 898 2742
rect 902 2698 906 2702
rect 886 2678 890 2682
rect 926 2738 930 2742
rect 918 2728 922 2732
rect 942 2718 946 2722
rect 934 2678 938 2682
rect 910 2658 914 2662
rect 1006 2758 1010 2762
rect 1094 2798 1098 2802
rect 1134 2868 1138 2872
rect 1190 2868 1194 2872
rect 1110 2848 1114 2852
rect 1150 2838 1154 2842
rect 1118 2808 1122 2812
rect 1142 2808 1146 2812
rect 1070 2788 1074 2792
rect 1102 2788 1106 2792
rect 1086 2758 1090 2762
rect 1118 2758 1122 2762
rect 1070 2748 1074 2752
rect 1078 2738 1082 2742
rect 1054 2708 1058 2712
rect 990 2698 994 2702
rect 950 2668 954 2672
rect 1070 2678 1074 2682
rect 1078 2678 1082 2682
rect 1022 2668 1026 2672
rect 1062 2668 1066 2672
rect 1158 2798 1162 2802
rect 1302 2898 1306 2902
rect 1374 2908 1378 2912
rect 1326 2888 1330 2892
rect 1286 2868 1290 2872
rect 1302 2868 1306 2872
rect 1294 2848 1298 2852
rect 1302 2848 1306 2852
rect 1310 2828 1314 2832
rect 1174 2768 1178 2772
rect 1270 2768 1274 2772
rect 1294 2768 1298 2772
rect 1150 2758 1154 2762
rect 1134 2748 1138 2752
rect 1150 2748 1154 2752
rect 1190 2758 1194 2762
rect 1110 2738 1114 2742
rect 1102 2728 1106 2732
rect 1126 2728 1130 2732
rect 1110 2718 1114 2722
rect 1118 2688 1122 2692
rect 1086 2668 1090 2672
rect 1126 2668 1130 2672
rect 918 2648 922 2652
rect 902 2638 906 2642
rect 926 2638 930 2642
rect 878 2568 882 2572
rect 870 2558 874 2562
rect 910 2558 914 2562
rect 854 2528 858 2532
rect 846 2518 850 2522
rect 850 2503 854 2507
rect 857 2503 861 2507
rect 878 2518 882 2522
rect 822 2468 826 2472
rect 846 2468 850 2472
rect 830 2458 834 2462
rect 838 2398 842 2402
rect 846 2378 850 2382
rect 830 2368 834 2372
rect 854 2318 858 2322
rect 850 2303 854 2307
rect 857 2303 861 2307
rect 806 2268 810 2272
rect 822 2268 826 2272
rect 670 2258 674 2262
rect 702 2258 706 2262
rect 758 2258 762 2262
rect 814 2258 818 2262
rect 686 2248 690 2252
rect 694 2178 698 2182
rect 446 2168 450 2172
rect 662 2158 666 2162
rect 686 2158 690 2162
rect 382 2148 386 2152
rect 790 2248 794 2252
rect 750 2218 754 2222
rect 766 2198 770 2202
rect 838 2238 842 2242
rect 886 2458 890 2462
rect 878 2448 882 2452
rect 894 2438 898 2442
rect 878 2398 882 2402
rect 894 2388 898 2392
rect 918 2468 922 2472
rect 974 2568 978 2572
rect 1014 2568 1018 2572
rect 990 2558 994 2562
rect 1006 2558 1010 2562
rect 974 2548 978 2552
rect 974 2528 978 2532
rect 958 2508 962 2512
rect 990 2468 994 2472
rect 934 2458 938 2462
rect 958 2458 962 2462
rect 926 2448 930 2452
rect 950 2438 954 2442
rect 926 2428 930 2432
rect 902 2358 906 2362
rect 1046 2648 1050 2652
rect 1094 2658 1098 2662
rect 1086 2638 1090 2642
rect 1086 2628 1090 2632
rect 1078 2568 1082 2572
rect 1062 2558 1066 2562
rect 1030 2538 1034 2542
rect 1062 2538 1066 2542
rect 1022 2518 1026 2522
rect 1022 2488 1026 2492
rect 982 2458 986 2462
rect 1006 2458 1010 2462
rect 1030 2468 1034 2472
rect 1062 2468 1066 2472
rect 1054 2458 1058 2462
rect 1102 2638 1106 2642
rect 1102 2538 1106 2542
rect 1094 2518 1098 2522
rect 1078 2508 1082 2512
rect 1070 2448 1074 2452
rect 990 2438 994 2442
rect 966 2388 970 2392
rect 1046 2438 1050 2442
rect 1054 2438 1058 2442
rect 1070 2438 1074 2442
rect 998 2378 1002 2382
rect 1022 2378 1026 2382
rect 934 2368 938 2372
rect 934 2348 938 2352
rect 910 2338 914 2342
rect 942 2338 946 2342
rect 1054 2398 1058 2402
rect 1038 2358 1042 2362
rect 1022 2348 1026 2352
rect 982 2328 986 2332
rect 886 2318 890 2322
rect 902 2318 906 2322
rect 982 2318 986 2322
rect 990 2298 994 2302
rect 1014 2318 1018 2322
rect 918 2268 922 2272
rect 990 2268 994 2272
rect 998 2268 1002 2272
rect 894 2259 898 2263
rect 958 2238 962 2242
rect 870 2228 874 2232
rect 790 2218 794 2222
rect 750 2188 754 2192
rect 974 2248 978 2252
rect 974 2208 978 2212
rect 982 2208 986 2212
rect 1046 2268 1050 2272
rect 1062 2358 1066 2362
rect 1190 2718 1194 2722
rect 1142 2698 1146 2702
rect 1150 2688 1154 2692
rect 1142 2668 1146 2672
rect 1134 2658 1138 2662
rect 1142 2628 1146 2632
rect 1134 2558 1138 2562
rect 1126 2538 1130 2542
rect 1198 2708 1202 2712
rect 1254 2708 1258 2712
rect 1166 2668 1170 2672
rect 1150 2558 1154 2562
rect 1270 2688 1274 2692
rect 1206 2668 1210 2672
rect 1518 3258 1522 3262
rect 1534 3248 1538 3252
rect 1590 3318 1594 3322
rect 1582 3288 1586 3292
rect 1566 3248 1570 3252
rect 1542 3238 1546 3242
rect 1550 3238 1554 3242
rect 1510 3218 1514 3222
rect 1574 3168 1578 3172
rect 1550 3158 1554 3162
rect 1422 3148 1426 3152
rect 1566 3148 1570 3152
rect 1438 3138 1442 3142
rect 1462 3138 1466 3142
rect 1478 3138 1482 3142
rect 1558 3138 1562 3142
rect 1406 3128 1410 3132
rect 1526 3128 1530 3132
rect 1542 3128 1546 3132
rect 1446 3118 1450 3122
rect 1494 3118 1498 3122
rect 1502 3108 1506 3112
rect 1462 3098 1466 3102
rect 1438 3088 1442 3092
rect 1478 3088 1482 3092
rect 1414 3078 1418 3082
rect 1398 3058 1402 3062
rect 1414 3058 1418 3062
rect 1438 3058 1442 3062
rect 1454 3058 1458 3062
rect 1470 3058 1474 3062
rect 1454 3048 1458 3052
rect 1486 3048 1490 3052
rect 1422 3038 1426 3042
rect 1438 3038 1442 3042
rect 1422 3008 1426 3012
rect 1390 2998 1394 3002
rect 1462 2988 1466 2992
rect 1590 3248 1594 3252
rect 1590 3178 1594 3182
rect 1646 3448 1650 3452
rect 1630 3388 1634 3392
rect 1622 3328 1626 3332
rect 1614 3308 1618 3312
rect 1646 3358 1650 3362
rect 1662 3358 1666 3362
rect 1646 3288 1650 3292
rect 1622 3278 1626 3282
rect 1606 3268 1610 3272
rect 1606 3238 1610 3242
rect 1614 3198 1618 3202
rect 1606 3148 1610 3152
rect 1854 3548 1858 3552
rect 1886 3608 1890 3612
rect 1990 3738 1994 3742
rect 2022 3728 2026 3732
rect 1990 3708 1994 3712
rect 2014 3708 2018 3712
rect 1998 3688 2002 3692
rect 1902 3648 1906 3652
rect 1926 3648 1930 3652
rect 1990 3658 1994 3662
rect 1974 3608 1978 3612
rect 2038 3738 2042 3742
rect 2110 3738 2114 3742
rect 2126 3728 2130 3732
rect 2150 3728 2154 3732
rect 2134 3718 2138 3722
rect 2030 3698 2034 3702
rect 2038 3698 2042 3702
rect 2078 3698 2082 3702
rect 2110 3698 2114 3702
rect 2118 3698 2122 3702
rect 2102 3668 2106 3672
rect 2158 3668 2162 3672
rect 2022 3658 2026 3662
rect 2062 3658 2066 3662
rect 2110 3658 2114 3662
rect 2150 3658 2154 3662
rect 1998 3568 2002 3572
rect 1982 3558 1986 3562
rect 2030 3558 2034 3562
rect 1966 3548 1970 3552
rect 1974 3548 1978 3552
rect 1998 3548 2002 3552
rect 2030 3548 2034 3552
rect 1902 3538 1906 3542
rect 1870 3528 1874 3532
rect 1874 3503 1878 3507
rect 1881 3503 1885 3507
rect 1918 3498 1922 3502
rect 1902 3488 1906 3492
rect 1854 3478 1858 3482
rect 1870 3468 1874 3472
rect 1918 3468 1922 3472
rect 1974 3468 1978 3472
rect 1718 3458 1722 3462
rect 1750 3458 1754 3462
rect 1774 3458 1778 3462
rect 1790 3458 1794 3462
rect 1806 3458 1810 3462
rect 1902 3458 1906 3462
rect 1846 3448 1850 3452
rect 1766 3438 1770 3442
rect 1854 3398 1858 3402
rect 1790 3378 1794 3382
rect 1822 3378 1826 3382
rect 1766 3368 1770 3372
rect 1710 3358 1714 3362
rect 1766 3358 1770 3362
rect 1726 3288 1730 3292
rect 1758 3288 1762 3292
rect 1718 3268 1722 3272
rect 1758 3268 1762 3272
rect 1814 3368 1818 3372
rect 1798 3358 1802 3362
rect 1958 3459 1962 3463
rect 1990 3538 1994 3542
rect 2014 3538 2018 3542
rect 2030 3528 2034 3532
rect 2030 3508 2034 3512
rect 2126 3638 2130 3642
rect 2086 3628 2090 3632
rect 2110 3588 2114 3592
rect 2454 4078 2458 4082
rect 2462 4078 2466 4082
rect 2446 4058 2450 4062
rect 2302 4048 2306 4052
rect 2318 4048 2322 4052
rect 2342 4048 2346 4052
rect 2382 4038 2386 4042
rect 2414 4028 2418 4032
rect 2206 4018 2210 4022
rect 2214 4018 2218 4022
rect 2198 3968 2202 3972
rect 2190 3958 2194 3962
rect 2182 3948 2186 3952
rect 2190 3928 2194 3932
rect 2174 3798 2178 3802
rect 2182 3788 2186 3792
rect 2310 3988 2314 3992
rect 2222 3968 2226 3972
rect 2294 3968 2298 3972
rect 2230 3948 2234 3952
rect 2246 3938 2250 3942
rect 2230 3928 2234 3932
rect 2334 3978 2338 3982
rect 2334 3958 2338 3962
rect 2334 3938 2338 3942
rect 2358 3928 2362 3932
rect 2326 3908 2330 3912
rect 2222 3878 2226 3882
rect 2286 3888 2290 3892
rect 2318 3888 2322 3892
rect 2278 3878 2282 3882
rect 2270 3858 2274 3862
rect 2214 3848 2218 3852
rect 2254 3848 2258 3852
rect 2262 3848 2266 3852
rect 2246 3838 2250 3842
rect 2302 3848 2306 3852
rect 2310 3758 2314 3762
rect 2350 3868 2354 3872
rect 2386 4003 2390 4007
rect 2393 4003 2397 4007
rect 2374 3978 2378 3982
rect 2422 3968 2426 3972
rect 2398 3948 2402 3952
rect 2494 4058 2498 4062
rect 2510 4018 2514 4022
rect 2478 3988 2482 3992
rect 2486 3958 2490 3962
rect 2430 3938 2434 3942
rect 2438 3938 2442 3942
rect 2470 3928 2474 3932
rect 2382 3888 2386 3892
rect 2414 3878 2418 3882
rect 2438 3878 2442 3882
rect 2414 3868 2418 3872
rect 2382 3858 2386 3862
rect 2342 3818 2346 3822
rect 2334 3758 2338 3762
rect 2246 3738 2250 3742
rect 2206 3708 2210 3712
rect 2262 3698 2266 3702
rect 2222 3688 2226 3692
rect 2246 3668 2250 3672
rect 2174 3578 2178 3582
rect 2054 3558 2058 3562
rect 2134 3558 2138 3562
rect 2166 3558 2170 3562
rect 2062 3548 2066 3552
rect 2094 3548 2098 3552
rect 2102 3538 2106 3542
rect 2054 3528 2058 3532
rect 2046 3518 2050 3522
rect 2110 3528 2114 3532
rect 2142 3538 2146 3542
rect 2174 3538 2178 3542
rect 2086 3518 2090 3522
rect 2126 3518 2130 3522
rect 2062 3498 2066 3502
rect 2006 3488 2010 3492
rect 2038 3468 2042 3472
rect 2086 3508 2090 3512
rect 1982 3458 1986 3462
rect 1830 3358 1834 3362
rect 1918 3358 1922 3362
rect 1934 3358 1938 3362
rect 1774 3338 1778 3342
rect 1782 3268 1786 3272
rect 1670 3248 1674 3252
rect 1702 3248 1706 3252
rect 1702 3228 1706 3232
rect 1670 3208 1674 3212
rect 1630 3148 1634 3152
rect 1638 3138 1642 3142
rect 1598 3128 1602 3132
rect 1582 3108 1586 3112
rect 1574 3098 1578 3102
rect 1606 3098 1610 3102
rect 1574 3088 1578 3092
rect 1582 3088 1586 3092
rect 1550 3078 1554 3082
rect 1558 3078 1562 3082
rect 1526 3028 1530 3032
rect 1518 2968 1522 2972
rect 1462 2948 1466 2952
rect 1406 2938 1410 2942
rect 1422 2938 1426 2942
rect 1390 2888 1394 2892
rect 1590 3078 1594 3082
rect 1598 3058 1602 3062
rect 1582 3028 1586 3032
rect 1606 3038 1610 3042
rect 1606 3028 1610 3032
rect 1630 3128 1634 3132
rect 1662 3148 1666 3152
rect 1654 3138 1658 3142
rect 1670 3138 1674 3142
rect 1734 3198 1738 3202
rect 1702 3188 1706 3192
rect 1846 3328 1850 3332
rect 1822 3308 1826 3312
rect 1830 3278 1834 3282
rect 1822 3268 1826 3272
rect 1846 3248 1850 3252
rect 1822 3218 1826 3222
rect 1806 3208 1810 3212
rect 1790 3198 1794 3202
rect 1782 3188 1786 3192
rect 1694 3178 1698 3182
rect 1774 3168 1778 3172
rect 1694 3158 1698 3162
rect 1710 3158 1714 3162
rect 1806 3158 1810 3162
rect 1662 3078 1666 3082
rect 1622 3058 1626 3062
rect 1622 3038 1626 3042
rect 1614 2998 1618 3002
rect 1630 2988 1634 2992
rect 1742 3148 1746 3152
rect 1774 3148 1778 3152
rect 1894 3318 1898 3322
rect 1874 3303 1878 3307
rect 1881 3303 1885 3307
rect 1894 3288 1898 3292
rect 1918 3288 1922 3292
rect 1910 3278 1914 3282
rect 1870 3238 1874 3242
rect 1870 3218 1874 3222
rect 1862 3208 1866 3212
rect 2038 3438 2042 3442
rect 2150 3528 2154 3532
rect 2102 3418 2106 3422
rect 2110 3378 2114 3382
rect 2014 3368 2018 3372
rect 2030 3368 2034 3372
rect 1958 3358 1962 3362
rect 1982 3358 1986 3362
rect 1966 3348 1970 3352
rect 1950 3338 1954 3342
rect 1974 3328 1978 3332
rect 1958 3248 1962 3252
rect 1934 3188 1938 3192
rect 1902 3158 1906 3162
rect 2054 3358 2058 3362
rect 1998 3348 2002 3352
rect 2006 3338 2010 3342
rect 2038 3338 2042 3342
rect 2030 3288 2034 3292
rect 2046 3278 2050 3282
rect 2030 3258 2034 3262
rect 2006 3218 2010 3222
rect 1998 3178 2002 3182
rect 2014 3178 2018 3182
rect 1990 3158 1994 3162
rect 1942 3148 1946 3152
rect 1806 3138 1810 3142
rect 1846 3138 1850 3142
rect 1982 3138 1986 3142
rect 1798 3128 1802 3132
rect 2014 3118 2018 3122
rect 1798 3108 1802 3112
rect 1950 3108 1954 3112
rect 2038 3248 2042 3252
rect 2046 3228 2050 3232
rect 2078 3338 2082 3342
rect 2102 3338 2106 3342
rect 2102 3308 2106 3312
rect 2142 3488 2146 3492
rect 2142 3428 2146 3432
rect 2174 3458 2178 3462
rect 2166 3408 2170 3412
rect 2158 3398 2162 3402
rect 2142 3368 2146 3372
rect 2126 3338 2130 3342
rect 2166 3338 2170 3342
rect 2134 3318 2138 3322
rect 2094 3238 2098 3242
rect 2110 3238 2114 3242
rect 2070 3218 2074 3222
rect 2062 3188 2066 3192
rect 2038 3178 2042 3182
rect 2070 3168 2074 3172
rect 2078 3168 2082 3172
rect 1874 3103 1878 3107
rect 1881 3103 1885 3107
rect 1822 3098 1826 3102
rect 1934 3098 1938 3102
rect 1726 3078 1730 3082
rect 1846 3078 1850 3082
rect 1934 3078 1938 3082
rect 1694 3068 1698 3072
rect 1886 3068 1890 3072
rect 1918 3068 1922 3072
rect 1654 2998 1658 3002
rect 1646 2968 1650 2972
rect 1838 3058 1842 3062
rect 1702 3048 1706 3052
rect 1726 3048 1730 3052
rect 1678 3028 1682 3032
rect 1686 3018 1690 3022
rect 1678 2968 1682 2972
rect 1582 2948 1586 2952
rect 1718 2948 1722 2952
rect 1574 2938 1578 2942
rect 1662 2938 1666 2942
rect 1526 2928 1530 2932
rect 1534 2928 1538 2932
rect 1486 2898 1490 2902
rect 1422 2878 1426 2882
rect 1438 2878 1442 2882
rect 1406 2868 1410 2872
rect 1390 2848 1394 2852
rect 1382 2838 1386 2842
rect 1510 2878 1514 2882
rect 1454 2868 1458 2872
rect 1598 2898 1602 2902
rect 1582 2888 1586 2892
rect 1622 2868 1626 2872
rect 1438 2848 1442 2852
rect 1558 2848 1562 2852
rect 1438 2838 1442 2842
rect 1566 2838 1570 2842
rect 1422 2828 1426 2832
rect 1354 2803 1358 2807
rect 1361 2803 1365 2807
rect 1406 2808 1410 2812
rect 1422 2808 1426 2812
rect 1398 2788 1402 2792
rect 1350 2758 1354 2762
rect 1366 2728 1370 2732
rect 1374 2728 1378 2732
rect 1334 2688 1338 2692
rect 1326 2668 1330 2672
rect 1350 2668 1354 2672
rect 1302 2658 1306 2662
rect 1182 2638 1186 2642
rect 1198 2548 1202 2552
rect 1390 2698 1394 2702
rect 1382 2668 1386 2672
rect 1342 2638 1346 2642
rect 1350 2638 1354 2642
rect 1302 2618 1306 2622
rect 1318 2618 1322 2622
rect 1294 2558 1298 2562
rect 1310 2558 1314 2562
rect 1354 2603 1358 2607
rect 1361 2603 1365 2607
rect 1382 2558 1386 2562
rect 1334 2548 1338 2552
rect 1166 2538 1170 2542
rect 1174 2538 1178 2542
rect 1190 2538 1194 2542
rect 1206 2538 1210 2542
rect 1254 2538 1258 2542
rect 1262 2538 1266 2542
rect 1142 2508 1146 2512
rect 1150 2498 1154 2502
rect 1174 2498 1178 2502
rect 1134 2458 1138 2462
rect 1126 2368 1130 2372
rect 1126 2358 1130 2362
rect 1126 2348 1130 2352
rect 1214 2518 1218 2522
rect 1206 2498 1210 2502
rect 1198 2468 1202 2472
rect 1182 2438 1186 2442
rect 1182 2368 1186 2372
rect 1190 2358 1194 2362
rect 1182 2348 1186 2352
rect 1134 2338 1138 2342
rect 1142 2338 1146 2342
rect 1110 2328 1114 2332
rect 1102 2278 1106 2282
rect 1214 2468 1218 2472
rect 1214 2458 1218 2462
rect 1206 2358 1210 2362
rect 1206 2348 1210 2352
rect 1254 2528 1258 2532
rect 1238 2468 1242 2472
rect 1238 2448 1242 2452
rect 1318 2498 1322 2502
rect 1302 2468 1306 2472
rect 1246 2438 1250 2442
rect 1254 2438 1258 2442
rect 1270 2438 1274 2442
rect 1166 2328 1170 2332
rect 1230 2328 1234 2332
rect 1158 2298 1162 2302
rect 1198 2288 1202 2292
rect 1198 2278 1202 2282
rect 1206 2278 1210 2282
rect 1086 2268 1090 2272
rect 1214 2268 1218 2272
rect 1062 2258 1066 2262
rect 1086 2258 1090 2262
rect 1022 2218 1026 2222
rect 1038 2218 1042 2222
rect 1014 2188 1018 2192
rect 966 2178 970 2182
rect 774 2168 778 2172
rect 1046 2168 1050 2172
rect 854 2158 858 2162
rect 422 2138 426 2142
rect 486 2138 490 2142
rect 550 2138 554 2142
rect 670 2138 674 2142
rect 734 2138 738 2142
rect 358 2118 362 2122
rect 350 2038 354 2042
rect 330 2003 334 2007
rect 337 2003 341 2007
rect 318 1998 322 2002
rect 286 1988 290 1992
rect 342 1988 346 1992
rect 286 1968 290 1972
rect 270 1958 274 1962
rect 222 1948 226 1952
rect 254 1948 258 1952
rect 118 1908 122 1912
rect 142 1908 146 1912
rect 102 1888 106 1892
rect 70 1878 74 1882
rect 182 1888 186 1892
rect 150 1868 154 1872
rect 190 1868 194 1872
rect 126 1858 130 1862
rect 70 1848 74 1852
rect 62 1818 66 1822
rect 142 1748 146 1752
rect 14 1738 18 1742
rect 70 1738 74 1742
rect 62 1728 66 1732
rect 54 1658 58 1662
rect 38 1538 42 1542
rect 54 1458 58 1462
rect 158 1728 162 1732
rect 158 1718 162 1722
rect 94 1708 98 1712
rect 134 1708 138 1712
rect 118 1688 122 1692
rect 102 1658 106 1662
rect 110 1648 114 1652
rect 222 1928 226 1932
rect 254 1888 258 1892
rect 278 1948 282 1952
rect 326 1948 330 1952
rect 462 2098 466 2102
rect 390 2078 394 2082
rect 382 2068 386 2072
rect 334 1938 338 1942
rect 286 1918 290 1922
rect 318 1918 322 1922
rect 318 1888 322 1892
rect 262 1878 266 1882
rect 286 1878 290 1882
rect 398 2058 402 2062
rect 638 2108 642 2112
rect 542 2098 546 2102
rect 566 2098 570 2102
rect 574 2098 578 2102
rect 526 2088 530 2092
rect 550 2088 554 2092
rect 558 2088 562 2092
rect 526 2078 530 2082
rect 582 2078 586 2082
rect 606 2058 610 2062
rect 494 2048 498 2052
rect 614 2048 618 2052
rect 638 2048 642 2052
rect 726 2088 730 2092
rect 678 2038 682 2042
rect 710 2038 714 2042
rect 662 2028 666 2032
rect 486 1988 490 1992
rect 470 1978 474 1982
rect 422 1968 426 1972
rect 430 1968 434 1972
rect 758 2098 762 2102
rect 766 2048 770 2052
rect 750 2028 754 2032
rect 758 1988 762 1992
rect 630 1968 634 1972
rect 758 1968 762 1972
rect 654 1958 658 1962
rect 790 2128 794 2132
rect 798 2108 802 2112
rect 790 2078 794 2082
rect 854 2148 858 2152
rect 822 2138 826 2142
rect 934 2158 938 2162
rect 1022 2148 1026 2152
rect 862 2138 866 2142
rect 934 2138 938 2142
rect 846 2118 850 2122
rect 850 2103 854 2107
rect 857 2103 861 2107
rect 838 2088 842 2092
rect 822 2078 826 2082
rect 798 2058 802 2062
rect 806 2058 810 2062
rect 822 2058 826 2062
rect 798 2048 802 2052
rect 822 2048 826 2052
rect 814 2038 818 2042
rect 814 1998 818 2002
rect 782 1968 786 1972
rect 790 1968 794 1972
rect 398 1948 402 1952
rect 398 1928 402 1932
rect 382 1908 386 1912
rect 398 1908 402 1912
rect 422 1908 426 1912
rect 382 1878 386 1882
rect 286 1868 290 1872
rect 374 1868 378 1872
rect 254 1848 258 1852
rect 206 1798 210 1802
rect 238 1798 242 1802
rect 454 1908 458 1912
rect 646 1948 650 1952
rect 766 1948 770 1952
rect 574 1938 578 1942
rect 590 1938 594 1942
rect 646 1928 650 1932
rect 670 1928 674 1932
rect 694 1928 698 1932
rect 502 1918 506 1922
rect 766 1918 770 1922
rect 606 1888 610 1892
rect 614 1878 618 1882
rect 638 1878 642 1882
rect 702 1878 706 1882
rect 750 1878 754 1882
rect 462 1868 466 1872
rect 510 1868 514 1872
rect 694 1868 698 1872
rect 718 1868 722 1872
rect 334 1858 338 1862
rect 350 1858 354 1862
rect 374 1858 378 1862
rect 430 1858 434 1862
rect 510 1858 514 1862
rect 542 1858 546 1862
rect 614 1858 618 1862
rect 686 1858 690 1862
rect 702 1858 706 1862
rect 710 1858 714 1862
rect 286 1808 290 1812
rect 262 1788 266 1792
rect 254 1748 258 1752
rect 286 1748 290 1752
rect 238 1728 242 1732
rect 198 1718 202 1722
rect 166 1678 170 1682
rect 158 1658 162 1662
rect 190 1658 194 1662
rect 142 1648 146 1652
rect 126 1638 130 1642
rect 174 1638 178 1642
rect 494 1838 498 1842
rect 330 1803 334 1807
rect 337 1803 341 1807
rect 358 1748 362 1752
rect 294 1708 298 1712
rect 334 1708 338 1712
rect 254 1698 258 1702
rect 214 1668 218 1672
rect 222 1658 226 1662
rect 214 1648 218 1652
rect 206 1638 210 1642
rect 190 1618 194 1622
rect 102 1568 106 1572
rect 134 1568 138 1572
rect 142 1558 146 1562
rect 166 1558 170 1562
rect 102 1548 106 1552
rect 126 1548 130 1552
rect 110 1538 114 1542
rect 118 1538 122 1542
rect 118 1508 122 1512
rect 94 1478 98 1482
rect 102 1468 106 1472
rect 126 1498 130 1502
rect 134 1478 138 1482
rect 110 1448 114 1452
rect 110 1358 114 1362
rect 70 1328 74 1332
rect 14 1318 18 1322
rect 86 1318 90 1322
rect 38 1268 42 1272
rect 110 1268 114 1272
rect 254 1648 258 1652
rect 254 1568 258 1572
rect 246 1558 250 1562
rect 214 1548 218 1552
rect 246 1548 250 1552
rect 174 1528 178 1532
rect 222 1528 226 1532
rect 166 1478 170 1482
rect 198 1468 202 1472
rect 142 1458 146 1462
rect 158 1458 162 1462
rect 190 1458 194 1462
rect 126 1338 130 1342
rect 174 1448 178 1452
rect 174 1368 178 1372
rect 206 1358 210 1362
rect 198 1348 202 1352
rect 166 1338 170 1342
rect 238 1498 242 1502
rect 350 1658 354 1662
rect 334 1648 338 1652
rect 310 1588 314 1592
rect 270 1578 274 1582
rect 330 1603 334 1607
rect 337 1603 341 1607
rect 318 1578 322 1582
rect 278 1548 282 1552
rect 334 1548 338 1552
rect 230 1458 234 1462
rect 246 1458 250 1462
rect 222 1358 226 1362
rect 214 1318 218 1322
rect 182 1298 186 1302
rect 150 1288 154 1292
rect 182 1288 186 1292
rect 246 1438 250 1442
rect 518 1828 522 1832
rect 430 1778 434 1782
rect 398 1768 402 1772
rect 382 1758 386 1762
rect 422 1758 426 1762
rect 438 1748 442 1752
rect 374 1738 378 1742
rect 414 1738 418 1742
rect 438 1738 442 1742
rect 398 1718 402 1722
rect 390 1708 394 1712
rect 382 1688 386 1692
rect 374 1648 378 1652
rect 398 1688 402 1692
rect 438 1698 442 1702
rect 406 1678 410 1682
rect 422 1678 426 1682
rect 438 1648 442 1652
rect 398 1618 402 1622
rect 382 1608 386 1612
rect 430 1608 434 1612
rect 406 1578 410 1582
rect 422 1578 426 1582
rect 398 1568 402 1572
rect 374 1558 378 1562
rect 382 1558 386 1562
rect 414 1548 418 1552
rect 574 1848 578 1852
rect 550 1828 554 1832
rect 526 1798 530 1802
rect 598 1838 602 1842
rect 526 1778 530 1782
rect 582 1778 586 1782
rect 518 1748 522 1752
rect 510 1738 514 1742
rect 478 1698 482 1702
rect 462 1648 466 1652
rect 478 1648 482 1652
rect 454 1638 458 1642
rect 342 1528 346 1532
rect 366 1528 370 1532
rect 390 1518 394 1522
rect 342 1508 346 1512
rect 326 1498 330 1502
rect 350 1498 354 1502
rect 302 1488 306 1492
rect 310 1488 314 1492
rect 318 1488 322 1492
rect 382 1488 386 1492
rect 302 1478 306 1482
rect 278 1358 282 1362
rect 310 1358 314 1362
rect 270 1348 274 1352
rect 374 1478 378 1482
rect 414 1478 418 1482
rect 390 1468 394 1472
rect 542 1758 546 1762
rect 590 1758 594 1762
rect 590 1748 594 1752
rect 582 1738 586 1742
rect 558 1728 562 1732
rect 590 1698 594 1702
rect 558 1688 562 1692
rect 518 1678 522 1682
rect 542 1678 546 1682
rect 566 1668 570 1672
rect 614 1728 618 1732
rect 670 1808 674 1812
rect 710 1808 714 1812
rect 726 1808 730 1812
rect 766 1858 770 1862
rect 766 1838 770 1842
rect 750 1808 754 1812
rect 830 1978 834 1982
rect 806 1948 810 1952
rect 782 1908 786 1912
rect 774 1808 778 1812
rect 766 1788 770 1792
rect 806 1928 810 1932
rect 1006 2128 1010 2132
rect 878 2088 882 2092
rect 878 2078 882 2082
rect 926 2078 930 2082
rect 934 2078 938 2082
rect 878 2058 882 2062
rect 910 2058 914 2062
rect 958 2058 962 2062
rect 862 1968 866 1972
rect 870 1938 874 1942
rect 862 1928 866 1932
rect 850 1903 854 1907
rect 857 1903 861 1907
rect 838 1898 842 1902
rect 838 1878 842 1882
rect 926 2048 930 2052
rect 950 2038 954 2042
rect 902 2008 906 2012
rect 886 1998 890 2002
rect 902 1988 906 1992
rect 942 1958 946 1962
rect 934 1928 938 1932
rect 814 1868 818 1872
rect 942 1868 946 1872
rect 814 1858 818 1862
rect 878 1858 882 1862
rect 846 1848 850 1852
rect 822 1838 826 1842
rect 854 1828 858 1832
rect 830 1818 834 1822
rect 798 1768 802 1772
rect 758 1758 762 1762
rect 734 1748 738 1752
rect 646 1678 650 1682
rect 606 1668 610 1672
rect 638 1668 642 1672
rect 614 1658 618 1662
rect 646 1658 650 1662
rect 582 1648 586 1652
rect 550 1638 554 1642
rect 590 1638 594 1642
rect 574 1628 578 1632
rect 518 1578 522 1582
rect 614 1628 618 1632
rect 622 1598 626 1602
rect 686 1628 690 1632
rect 654 1618 658 1622
rect 646 1608 650 1612
rect 598 1578 602 1582
rect 606 1578 610 1582
rect 638 1578 642 1582
rect 558 1548 562 1552
rect 590 1548 594 1552
rect 630 1548 634 1552
rect 454 1538 458 1542
rect 438 1528 442 1532
rect 478 1528 482 1532
rect 462 1488 466 1492
rect 446 1478 450 1482
rect 350 1458 354 1462
rect 358 1458 362 1462
rect 446 1458 450 1462
rect 502 1458 506 1462
rect 430 1448 434 1452
rect 438 1448 442 1452
rect 350 1438 354 1442
rect 366 1438 370 1442
rect 330 1403 334 1407
rect 337 1403 341 1407
rect 238 1338 242 1342
rect 262 1338 266 1342
rect 278 1338 282 1342
rect 318 1338 322 1342
rect 238 1318 242 1322
rect 222 1278 226 1282
rect 134 1268 138 1272
rect 102 1258 106 1262
rect 126 1258 130 1262
rect 94 1248 98 1252
rect 142 1248 146 1252
rect 246 1298 250 1302
rect 206 1258 210 1262
rect 254 1258 258 1262
rect 190 1248 194 1252
rect 166 1238 170 1242
rect 158 1228 162 1232
rect 150 1178 154 1182
rect 158 1178 162 1182
rect 94 1168 98 1172
rect 102 1168 106 1172
rect 126 1158 130 1162
rect 166 1158 170 1162
rect 54 1148 58 1152
rect 94 1148 98 1152
rect 126 1148 130 1152
rect 134 1138 138 1142
rect 158 1128 162 1132
rect 78 1118 82 1122
rect 38 1078 42 1082
rect 62 1068 66 1072
rect 38 958 42 962
rect 46 858 50 862
rect 150 1088 154 1092
rect 118 1078 122 1082
rect 126 1078 130 1082
rect 214 1178 218 1182
rect 230 1178 234 1182
rect 182 1168 186 1172
rect 190 1168 194 1172
rect 198 1148 202 1152
rect 230 1138 234 1142
rect 214 1118 218 1122
rect 182 1108 186 1112
rect 158 1078 162 1082
rect 174 1078 178 1082
rect 270 1268 274 1272
rect 286 1258 290 1262
rect 278 1238 282 1242
rect 330 1203 334 1207
rect 337 1203 341 1207
rect 326 1178 330 1182
rect 278 1148 282 1152
rect 262 1138 266 1142
rect 262 1118 266 1122
rect 270 1098 274 1102
rect 262 1068 266 1072
rect 110 1058 114 1062
rect 142 1058 146 1062
rect 174 1058 178 1062
rect 262 1058 266 1062
rect 222 1028 226 1032
rect 206 1018 210 1022
rect 158 998 162 1002
rect 102 968 106 972
rect 118 958 122 962
rect 134 958 138 962
rect 110 938 114 942
rect 182 968 186 972
rect 198 968 202 972
rect 166 958 170 962
rect 150 918 154 922
rect 118 908 122 912
rect 254 968 258 972
rect 262 958 266 962
rect 270 958 274 962
rect 230 948 234 952
rect 166 918 170 922
rect 158 898 162 902
rect 102 888 106 892
rect 150 888 154 892
rect 102 848 106 852
rect 174 878 178 882
rect 182 868 186 872
rect 254 948 258 952
rect 302 1138 306 1142
rect 302 1098 306 1102
rect 294 1078 298 1082
rect 430 1428 434 1432
rect 430 1408 434 1412
rect 406 1398 410 1402
rect 374 1347 378 1351
rect 398 1348 402 1352
rect 414 1348 418 1352
rect 478 1408 482 1412
rect 470 1388 474 1392
rect 486 1388 490 1392
rect 454 1378 458 1382
rect 502 1378 506 1382
rect 494 1348 498 1352
rect 478 1328 482 1332
rect 454 1288 458 1292
rect 486 1288 490 1292
rect 590 1538 594 1542
rect 582 1518 586 1522
rect 590 1518 594 1522
rect 582 1508 586 1512
rect 566 1478 570 1482
rect 686 1608 690 1612
rect 702 1588 706 1592
rect 750 1738 754 1742
rect 790 1748 794 1752
rect 902 1808 906 1812
rect 990 1998 994 2002
rect 982 1958 986 1962
rect 998 1948 1002 1952
rect 966 1938 970 1942
rect 1022 2058 1026 2062
rect 1142 2259 1146 2263
rect 1270 2408 1274 2412
rect 1254 2358 1258 2362
rect 1246 2298 1250 2302
rect 1262 2278 1266 2282
rect 1406 2778 1410 2782
rect 1534 2828 1538 2832
rect 1518 2808 1522 2812
rect 1574 2788 1578 2792
rect 1550 2778 1554 2782
rect 1454 2768 1458 2772
rect 1478 2758 1482 2762
rect 1502 2758 1506 2762
rect 1542 2758 1546 2762
rect 1438 2748 1442 2752
rect 1462 2748 1466 2752
rect 1406 2718 1410 2722
rect 1430 2738 1434 2742
rect 1438 2728 1442 2732
rect 1430 2708 1434 2712
rect 1406 2658 1410 2662
rect 1406 2648 1410 2652
rect 1342 2538 1346 2542
rect 1366 2528 1370 2532
rect 1486 2738 1490 2742
rect 1502 2718 1506 2722
rect 1478 2688 1482 2692
rect 1782 3028 1786 3032
rect 1822 3028 1826 3032
rect 1798 2978 1802 2982
rect 1822 2948 1826 2952
rect 1782 2938 1786 2942
rect 1814 2938 1818 2942
rect 1742 2928 1746 2932
rect 1710 2898 1714 2902
rect 1702 2868 1706 2872
rect 1774 2918 1778 2922
rect 1766 2888 1770 2892
rect 1750 2868 1754 2872
rect 1758 2868 1762 2872
rect 1694 2848 1698 2852
rect 1734 2848 1738 2852
rect 1678 2828 1682 2832
rect 1670 2808 1674 2812
rect 1726 2808 1730 2812
rect 1574 2768 1578 2772
rect 1638 2768 1642 2772
rect 1718 2768 1722 2772
rect 1558 2758 1562 2762
rect 1566 2748 1570 2752
rect 1574 2738 1578 2742
rect 1542 2728 1546 2732
rect 1606 2728 1610 2732
rect 1582 2718 1586 2722
rect 1590 2708 1594 2712
rect 1526 2688 1530 2692
rect 1574 2688 1578 2692
rect 1518 2678 1522 2682
rect 1446 2658 1450 2662
rect 1446 2648 1450 2652
rect 1422 2638 1426 2642
rect 1414 2628 1418 2632
rect 1510 2659 1514 2663
rect 1510 2638 1514 2642
rect 1478 2628 1482 2632
rect 1470 2618 1474 2622
rect 1422 2608 1426 2612
rect 1430 2558 1434 2562
rect 1414 2548 1418 2552
rect 1366 2478 1370 2482
rect 1414 2478 1418 2482
rect 1398 2468 1402 2472
rect 1326 2458 1330 2462
rect 1406 2458 1410 2462
rect 1358 2448 1362 2452
rect 1398 2408 1402 2412
rect 1354 2403 1358 2407
rect 1361 2403 1365 2407
rect 1390 2398 1394 2402
rect 1326 2388 1330 2392
rect 1318 2378 1322 2382
rect 1390 2378 1394 2382
rect 1374 2348 1378 2352
rect 1342 2338 1346 2342
rect 1382 2328 1386 2332
rect 1446 2538 1450 2542
rect 1446 2468 1450 2472
rect 1438 2428 1442 2432
rect 1430 2408 1434 2412
rect 1654 2708 1658 2712
rect 1646 2688 1650 2692
rect 1662 2688 1666 2692
rect 1598 2668 1602 2672
rect 1622 2668 1626 2672
rect 1606 2658 1610 2662
rect 1566 2648 1570 2652
rect 1526 2628 1530 2632
rect 1582 2628 1586 2632
rect 1542 2618 1546 2622
rect 1566 2608 1570 2612
rect 1518 2568 1522 2572
rect 1534 2568 1538 2572
rect 1558 2558 1562 2562
rect 1590 2608 1594 2612
rect 1630 2648 1634 2652
rect 1702 2738 1706 2742
rect 1710 2678 1714 2682
rect 1686 2668 1690 2672
rect 1702 2668 1706 2672
rect 1694 2658 1698 2662
rect 1710 2658 1714 2662
rect 1622 2558 1626 2562
rect 1670 2618 1674 2622
rect 1534 2548 1538 2552
rect 1590 2548 1594 2552
rect 1614 2548 1618 2552
rect 1486 2538 1490 2542
rect 1566 2538 1570 2542
rect 1462 2508 1466 2512
rect 1486 2498 1490 2502
rect 1494 2498 1498 2502
rect 1526 2498 1530 2502
rect 1470 2468 1474 2472
rect 1454 2438 1458 2442
rect 1470 2438 1474 2442
rect 1454 2428 1458 2432
rect 1486 2398 1490 2402
rect 1446 2348 1450 2352
rect 1478 2348 1482 2352
rect 1294 2288 1298 2292
rect 1398 2308 1402 2312
rect 1278 2278 1282 2282
rect 1342 2278 1346 2282
rect 1366 2278 1370 2282
rect 1230 2258 1234 2262
rect 1246 2258 1250 2262
rect 1262 2258 1266 2262
rect 1278 2258 1282 2262
rect 1286 2258 1290 2262
rect 1118 2248 1122 2252
rect 1086 2178 1090 2182
rect 1126 2178 1130 2182
rect 1206 2178 1210 2182
rect 1086 2148 1090 2152
rect 1070 2138 1074 2142
rect 1062 2098 1066 2102
rect 1062 2088 1066 2092
rect 1086 2098 1090 2102
rect 1110 2138 1114 2142
rect 1110 2078 1114 2082
rect 1238 2188 1242 2192
rect 1166 2148 1170 2152
rect 1214 2148 1218 2152
rect 1230 2148 1234 2152
rect 1286 2238 1290 2242
rect 1278 2158 1282 2162
rect 1246 2138 1250 2142
rect 1142 2118 1146 2122
rect 1158 2088 1162 2092
rect 1126 2068 1130 2072
rect 1142 2068 1146 2072
rect 1190 2068 1194 2072
rect 1206 2068 1210 2072
rect 1222 2068 1226 2072
rect 1134 2058 1138 2062
rect 1126 1988 1130 1992
rect 1126 1968 1130 1972
rect 1054 1948 1058 1952
rect 1070 1948 1074 1952
rect 1118 1948 1122 1952
rect 1126 1948 1130 1952
rect 1006 1928 1010 1932
rect 958 1918 962 1922
rect 1118 1938 1122 1942
rect 1022 1898 1026 1902
rect 1022 1888 1026 1892
rect 1030 1868 1034 1872
rect 1086 1928 1090 1932
rect 1078 1898 1082 1902
rect 1070 1888 1074 1892
rect 1062 1868 1066 1872
rect 1046 1858 1050 1862
rect 1038 1818 1042 1822
rect 958 1798 962 1802
rect 910 1758 914 1762
rect 854 1747 858 1751
rect 974 1748 978 1752
rect 1022 1748 1026 1752
rect 806 1738 810 1742
rect 902 1738 906 1742
rect 934 1738 938 1742
rect 766 1718 770 1722
rect 718 1708 722 1712
rect 750 1688 754 1692
rect 782 1688 786 1692
rect 750 1678 754 1682
rect 750 1658 754 1662
rect 758 1638 762 1642
rect 766 1628 770 1632
rect 798 1608 802 1612
rect 710 1568 714 1572
rect 646 1548 650 1552
rect 670 1548 674 1552
rect 654 1538 658 1542
rect 662 1538 666 1542
rect 654 1528 658 1532
rect 654 1488 658 1492
rect 678 1488 682 1492
rect 614 1478 618 1482
rect 614 1458 618 1462
rect 590 1418 594 1422
rect 526 1358 530 1362
rect 558 1358 562 1362
rect 526 1348 530 1352
rect 534 1338 538 1342
rect 622 1338 626 1342
rect 510 1328 514 1332
rect 422 1268 426 1272
rect 438 1268 442 1272
rect 558 1328 562 1332
rect 526 1308 530 1312
rect 614 1278 618 1282
rect 598 1268 602 1272
rect 422 1258 426 1262
rect 374 1248 378 1252
rect 438 1168 442 1172
rect 454 1168 458 1172
rect 406 1158 410 1162
rect 430 1158 434 1162
rect 390 1148 394 1152
rect 374 1098 378 1102
rect 334 1088 338 1092
rect 342 1088 346 1092
rect 294 1048 298 1052
rect 318 1038 322 1042
rect 550 1238 554 1242
rect 494 1158 498 1162
rect 422 1138 426 1142
rect 494 1138 498 1142
rect 398 1128 402 1132
rect 430 1118 434 1122
rect 454 1118 458 1122
rect 438 1078 442 1082
rect 414 1068 418 1072
rect 430 1068 434 1072
rect 374 1058 378 1062
rect 326 1018 330 1022
rect 330 1003 334 1007
rect 337 1003 341 1007
rect 310 968 314 972
rect 326 968 330 972
rect 286 958 290 962
rect 334 958 338 962
rect 350 958 354 962
rect 222 938 226 942
rect 238 938 242 942
rect 286 938 290 942
rect 206 918 210 922
rect 238 888 242 892
rect 246 878 250 882
rect 126 858 130 862
rect 214 858 218 862
rect 110 838 114 842
rect 134 838 138 842
rect 78 828 82 832
rect 38 748 42 752
rect 62 748 66 752
rect 14 738 18 742
rect 30 738 34 742
rect 38 668 42 672
rect 62 668 66 672
rect 118 768 122 772
rect 166 758 170 762
rect 102 748 106 752
rect 118 748 122 752
rect 158 748 162 752
rect 198 758 202 762
rect 206 738 210 742
rect 182 718 186 722
rect 190 718 194 722
rect 174 708 178 712
rect 246 788 250 792
rect 230 748 234 752
rect 230 728 234 732
rect 230 698 234 702
rect 222 688 226 692
rect 126 678 130 682
rect 94 668 98 672
rect 102 668 106 672
rect 134 668 138 672
rect 158 668 162 672
rect 206 668 210 672
rect 54 658 58 662
rect 70 658 74 662
rect 46 648 50 652
rect 54 638 58 642
rect 78 638 82 642
rect 46 488 50 492
rect 14 458 18 462
rect 6 348 10 352
rect 38 318 42 322
rect 6 308 10 312
rect 22 288 26 292
rect 126 658 130 662
rect 174 638 178 642
rect 198 608 202 612
rect 190 598 194 602
rect 134 588 138 592
rect 182 588 186 592
rect 262 768 266 772
rect 294 898 298 902
rect 278 748 282 752
rect 270 718 274 722
rect 262 678 266 682
rect 374 1008 378 1012
rect 342 948 346 952
rect 334 888 338 892
rect 326 858 330 862
rect 350 808 354 812
rect 330 803 334 807
rect 337 803 341 807
rect 318 778 322 782
rect 270 668 274 672
rect 294 668 298 672
rect 302 668 306 672
rect 278 658 282 662
rect 238 568 242 572
rect 126 558 130 562
rect 206 558 210 562
rect 78 548 82 552
rect 62 538 66 542
rect 230 538 234 542
rect 110 528 114 532
rect 206 528 210 532
rect 126 508 130 512
rect 118 468 122 472
rect 182 488 186 492
rect 254 638 258 642
rect 270 628 274 632
rect 286 588 290 592
rect 510 1128 514 1132
rect 526 1088 530 1092
rect 486 1078 490 1082
rect 542 1058 546 1062
rect 398 968 402 972
rect 390 948 394 952
rect 398 928 402 932
rect 438 978 442 982
rect 414 958 418 962
rect 470 958 474 962
rect 574 1228 578 1232
rect 566 1158 570 1162
rect 606 1158 610 1162
rect 654 1398 658 1402
rect 750 1498 754 1502
rect 734 1468 738 1472
rect 774 1478 778 1482
rect 790 1468 794 1472
rect 790 1458 794 1462
rect 758 1378 762 1382
rect 766 1358 770 1362
rect 670 1348 674 1352
rect 702 1348 706 1352
rect 758 1348 762 1352
rect 718 1338 722 1342
rect 782 1418 786 1422
rect 790 1378 794 1382
rect 782 1348 786 1352
rect 774 1318 778 1322
rect 750 1298 754 1302
rect 734 1288 738 1292
rect 702 1278 706 1282
rect 774 1278 778 1282
rect 750 1268 754 1272
rect 830 1728 834 1732
rect 850 1703 854 1707
rect 857 1703 861 1707
rect 918 1718 922 1722
rect 926 1718 930 1722
rect 894 1688 898 1692
rect 870 1678 874 1682
rect 950 1678 954 1682
rect 910 1668 914 1672
rect 926 1668 930 1672
rect 942 1668 946 1672
rect 846 1648 850 1652
rect 878 1638 882 1642
rect 814 1628 818 1632
rect 838 1628 842 1632
rect 814 1548 818 1552
rect 878 1528 882 1532
rect 814 1498 818 1502
rect 806 1418 810 1422
rect 830 1488 834 1492
rect 850 1503 854 1507
rect 857 1503 861 1507
rect 846 1488 850 1492
rect 814 1358 818 1362
rect 910 1548 914 1552
rect 918 1528 922 1532
rect 958 1608 962 1612
rect 894 1478 898 1482
rect 870 1468 874 1472
rect 918 1468 922 1472
rect 846 1458 850 1462
rect 838 1438 842 1442
rect 886 1438 890 1442
rect 838 1418 842 1422
rect 870 1338 874 1342
rect 798 1288 802 1292
rect 806 1288 810 1292
rect 846 1328 850 1332
rect 1078 1768 1082 1772
rect 1110 1898 1114 1902
rect 1102 1878 1106 1882
rect 1094 1868 1098 1872
rect 1134 1928 1138 1932
rect 1126 1918 1130 1922
rect 1134 1908 1138 1912
rect 1182 2058 1186 2062
rect 1214 2058 1218 2062
rect 1190 2038 1194 2042
rect 1182 2028 1186 2032
rect 1270 2128 1274 2132
rect 1270 2118 1274 2122
rect 1246 2078 1250 2082
rect 1254 2078 1258 2082
rect 1238 2068 1242 2072
rect 1246 2068 1250 2072
rect 1318 2248 1322 2252
rect 1342 2238 1346 2242
rect 1406 2298 1410 2302
rect 1406 2278 1410 2282
rect 1318 2178 1322 2182
rect 1310 2108 1314 2112
rect 1374 2208 1378 2212
rect 1354 2203 1358 2207
rect 1361 2203 1365 2207
rect 1430 2338 1434 2342
rect 1446 2338 1450 2342
rect 1518 2488 1522 2492
rect 1510 2468 1514 2472
rect 1550 2528 1554 2532
rect 1590 2528 1594 2532
rect 1590 2518 1594 2522
rect 1558 2508 1562 2512
rect 1534 2468 1538 2472
rect 1510 2448 1514 2452
rect 1502 2408 1506 2412
rect 1518 2398 1522 2402
rect 1502 2348 1506 2352
rect 1550 2458 1554 2462
rect 1574 2458 1578 2462
rect 1534 2398 1538 2402
rect 1526 2358 1530 2362
rect 1558 2368 1562 2372
rect 1630 2538 1634 2542
rect 1662 2538 1666 2542
rect 1630 2518 1634 2522
rect 1598 2498 1602 2502
rect 1606 2468 1610 2472
rect 1614 2468 1618 2472
rect 1694 2558 1698 2562
rect 1678 2508 1682 2512
rect 1646 2488 1650 2492
rect 1638 2458 1642 2462
rect 1646 2438 1650 2442
rect 1686 2448 1690 2452
rect 1798 2898 1802 2902
rect 1822 2898 1826 2902
rect 1782 2868 1786 2872
rect 1798 2868 1802 2872
rect 1774 2858 1778 2862
rect 1782 2848 1786 2852
rect 1830 2848 1834 2852
rect 1806 2818 1810 2822
rect 1742 2798 1746 2802
rect 1758 2798 1762 2802
rect 1734 2778 1738 2782
rect 1758 2788 1762 2792
rect 1822 2808 1826 2812
rect 1814 2798 1818 2802
rect 1734 2738 1738 2742
rect 1766 2738 1770 2742
rect 1750 2728 1754 2732
rect 1758 2728 1762 2732
rect 1774 2718 1778 2722
rect 1734 2698 1738 2702
rect 1806 2738 1810 2742
rect 1870 3058 1874 3062
rect 1878 3058 1882 3062
rect 1854 3048 1858 3052
rect 1886 3048 1890 3052
rect 1902 3048 1906 3052
rect 1886 3028 1890 3032
rect 1910 2978 1914 2982
rect 1874 2903 1878 2907
rect 1881 2903 1885 2907
rect 1942 2928 1946 2932
rect 1910 2898 1914 2902
rect 1862 2888 1866 2892
rect 1894 2868 1898 2872
rect 1838 2788 1842 2792
rect 1934 2808 1938 2812
rect 1830 2738 1834 2742
rect 1838 2738 1842 2742
rect 1886 2738 1890 2742
rect 1782 2688 1786 2692
rect 1750 2678 1754 2682
rect 1758 2658 1762 2662
rect 1782 2658 1786 2662
rect 1790 2658 1794 2662
rect 1718 2538 1722 2542
rect 1686 2438 1690 2442
rect 1710 2438 1714 2442
rect 1630 2388 1634 2392
rect 1614 2368 1618 2372
rect 1598 2358 1602 2362
rect 1494 2338 1498 2342
rect 1582 2338 1586 2342
rect 1462 2328 1466 2332
rect 1454 2298 1458 2302
rect 1430 2258 1434 2262
rect 1438 2258 1442 2262
rect 1430 2218 1434 2222
rect 1422 2198 1426 2202
rect 1406 2158 1410 2162
rect 1478 2288 1482 2292
rect 1534 2328 1538 2332
rect 1566 2328 1570 2332
rect 1502 2308 1506 2312
rect 1630 2348 1634 2352
rect 1622 2338 1626 2342
rect 1638 2338 1642 2342
rect 1606 2328 1610 2332
rect 1598 2318 1602 2322
rect 1614 2318 1618 2322
rect 1614 2308 1618 2312
rect 1566 2288 1570 2292
rect 1518 2268 1522 2272
rect 1534 2268 1538 2272
rect 1558 2268 1562 2272
rect 1462 2258 1466 2262
rect 1478 2258 1482 2262
rect 1478 2218 1482 2222
rect 1526 2258 1530 2262
rect 1558 2238 1562 2242
rect 1542 2218 1546 2222
rect 1566 2218 1570 2222
rect 1502 2208 1506 2212
rect 1710 2398 1714 2402
rect 1758 2628 1762 2632
rect 1766 2628 1770 2632
rect 1750 2598 1754 2602
rect 1862 2728 1866 2732
rect 1902 2718 1906 2722
rect 1874 2703 1878 2707
rect 1881 2703 1885 2707
rect 1998 3068 2002 3072
rect 1958 3018 1962 3022
rect 1990 3018 1994 3022
rect 1966 2978 1970 2982
rect 2006 2958 2010 2962
rect 2022 3098 2026 3102
rect 2038 3108 2042 3112
rect 1966 2948 1970 2952
rect 1998 2948 2002 2952
rect 2014 2948 2018 2952
rect 2094 3148 2098 3152
rect 2086 3138 2090 3142
rect 2134 3278 2138 3282
rect 2286 3738 2290 3742
rect 2318 3738 2322 3742
rect 2374 3848 2378 3852
rect 2446 3868 2450 3872
rect 2438 3828 2442 3832
rect 2386 3803 2390 3807
rect 2393 3803 2397 3807
rect 2366 3798 2370 3802
rect 2358 3768 2362 3772
rect 2390 3778 2394 3782
rect 2358 3738 2362 3742
rect 2278 3728 2282 3732
rect 2310 3728 2314 3732
rect 2326 3728 2330 3732
rect 2342 3728 2346 3732
rect 2334 3718 2338 3722
rect 2286 3688 2290 3692
rect 2294 3658 2298 3662
rect 2326 3658 2330 3662
rect 2270 3628 2274 3632
rect 2230 3598 2234 3602
rect 2326 3588 2330 3592
rect 2238 3568 2242 3572
rect 2206 3548 2210 3552
rect 2222 3548 2226 3552
rect 2254 3558 2258 3562
rect 2278 3558 2282 3562
rect 2326 3558 2330 3562
rect 2254 3548 2258 3552
rect 2270 3548 2274 3552
rect 2190 3518 2194 3522
rect 2310 3548 2314 3552
rect 2278 3508 2282 3512
rect 2358 3608 2362 3612
rect 2342 3598 2346 3602
rect 2350 3558 2354 3562
rect 2358 3548 2362 3552
rect 2326 3528 2330 3532
rect 2302 3518 2306 3522
rect 2334 3508 2338 3512
rect 2214 3498 2218 3502
rect 2294 3498 2298 3502
rect 2358 3528 2362 3532
rect 2374 3698 2378 3702
rect 2502 3938 2506 3942
rect 2566 4378 2570 4382
rect 2590 4408 2594 4412
rect 2566 4368 2570 4372
rect 2582 4368 2586 4372
rect 2550 4308 2554 4312
rect 2558 4288 2562 4292
rect 2566 4278 2570 4282
rect 2574 4258 2578 4262
rect 2534 4248 2538 4252
rect 2606 4358 2610 4362
rect 2590 4228 2594 4232
rect 2582 4208 2586 4212
rect 2550 4188 2554 4192
rect 2526 4178 2530 4182
rect 2598 4168 2602 4172
rect 2558 4148 2562 4152
rect 2622 4148 2626 4152
rect 2702 4598 2706 4602
rect 2742 4588 2746 4592
rect 2758 4568 2762 4572
rect 2766 4558 2770 4562
rect 2782 4558 2786 4562
rect 2798 4558 2802 4562
rect 2782 4548 2786 4552
rect 2846 4648 2850 4652
rect 2846 4628 2850 4632
rect 2838 4548 2842 4552
rect 2798 4538 2802 4542
rect 2814 4538 2818 4542
rect 2742 4518 2746 4522
rect 2726 4488 2730 4492
rect 2702 4468 2706 4472
rect 2710 4468 2714 4472
rect 2742 4478 2746 4482
rect 2694 4438 2698 4442
rect 2662 4428 2666 4432
rect 2670 4378 2674 4382
rect 2790 4508 2794 4512
rect 2830 4498 2834 4502
rect 2814 4488 2818 4492
rect 2822 4488 2826 4492
rect 2846 4488 2850 4492
rect 2758 4448 2762 4452
rect 2718 4418 2722 4422
rect 2734 4418 2738 4422
rect 2766 4418 2770 4422
rect 2710 4388 2714 4392
rect 2718 4378 2722 4382
rect 2662 4368 2666 4372
rect 2638 4358 2642 4362
rect 2686 4368 2690 4372
rect 2694 4358 2698 4362
rect 2758 4388 2762 4392
rect 2838 4468 2842 4472
rect 2870 4558 2874 4562
rect 2950 4608 2954 4612
rect 2950 4548 2954 4552
rect 2998 4658 3002 4662
rect 3014 4628 3018 4632
rect 3054 4758 3058 4762
rect 3062 4748 3066 4752
rect 3070 4738 3074 4742
rect 3070 4658 3074 4662
rect 3054 4648 3058 4652
rect 3046 4628 3050 4632
rect 3030 4568 3034 4572
rect 3046 4558 3050 4562
rect 3030 4548 3034 4552
rect 2982 4538 2986 4542
rect 2870 4528 2874 4532
rect 2910 4528 2914 4532
rect 3006 4528 3010 4532
rect 2890 4503 2894 4507
rect 2897 4503 2901 4507
rect 2894 4488 2898 4492
rect 3030 4508 3034 4512
rect 3006 4488 3010 4492
rect 2910 4478 2914 4482
rect 2854 4468 2858 4472
rect 2878 4468 2882 4472
rect 2974 4468 2978 4472
rect 3022 4468 3026 4472
rect 2830 4458 2834 4462
rect 2814 4438 2818 4442
rect 2806 4428 2810 4432
rect 2774 4368 2778 4372
rect 2798 4368 2802 4372
rect 2734 4348 2738 4352
rect 2750 4348 2754 4352
rect 2766 4348 2770 4352
rect 2798 4348 2802 4352
rect 2694 4308 2698 4312
rect 2678 4288 2682 4292
rect 2662 4218 2666 4222
rect 2710 4338 2714 4342
rect 2718 4338 2722 4342
rect 2758 4338 2762 4342
rect 2734 4318 2738 4322
rect 2774 4318 2778 4322
rect 2726 4308 2730 4312
rect 2710 4248 2714 4252
rect 2702 4208 2706 4212
rect 2646 4148 2650 4152
rect 2614 4138 2618 4142
rect 2558 4128 2562 4132
rect 2694 4138 2698 4142
rect 2566 4118 2570 4122
rect 2630 4118 2634 4122
rect 2638 4118 2642 4122
rect 2678 4118 2682 4122
rect 2534 4108 2538 4112
rect 2526 4098 2530 4102
rect 2550 4098 2554 4102
rect 2534 3968 2538 3972
rect 2558 4068 2562 4072
rect 2622 4098 2626 4102
rect 2598 4078 2602 4082
rect 2686 4098 2690 4102
rect 2630 4088 2634 4092
rect 2718 4168 2722 4172
rect 2774 4288 2778 4292
rect 2774 4278 2778 4282
rect 2870 4458 2874 4462
rect 2870 4378 2874 4382
rect 2830 4348 2834 4352
rect 2854 4338 2858 4342
rect 2798 4328 2802 4332
rect 2822 4328 2826 4332
rect 2830 4318 2834 4322
rect 2806 4278 2810 4282
rect 2838 4278 2842 4282
rect 2798 4268 2802 4272
rect 2814 4268 2818 4272
rect 2782 4238 2786 4242
rect 2814 4238 2818 4242
rect 2774 4228 2778 4232
rect 2798 4228 2802 4232
rect 2750 4198 2754 4202
rect 2774 4178 2778 4182
rect 2758 4168 2762 4172
rect 2742 4158 2746 4162
rect 2782 4158 2786 4162
rect 2598 4068 2602 4072
rect 2694 4068 2698 4072
rect 2702 4068 2706 4072
rect 2590 4058 2594 4062
rect 2574 4048 2578 4052
rect 2582 3978 2586 3982
rect 2534 3938 2538 3942
rect 2518 3928 2522 3932
rect 2486 3878 2490 3882
rect 2622 3958 2626 3962
rect 2582 3938 2586 3942
rect 2558 3918 2562 3922
rect 2566 3918 2570 3922
rect 2566 3908 2570 3912
rect 2590 3908 2594 3912
rect 2574 3898 2578 3902
rect 2510 3888 2514 3892
rect 2550 3878 2554 3882
rect 2502 3868 2506 3872
rect 2574 3868 2578 3872
rect 2486 3838 2490 3842
rect 2574 3848 2578 3852
rect 2566 3838 2570 3842
rect 2502 3808 2506 3812
rect 2502 3798 2506 3802
rect 2478 3758 2482 3762
rect 2502 3748 2506 3752
rect 2414 3728 2418 3732
rect 2422 3728 2426 3732
rect 2398 3688 2402 3692
rect 2446 3738 2450 3742
rect 2502 3738 2506 3742
rect 2558 3738 2562 3742
rect 2486 3728 2490 3732
rect 2494 3708 2498 3712
rect 2462 3698 2466 3702
rect 2430 3678 2434 3682
rect 2414 3668 2418 3672
rect 2386 3603 2390 3607
rect 2393 3603 2397 3607
rect 2374 3518 2378 3522
rect 2342 3488 2346 3492
rect 2366 3488 2370 3492
rect 2398 3488 2402 3492
rect 2198 3478 2202 3482
rect 2326 3478 2330 3482
rect 2446 3658 2450 3662
rect 2422 3648 2426 3652
rect 2438 3648 2442 3652
rect 2438 3628 2442 3632
rect 2422 3608 2426 3612
rect 2486 3658 2490 3662
rect 2494 3648 2498 3652
rect 2454 3588 2458 3592
rect 2478 3578 2482 3582
rect 2446 3518 2450 3522
rect 2350 3478 2354 3482
rect 2414 3478 2418 3482
rect 2206 3468 2210 3472
rect 2214 3468 2218 3472
rect 2342 3468 2346 3472
rect 2198 3438 2202 3442
rect 2286 3438 2290 3442
rect 2246 3418 2250 3422
rect 2310 3418 2314 3422
rect 2350 3448 2354 3452
rect 2374 3438 2378 3442
rect 2366 3408 2370 3412
rect 2326 3398 2330 3402
rect 2302 3378 2306 3382
rect 2254 3347 2258 3351
rect 2198 3338 2202 3342
rect 2182 3328 2186 3332
rect 2190 3318 2194 3322
rect 2206 3318 2210 3322
rect 2174 3308 2178 3312
rect 2166 3298 2170 3302
rect 2142 3168 2146 3172
rect 2182 3238 2186 3242
rect 2150 3148 2154 3152
rect 2086 3128 2090 3132
rect 2118 3128 2122 3132
rect 2070 3108 2074 3112
rect 2054 3088 2058 3092
rect 2062 3088 2066 3092
rect 2046 3068 2050 3072
rect 2054 3058 2058 3062
rect 2070 3058 2074 3062
rect 2078 3058 2082 3062
rect 2062 3048 2066 3052
rect 2070 2998 2074 3002
rect 2054 2968 2058 2972
rect 2078 2988 2082 2992
rect 2070 2938 2074 2942
rect 2134 3108 2138 3112
rect 2094 3078 2098 3082
rect 2126 3068 2130 3072
rect 2182 3088 2186 3092
rect 2150 3068 2154 3072
rect 2110 3058 2114 3062
rect 2134 3038 2138 3042
rect 2166 3038 2170 3042
rect 2110 3028 2114 3032
rect 2094 3018 2098 3022
rect 2126 3018 2130 3022
rect 2102 2948 2106 2952
rect 2070 2928 2074 2932
rect 2078 2928 2082 2932
rect 2086 2928 2090 2932
rect 1982 2918 1986 2922
rect 2022 2918 2026 2922
rect 1998 2898 2002 2902
rect 1974 2868 1978 2872
rect 2038 2888 2042 2892
rect 2038 2878 2042 2882
rect 2070 2868 2074 2872
rect 2094 2918 2098 2922
rect 2110 2918 2114 2922
rect 2086 2888 2090 2892
rect 2102 2888 2106 2892
rect 2054 2848 2058 2852
rect 2070 2848 2074 2852
rect 2078 2848 2082 2852
rect 1974 2838 1978 2842
rect 2006 2778 2010 2782
rect 1950 2748 1954 2752
rect 2038 2768 2042 2772
rect 1942 2728 1946 2732
rect 1998 2718 2002 2722
rect 1934 2688 1938 2692
rect 1998 2678 2002 2682
rect 1830 2668 1834 2672
rect 1862 2668 1866 2672
rect 1870 2668 1874 2672
rect 1838 2658 1842 2662
rect 1822 2648 1826 2652
rect 1822 2628 1826 2632
rect 1806 2608 1810 2612
rect 2038 2738 2042 2742
rect 2030 2708 2034 2712
rect 2046 2698 2050 2702
rect 2070 2838 2074 2842
rect 2062 2828 2066 2832
rect 2094 2808 2098 2812
rect 2118 2908 2122 2912
rect 2110 2848 2114 2852
rect 2118 2828 2122 2832
rect 2094 2798 2098 2802
rect 2102 2798 2106 2802
rect 2150 2888 2154 2892
rect 2142 2878 2146 2882
rect 2182 2998 2186 3002
rect 2174 2938 2178 2942
rect 2174 2898 2178 2902
rect 2174 2888 2178 2892
rect 2182 2878 2186 2882
rect 2142 2858 2146 2862
rect 2294 3318 2298 3322
rect 2262 3308 2266 3312
rect 2246 3298 2250 3302
rect 2198 3288 2202 3292
rect 2238 3288 2242 3292
rect 2254 3288 2258 3292
rect 2214 3278 2218 3282
rect 2270 3288 2274 3292
rect 2294 3288 2298 3292
rect 2246 3248 2250 3252
rect 2230 3228 2234 3232
rect 2230 3168 2234 3172
rect 2222 3148 2226 3152
rect 2198 3008 2202 3012
rect 2286 3238 2290 3242
rect 2318 3348 2322 3352
rect 2310 3338 2314 3342
rect 2326 3338 2330 3342
rect 2302 3238 2306 3242
rect 2294 3218 2298 3222
rect 2302 3168 2306 3172
rect 2342 3308 2346 3312
rect 2358 3258 2362 3262
rect 2438 3418 2442 3422
rect 2386 3403 2390 3407
rect 2393 3403 2397 3407
rect 2422 3398 2426 3402
rect 2398 3328 2402 3332
rect 2382 3288 2386 3292
rect 2462 3488 2466 3492
rect 2518 3708 2522 3712
rect 2542 3698 2546 3702
rect 2550 3698 2554 3702
rect 2526 3678 2530 3682
rect 2582 3808 2586 3812
rect 2646 3968 2650 3972
rect 2638 3928 2642 3932
rect 2638 3908 2642 3912
rect 2622 3888 2626 3892
rect 2598 3858 2602 3862
rect 2582 3738 2586 3742
rect 2566 3698 2570 3702
rect 2582 3698 2586 3702
rect 2558 3678 2562 3682
rect 2694 4048 2698 4052
rect 2726 4128 2730 4132
rect 2734 4118 2738 4122
rect 2790 4138 2794 4142
rect 2766 4118 2770 4122
rect 2718 4058 2722 4062
rect 2710 3958 2714 3962
rect 2694 3948 2698 3952
rect 2702 3928 2706 3932
rect 2662 3888 2666 3892
rect 2646 3868 2650 3872
rect 2662 3868 2666 3872
rect 2678 3868 2682 3872
rect 2670 3858 2674 3862
rect 2630 3838 2634 3842
rect 2630 3758 2634 3762
rect 2622 3748 2626 3752
rect 2606 3698 2610 3702
rect 2598 3668 2602 3672
rect 2534 3648 2538 3652
rect 2526 3638 2530 3642
rect 2534 3598 2538 3602
rect 2510 3588 2514 3592
rect 2574 3648 2578 3652
rect 2542 3568 2546 3572
rect 2550 3558 2554 3562
rect 2510 3548 2514 3552
rect 2646 3838 2650 3842
rect 2710 3838 2714 3842
rect 2734 4008 2738 4012
rect 2750 3968 2754 3972
rect 2726 3908 2730 3912
rect 2742 3908 2746 3912
rect 2742 3878 2746 3882
rect 2734 3868 2738 3872
rect 2718 3818 2722 3822
rect 2702 3768 2706 3772
rect 2670 3758 2674 3762
rect 2694 3758 2698 3762
rect 2982 4378 2986 4382
rect 2894 4348 2898 4352
rect 2870 4328 2874 4332
rect 2934 4318 2938 4322
rect 2890 4303 2894 4307
rect 2897 4303 2901 4307
rect 2878 4278 2882 4282
rect 2918 4278 2922 4282
rect 2910 4238 2914 4242
rect 2926 4238 2930 4242
rect 2934 4238 2938 4242
rect 2870 4228 2874 4232
rect 2862 4208 2866 4212
rect 2854 4198 2858 4202
rect 2814 4168 2818 4172
rect 2814 4158 2818 4162
rect 2814 4148 2818 4152
rect 2934 4218 2938 4222
rect 2878 4158 2882 4162
rect 3014 4358 3018 4362
rect 3446 5058 3450 5062
rect 3542 5058 3546 5062
rect 3574 5058 3578 5062
rect 3670 5058 3674 5062
rect 3950 5058 3954 5062
rect 3214 5048 3218 5052
rect 3342 5048 3346 5052
rect 3262 5038 3266 5042
rect 3430 5038 3434 5042
rect 3214 5008 3218 5012
rect 3206 4998 3210 5002
rect 3198 4948 3202 4952
rect 3206 4938 3210 4942
rect 3230 4978 3234 4982
rect 3254 4968 3258 4972
rect 3470 5008 3474 5012
rect 3494 5008 3498 5012
rect 3402 5003 3406 5007
rect 3409 5003 3413 5007
rect 3310 4988 3314 4992
rect 3294 4968 3298 4972
rect 3302 4958 3306 4962
rect 3278 4948 3282 4952
rect 3286 4948 3290 4952
rect 3246 4938 3250 4942
rect 3262 4938 3266 4942
rect 3166 4868 3170 4872
rect 3214 4868 3218 4872
rect 3150 4778 3154 4782
rect 3094 4758 3098 4762
rect 3150 4718 3154 4722
rect 3102 4698 3106 4702
rect 3206 4708 3210 4712
rect 3094 4688 3098 4692
rect 3110 4688 3114 4692
rect 3150 4688 3154 4692
rect 3158 4688 3162 4692
rect 3086 4648 3090 4652
rect 3078 4638 3082 4642
rect 3062 4558 3066 4562
rect 3118 4668 3122 4672
rect 3150 4668 3154 4672
rect 3110 4638 3114 4642
rect 3166 4658 3170 4662
rect 3190 4658 3194 4662
rect 3150 4538 3154 4542
rect 3134 4528 3138 4532
rect 3102 4508 3106 4512
rect 3110 4478 3114 4482
rect 3118 4478 3122 4482
rect 3078 4468 3082 4472
rect 3102 4468 3106 4472
rect 3110 4468 3114 4472
rect 3198 4648 3202 4652
rect 3230 4878 3234 4882
rect 3278 4928 3282 4932
rect 3350 4978 3354 4982
rect 3462 4978 3466 4982
rect 3334 4958 3338 4962
rect 3254 4868 3258 4872
rect 3286 4868 3290 4872
rect 3302 4868 3306 4872
rect 3246 4858 3250 4862
rect 3278 4858 3282 4862
rect 3238 4718 3242 4722
rect 3230 4678 3234 4682
rect 3262 4848 3266 4852
rect 3262 4838 3266 4842
rect 3254 4668 3258 4672
rect 3270 4828 3274 4832
rect 3310 4828 3314 4832
rect 3302 4788 3306 4792
rect 3286 4748 3290 4752
rect 3270 4728 3274 4732
rect 3310 4747 3314 4751
rect 3302 4688 3306 4692
rect 3438 4968 3442 4972
rect 3366 4948 3370 4952
rect 3382 4938 3386 4942
rect 3414 4898 3418 4902
rect 3438 4888 3442 4892
rect 3398 4858 3402 4862
rect 3350 4848 3354 4852
rect 3326 4828 3330 4832
rect 3402 4803 3406 4807
rect 3409 4803 3413 4807
rect 3430 4778 3434 4782
rect 3382 4768 3386 4772
rect 3414 4758 3418 4762
rect 3374 4748 3378 4752
rect 3350 4718 3354 4722
rect 3358 4718 3362 4722
rect 3398 4688 3402 4692
rect 3366 4678 3370 4682
rect 3270 4668 3274 4672
rect 3318 4668 3322 4672
rect 3350 4668 3354 4672
rect 3382 4668 3386 4672
rect 3422 4678 3426 4682
rect 3246 4658 3250 4662
rect 3254 4608 3258 4612
rect 3326 4648 3330 4652
rect 3382 4648 3386 4652
rect 3358 4638 3362 4642
rect 3406 4638 3410 4642
rect 3342 4618 3346 4622
rect 3262 4578 3266 4582
rect 3222 4558 3226 4562
rect 3294 4558 3298 4562
rect 3326 4558 3330 4562
rect 3358 4558 3362 4562
rect 3198 4548 3202 4552
rect 3182 4538 3186 4542
rect 3214 4508 3218 4512
rect 3230 4528 3234 4532
rect 3166 4498 3170 4502
rect 3222 4498 3226 4502
rect 3262 4518 3266 4522
rect 3270 4498 3274 4502
rect 3158 4478 3162 4482
rect 3246 4478 3250 4482
rect 3150 4468 3154 4472
rect 3174 4468 3178 4472
rect 3222 4468 3226 4472
rect 3070 4458 3074 4462
rect 3118 4458 3122 4462
rect 3054 4448 3058 4452
rect 3078 4448 3082 4452
rect 3046 4398 3050 4402
rect 3086 4398 3090 4402
rect 3070 4358 3074 4362
rect 3054 4328 3058 4332
rect 3038 4318 3042 4322
rect 2990 4308 2994 4312
rect 2982 4288 2986 4292
rect 2982 4278 2986 4282
rect 2950 4248 2954 4252
rect 3038 4288 3042 4292
rect 3014 4278 3018 4282
rect 3006 4268 3010 4272
rect 3014 4248 3018 4252
rect 3070 4268 3074 4272
rect 3030 4248 3034 4252
rect 2982 4208 2986 4212
rect 3022 4208 3026 4212
rect 3046 4188 3050 4192
rect 3022 4168 3026 4172
rect 3198 4458 3202 4462
rect 3230 4458 3234 4462
rect 3206 4448 3210 4452
rect 3134 4398 3138 4402
rect 3222 4438 3226 4442
rect 3254 4448 3258 4452
rect 3342 4548 3346 4552
rect 3318 4538 3322 4542
rect 3326 4528 3330 4532
rect 3374 4518 3378 4522
rect 3334 4488 3338 4492
rect 3382 4478 3386 4482
rect 3310 4468 3314 4472
rect 3350 4448 3354 4452
rect 3358 4448 3362 4452
rect 3286 4438 3290 4442
rect 3366 4438 3370 4442
rect 3190 4428 3194 4432
rect 3238 4428 3242 4432
rect 3150 4388 3154 4392
rect 3126 4378 3130 4382
rect 3102 4338 3106 4342
rect 3134 4338 3138 4342
rect 3118 4318 3122 4322
rect 3094 4218 3098 4222
rect 3046 4158 3050 4162
rect 3110 4158 3114 4162
rect 3126 4288 3130 4292
rect 3174 4288 3178 4292
rect 3166 4278 3170 4282
rect 3182 4268 3186 4272
rect 3150 4248 3154 4252
rect 3166 4238 3170 4242
rect 3182 4178 3186 4182
rect 3150 4158 3154 4162
rect 3134 4148 3138 4152
rect 3022 4138 3026 4142
rect 3086 4138 3090 4142
rect 3102 4138 3106 4142
rect 2870 4128 2874 4132
rect 2798 4108 2802 4112
rect 2814 4108 2818 4112
rect 2774 4098 2778 4102
rect 2830 4088 2834 4092
rect 2798 4078 2802 4082
rect 2782 4068 2786 4072
rect 2766 4048 2770 4052
rect 2830 4058 2834 4062
rect 2822 4038 2826 4042
rect 2830 4028 2834 4032
rect 2774 4018 2778 4022
rect 2890 4103 2894 4107
rect 2897 4103 2901 4107
rect 2918 4088 2922 4092
rect 2934 4088 2938 4092
rect 2926 4078 2930 4082
rect 2894 4068 2898 4072
rect 2950 4058 2954 4062
rect 2966 4058 2970 4062
rect 2862 4048 2866 4052
rect 2870 4048 2874 4052
rect 2894 4048 2898 4052
rect 2862 4028 2866 4032
rect 2846 3968 2850 3972
rect 2766 3958 2770 3962
rect 2830 3958 2834 3962
rect 2942 3978 2946 3982
rect 2782 3948 2786 3952
rect 2806 3948 2810 3952
rect 2838 3948 2842 3952
rect 2854 3948 2858 3952
rect 2766 3788 2770 3792
rect 2798 3938 2802 3942
rect 2918 3948 2922 3952
rect 3078 4128 3082 4132
rect 3022 4108 3026 4112
rect 3150 4138 3154 4142
rect 3326 4347 3330 4351
rect 3350 4348 3354 4352
rect 3198 4268 3202 4272
rect 3302 4338 3306 4342
rect 3254 4328 3258 4332
rect 3238 4318 3242 4322
rect 3254 4318 3258 4322
rect 3278 4318 3282 4322
rect 3286 4318 3290 4322
rect 3222 4288 3226 4292
rect 3270 4268 3274 4272
rect 3230 4258 3234 4262
rect 3262 4258 3266 4262
rect 3246 4248 3250 4252
rect 3278 4218 3282 4222
rect 3382 4458 3386 4462
rect 3402 4603 3406 4607
rect 3409 4603 3413 4607
rect 3414 4568 3418 4572
rect 3422 4548 3426 4552
rect 3406 4528 3410 4532
rect 3398 4508 3402 4512
rect 3414 4468 3418 4472
rect 3390 4448 3394 4452
rect 3390 4438 3394 4442
rect 3382 4378 3386 4382
rect 3398 4428 3402 4432
rect 3402 4403 3406 4407
rect 3409 4403 3413 4407
rect 3414 4368 3418 4372
rect 3374 4348 3378 4352
rect 3390 4348 3394 4352
rect 3398 4348 3402 4352
rect 3374 4338 3378 4342
rect 3366 4318 3370 4322
rect 3318 4258 3322 4262
rect 3286 4198 3290 4202
rect 3238 4138 3242 4142
rect 3246 4138 3250 4142
rect 3190 4118 3194 4122
rect 2998 4088 3002 4092
rect 3118 4088 3122 4092
rect 3006 4078 3010 4082
rect 3118 4078 3122 4082
rect 3206 4108 3210 4112
rect 3198 4098 3202 4102
rect 3022 4068 3026 4072
rect 3046 4068 3050 4072
rect 3094 4068 3098 4072
rect 3190 4068 3194 4072
rect 3006 4058 3010 4062
rect 3070 4058 3074 4062
rect 3102 4058 3106 4062
rect 3022 4048 3026 4052
rect 2990 4018 2994 4022
rect 3038 4008 3042 4012
rect 3006 3978 3010 3982
rect 3134 4038 3138 4042
rect 3150 4038 3154 4042
rect 3094 4028 3098 4032
rect 3118 4018 3122 4022
rect 3102 3978 3106 3982
rect 3142 3978 3146 3982
rect 3070 3948 3074 3952
rect 3086 3948 3090 3952
rect 3126 3948 3130 3952
rect 3150 3958 3154 3962
rect 3182 3958 3186 3962
rect 3222 4078 3226 4082
rect 3230 4078 3234 4082
rect 3214 4058 3218 4062
rect 3222 3988 3226 3992
rect 3214 3978 3218 3982
rect 3158 3948 3162 3952
rect 2878 3938 2882 3942
rect 3046 3938 3050 3942
rect 3110 3938 3114 3942
rect 3134 3938 3138 3942
rect 2870 3928 2874 3932
rect 2822 3888 2826 3892
rect 2838 3878 2842 3882
rect 2846 3878 2850 3882
rect 2838 3858 2842 3862
rect 2846 3858 2850 3862
rect 2806 3848 2810 3852
rect 2806 3768 2810 3772
rect 2822 3768 2826 3772
rect 2662 3748 2666 3752
rect 2694 3748 2698 3752
rect 2726 3748 2730 3752
rect 2742 3748 2746 3752
rect 2782 3748 2786 3752
rect 2638 3738 2642 3742
rect 2686 3738 2690 3742
rect 2702 3738 2706 3742
rect 2662 3728 2666 3732
rect 2654 3698 2658 3702
rect 2694 3708 2698 3712
rect 2718 3708 2722 3712
rect 2630 3688 2634 3692
rect 2646 3688 2650 3692
rect 2630 3658 2634 3662
rect 2590 3628 2594 3632
rect 2574 3588 2578 3592
rect 2654 3648 2658 3652
rect 2638 3638 2642 3642
rect 2606 3628 2610 3632
rect 2582 3578 2586 3582
rect 2598 3578 2602 3582
rect 2574 3558 2578 3562
rect 2614 3618 2618 3622
rect 2598 3558 2602 3562
rect 2590 3548 2594 3552
rect 2534 3518 2538 3522
rect 2662 3628 2666 3632
rect 2710 3658 2714 3662
rect 2702 3638 2706 3642
rect 2710 3628 2714 3632
rect 2718 3628 2722 3632
rect 2686 3598 2690 3602
rect 2638 3568 2642 3572
rect 2646 3558 2650 3562
rect 2686 3558 2690 3562
rect 2646 3548 2650 3552
rect 2518 3488 2522 3492
rect 2510 3458 2514 3462
rect 2566 3458 2570 3462
rect 2502 3438 2506 3442
rect 2550 3448 2554 3452
rect 2510 3408 2514 3412
rect 2446 3398 2450 3402
rect 2470 3348 2474 3352
rect 2470 3338 2474 3342
rect 2478 3338 2482 3342
rect 2486 3338 2490 3342
rect 2462 3308 2466 3312
rect 2438 3298 2442 3302
rect 2390 3278 2394 3282
rect 2438 3278 2442 3282
rect 2374 3218 2378 3222
rect 2386 3203 2390 3207
rect 2393 3203 2397 3207
rect 2278 3148 2282 3152
rect 2310 3148 2314 3152
rect 2262 3138 2266 3142
rect 2262 3058 2266 3062
rect 2326 3138 2330 3142
rect 2502 3328 2506 3332
rect 2510 3298 2514 3302
rect 2494 3288 2498 3292
rect 2582 3418 2586 3422
rect 2550 3338 2554 3342
rect 2470 3258 2474 3262
rect 2502 3258 2506 3262
rect 2518 3258 2522 3262
rect 2414 3238 2418 3242
rect 2358 3138 2362 3142
rect 2294 3118 2298 3122
rect 2326 3118 2330 3122
rect 2286 3098 2290 3102
rect 2294 3078 2298 3082
rect 2342 3078 2346 3082
rect 2310 3068 2314 3072
rect 2278 3048 2282 3052
rect 2270 3038 2274 3042
rect 2302 3038 2306 3042
rect 2270 2998 2274 3002
rect 2238 2988 2242 2992
rect 2246 2988 2250 2992
rect 2246 2978 2250 2982
rect 2350 3008 2354 3012
rect 2334 2988 2338 2992
rect 2318 2958 2322 2962
rect 2206 2948 2210 2952
rect 2262 2948 2266 2952
rect 2214 2938 2218 2942
rect 2214 2888 2218 2892
rect 2270 2888 2274 2892
rect 2278 2878 2282 2882
rect 2182 2848 2186 2852
rect 2190 2848 2194 2852
rect 2134 2838 2138 2842
rect 2094 2738 2098 2742
rect 2070 2728 2074 2732
rect 2030 2678 2034 2682
rect 2038 2678 2042 2682
rect 1926 2668 1930 2672
rect 2014 2668 2018 2672
rect 1878 2608 1882 2612
rect 1830 2598 1834 2602
rect 1766 2558 1770 2562
rect 1894 2558 1898 2562
rect 1798 2548 1802 2552
rect 1774 2528 1778 2532
rect 1758 2468 1762 2472
rect 1782 2468 1786 2472
rect 1814 2468 1818 2472
rect 1790 2458 1794 2462
rect 1806 2448 1810 2452
rect 1734 2418 1738 2422
rect 1774 2408 1778 2412
rect 1766 2398 1770 2402
rect 1662 2358 1666 2362
rect 1670 2358 1674 2362
rect 1726 2358 1730 2362
rect 1750 2358 1754 2362
rect 1998 2658 2002 2662
rect 2062 2658 2066 2662
rect 1918 2618 1922 2622
rect 1926 2608 1930 2612
rect 1990 2608 1994 2612
rect 2022 2588 2026 2592
rect 1974 2558 1978 2562
rect 2078 2658 2082 2662
rect 2070 2648 2074 2652
rect 2126 2768 2130 2772
rect 2246 2848 2250 2852
rect 2214 2808 2218 2812
rect 2214 2798 2218 2802
rect 2142 2768 2146 2772
rect 2158 2768 2162 2772
rect 2174 2768 2178 2772
rect 2206 2768 2210 2772
rect 2134 2748 2138 2752
rect 2142 2748 2146 2752
rect 2118 2738 2122 2742
rect 2134 2738 2138 2742
rect 2142 2718 2146 2722
rect 2110 2678 2114 2682
rect 2198 2738 2202 2742
rect 2174 2718 2178 2722
rect 2190 2708 2194 2712
rect 2182 2688 2186 2692
rect 2342 2958 2346 2962
rect 2318 2928 2322 2932
rect 2302 2898 2306 2902
rect 2294 2848 2298 2852
rect 2310 2808 2314 2812
rect 2286 2768 2290 2772
rect 2270 2758 2274 2762
rect 2238 2748 2242 2752
rect 2294 2748 2298 2752
rect 2094 2668 2098 2672
rect 2134 2668 2138 2672
rect 2110 2658 2114 2662
rect 2182 2658 2186 2662
rect 2230 2658 2234 2662
rect 2150 2648 2154 2652
rect 2166 2648 2170 2652
rect 2078 2638 2082 2642
rect 2086 2638 2090 2642
rect 2126 2628 2130 2632
rect 2070 2598 2074 2602
rect 2094 2598 2098 2602
rect 2134 2618 2138 2622
rect 2086 2558 2090 2562
rect 2110 2558 2114 2562
rect 1998 2548 2002 2552
rect 1838 2538 1842 2542
rect 1910 2538 1914 2542
rect 1942 2538 1946 2542
rect 1894 2528 1898 2532
rect 1902 2528 1906 2532
rect 1918 2528 1922 2532
rect 1926 2528 1930 2532
rect 1830 2518 1834 2522
rect 1894 2508 1898 2512
rect 1874 2503 1878 2507
rect 1881 2503 1885 2507
rect 1878 2468 1882 2472
rect 1830 2458 1834 2462
rect 1846 2458 1850 2462
rect 1822 2408 1826 2412
rect 1838 2438 1842 2442
rect 1886 2458 1890 2462
rect 1862 2418 1866 2422
rect 1854 2408 1858 2412
rect 1830 2398 1834 2402
rect 1782 2358 1786 2362
rect 1798 2358 1802 2362
rect 1886 2368 1890 2372
rect 1678 2348 1682 2352
rect 1710 2348 1714 2352
rect 1758 2348 1762 2352
rect 1782 2348 1786 2352
rect 1846 2348 1850 2352
rect 1886 2348 1890 2352
rect 1702 2338 1706 2342
rect 1766 2338 1770 2342
rect 1798 2338 1802 2342
rect 1830 2338 1834 2342
rect 1894 2338 1898 2342
rect 1758 2328 1762 2332
rect 1822 2328 1826 2332
rect 1678 2318 1682 2322
rect 1694 2318 1698 2322
rect 1750 2318 1754 2322
rect 1662 2308 1666 2312
rect 1734 2298 1738 2302
rect 1630 2278 1634 2282
rect 1654 2278 1658 2282
rect 1678 2268 1682 2272
rect 1694 2268 1698 2272
rect 1726 2268 1730 2272
rect 1790 2298 1794 2302
rect 1774 2278 1778 2282
rect 1742 2258 1746 2262
rect 1758 2258 1762 2262
rect 1918 2508 1922 2512
rect 1918 2448 1922 2452
rect 1902 2318 1906 2322
rect 1894 2308 1898 2312
rect 1874 2303 1878 2307
rect 1881 2303 1885 2307
rect 1862 2268 1866 2272
rect 1678 2238 1682 2242
rect 1686 2218 1690 2222
rect 1678 2208 1682 2212
rect 1710 2218 1714 2222
rect 1694 2188 1698 2192
rect 1446 2178 1450 2182
rect 1486 2178 1490 2182
rect 1478 2168 1482 2172
rect 1350 2148 1354 2152
rect 1366 2148 1370 2152
rect 1390 2148 1394 2152
rect 1414 2148 1418 2152
rect 1374 2128 1378 2132
rect 1398 2128 1402 2132
rect 1342 2118 1346 2122
rect 1390 2118 1394 2122
rect 1358 2108 1362 2112
rect 1334 2088 1338 2092
rect 1334 2068 1338 2072
rect 1454 2148 1458 2152
rect 1454 2108 1458 2112
rect 1422 2088 1426 2092
rect 1366 2078 1370 2082
rect 1406 2068 1410 2072
rect 1446 2068 1450 2072
rect 1310 2058 1314 2062
rect 1366 2058 1370 2062
rect 1382 2058 1386 2062
rect 1430 2058 1434 2062
rect 1230 2018 1234 2022
rect 1166 2008 1170 2012
rect 1158 1988 1162 1992
rect 1206 1988 1210 1992
rect 1214 1978 1218 1982
rect 1158 1968 1162 1972
rect 1190 1948 1194 1952
rect 1150 1898 1154 1902
rect 1142 1878 1146 1882
rect 1126 1868 1130 1872
rect 1118 1858 1122 1862
rect 1126 1858 1130 1862
rect 1158 1858 1162 1862
rect 1094 1848 1098 1852
rect 1126 1848 1130 1852
rect 1142 1808 1146 1812
rect 1094 1798 1098 1802
rect 1102 1768 1106 1772
rect 1086 1758 1090 1762
rect 1054 1738 1058 1742
rect 1070 1738 1074 1742
rect 1094 1738 1098 1742
rect 990 1728 994 1732
rect 974 1698 978 1702
rect 1014 1698 1018 1702
rect 1262 1948 1266 1952
rect 1198 1938 1202 1942
rect 1214 1938 1218 1942
rect 1246 1938 1250 1942
rect 1182 1928 1186 1932
rect 1206 1858 1210 1862
rect 1358 2038 1362 2042
rect 1390 2038 1394 2042
rect 1294 2028 1298 2032
rect 1354 2003 1358 2007
rect 1361 2003 1365 2007
rect 1342 1978 1346 1982
rect 1318 1958 1322 1962
rect 1374 1958 1378 1962
rect 1350 1938 1354 1942
rect 1406 2028 1410 2032
rect 1422 2028 1426 2032
rect 1422 2008 1426 2012
rect 1398 1968 1402 1972
rect 1422 1968 1426 1972
rect 1446 2038 1450 2042
rect 1558 2168 1562 2172
rect 1566 2168 1570 2172
rect 1590 2168 1594 2172
rect 1678 2168 1682 2172
rect 1702 2168 1706 2172
rect 1734 2198 1738 2202
rect 1726 2178 1730 2182
rect 1694 2158 1698 2162
rect 1758 2248 1762 2252
rect 1742 2178 1746 2182
rect 1750 2168 1754 2172
rect 1558 2148 1562 2152
rect 1566 2148 1570 2152
rect 1638 2148 1642 2152
rect 1734 2148 1738 2152
rect 1534 2138 1538 2142
rect 1606 2138 1610 2142
rect 1598 2128 1602 2132
rect 1662 2128 1666 2132
rect 1710 2128 1714 2132
rect 1542 2118 1546 2122
rect 1574 2118 1578 2122
rect 1598 2108 1602 2112
rect 1606 2098 1610 2102
rect 1582 2088 1586 2092
rect 1654 2118 1658 2122
rect 1494 2078 1498 2082
rect 1558 2078 1562 2082
rect 1614 2078 1618 2082
rect 1622 2078 1626 2082
rect 1646 2078 1650 2082
rect 1566 2068 1570 2072
rect 1574 2068 1578 2072
rect 1510 2058 1514 2062
rect 1550 2058 1554 2062
rect 1726 2108 1730 2112
rect 1734 2098 1738 2102
rect 1630 2058 1634 2062
rect 1662 2058 1666 2062
rect 1574 2048 1578 2052
rect 1534 2008 1538 2012
rect 1470 1998 1474 2002
rect 1518 1998 1522 2002
rect 1526 1978 1530 1982
rect 1566 1978 1570 1982
rect 1454 1968 1458 1972
rect 1406 1958 1410 1962
rect 1438 1958 1442 1962
rect 1446 1958 1450 1962
rect 1278 1918 1282 1922
rect 1310 1918 1314 1922
rect 1334 1918 1338 1922
rect 1270 1878 1274 1882
rect 1278 1868 1282 1872
rect 1398 1918 1402 1922
rect 1358 1898 1362 1902
rect 1366 1898 1370 1902
rect 1318 1878 1322 1882
rect 1350 1878 1354 1882
rect 1334 1868 1338 1872
rect 1294 1848 1298 1852
rect 1262 1838 1266 1842
rect 1190 1818 1194 1822
rect 1238 1818 1242 1822
rect 1158 1798 1162 1802
rect 1174 1798 1178 1802
rect 1182 1768 1186 1772
rect 1134 1748 1138 1752
rect 1158 1748 1162 1752
rect 1142 1738 1146 1742
rect 1174 1738 1178 1742
rect 1206 1768 1210 1772
rect 1374 1868 1378 1872
rect 1326 1848 1330 1852
rect 1342 1838 1346 1842
rect 1310 1798 1314 1802
rect 1286 1778 1290 1782
rect 1270 1748 1274 1752
rect 1222 1728 1226 1732
rect 1254 1728 1258 1732
rect 1110 1678 1114 1682
rect 1134 1678 1138 1682
rect 1046 1668 1050 1672
rect 1078 1668 1082 1672
rect 1110 1668 1114 1672
rect 1126 1668 1130 1672
rect 1126 1658 1130 1662
rect 1006 1648 1010 1652
rect 1054 1628 1058 1632
rect 1054 1598 1058 1602
rect 1014 1578 1018 1582
rect 1046 1568 1050 1572
rect 1134 1598 1138 1602
rect 1086 1578 1090 1582
rect 1134 1578 1138 1582
rect 1118 1568 1122 1572
rect 990 1548 994 1552
rect 1022 1548 1026 1552
rect 1078 1548 1082 1552
rect 1094 1548 1098 1552
rect 982 1538 986 1542
rect 1014 1538 1018 1542
rect 982 1458 986 1462
rect 1006 1448 1010 1452
rect 1014 1438 1018 1442
rect 1118 1538 1122 1542
rect 1102 1508 1106 1512
rect 1350 1828 1354 1832
rect 1342 1808 1346 1812
rect 1354 1803 1358 1807
rect 1361 1803 1365 1807
rect 1318 1748 1322 1752
rect 1326 1748 1330 1752
rect 1334 1738 1338 1742
rect 1318 1728 1322 1732
rect 1334 1688 1338 1692
rect 1302 1678 1306 1682
rect 1278 1668 1282 1672
rect 1326 1668 1330 1672
rect 1262 1658 1266 1662
rect 1438 1938 1442 1942
rect 1422 1918 1426 1922
rect 1406 1858 1410 1862
rect 1422 1828 1426 1832
rect 1430 1758 1434 1762
rect 1430 1748 1434 1752
rect 1406 1738 1410 1742
rect 1422 1738 1426 1742
rect 1374 1728 1378 1732
rect 1366 1678 1370 1682
rect 1358 1668 1362 1672
rect 1414 1718 1418 1722
rect 1406 1708 1410 1712
rect 1414 1698 1418 1702
rect 1406 1678 1410 1682
rect 1390 1658 1394 1662
rect 1310 1648 1314 1652
rect 1302 1618 1306 1622
rect 1278 1608 1282 1612
rect 1182 1588 1186 1592
rect 1166 1578 1170 1582
rect 1422 1668 1426 1672
rect 1430 1658 1434 1662
rect 1390 1608 1394 1612
rect 1354 1603 1358 1607
rect 1361 1603 1365 1607
rect 1406 1598 1410 1602
rect 1398 1578 1402 1582
rect 1342 1568 1346 1572
rect 1318 1558 1322 1562
rect 1358 1558 1362 1562
rect 1174 1548 1178 1552
rect 1286 1548 1290 1552
rect 1342 1548 1346 1552
rect 1158 1538 1162 1542
rect 1166 1538 1170 1542
rect 1246 1538 1250 1542
rect 1150 1528 1154 1532
rect 1142 1518 1146 1522
rect 1094 1478 1098 1482
rect 1046 1468 1050 1472
rect 1070 1458 1074 1462
rect 1102 1458 1106 1462
rect 1118 1458 1122 1462
rect 1174 1458 1178 1462
rect 1142 1448 1146 1452
rect 1054 1438 1058 1442
rect 1078 1438 1082 1442
rect 1126 1428 1130 1432
rect 1030 1418 1034 1422
rect 1134 1418 1138 1422
rect 1078 1408 1082 1412
rect 1102 1398 1106 1402
rect 1030 1388 1034 1392
rect 966 1378 970 1382
rect 1014 1368 1018 1372
rect 942 1348 946 1352
rect 974 1348 978 1352
rect 950 1338 954 1342
rect 850 1303 854 1307
rect 857 1303 861 1307
rect 870 1288 874 1292
rect 878 1288 882 1292
rect 790 1278 794 1282
rect 830 1278 834 1282
rect 822 1268 826 1272
rect 886 1268 890 1272
rect 902 1268 906 1272
rect 662 1258 666 1262
rect 758 1258 762 1262
rect 774 1258 778 1262
rect 806 1258 810 1262
rect 838 1258 842 1262
rect 638 1248 642 1252
rect 662 1248 666 1252
rect 638 1228 642 1232
rect 646 1228 650 1232
rect 574 1148 578 1152
rect 638 1148 642 1152
rect 646 1148 650 1152
rect 582 1128 586 1132
rect 558 1098 562 1102
rect 422 948 426 952
rect 550 948 554 952
rect 406 908 410 912
rect 398 848 402 852
rect 422 878 426 882
rect 462 928 466 932
rect 510 928 514 932
rect 446 908 450 912
rect 486 908 490 912
rect 486 878 490 882
rect 462 868 466 872
rect 430 848 434 852
rect 470 848 474 852
rect 422 838 426 842
rect 414 778 418 782
rect 406 768 410 772
rect 358 758 362 762
rect 358 748 362 752
rect 374 738 378 742
rect 390 718 394 722
rect 366 708 370 712
rect 366 698 370 702
rect 374 678 378 682
rect 390 678 394 682
rect 366 658 370 662
rect 390 648 394 652
rect 334 618 338 622
rect 330 603 334 607
rect 337 603 341 607
rect 358 578 362 582
rect 398 568 402 572
rect 302 548 306 552
rect 334 548 338 552
rect 358 548 362 552
rect 302 538 306 542
rect 382 528 386 532
rect 246 508 250 512
rect 246 498 250 502
rect 326 498 330 502
rect 166 478 170 482
rect 174 468 178 472
rect 310 488 314 492
rect 342 488 346 492
rect 326 468 330 472
rect 374 468 378 472
rect 198 458 202 462
rect 302 458 306 462
rect 150 448 154 452
rect 182 448 186 452
rect 198 448 202 452
rect 398 458 402 462
rect 382 438 386 442
rect 198 428 202 432
rect 390 408 394 412
rect 330 403 334 407
rect 337 403 341 407
rect 350 368 354 372
rect 214 358 218 362
rect 86 348 90 352
rect 222 348 226 352
rect 334 348 338 352
rect 62 338 66 342
rect 198 338 202 342
rect 206 338 210 342
rect 70 308 74 312
rect 94 308 98 312
rect 110 298 114 302
rect 166 298 170 302
rect 158 278 162 282
rect 142 268 146 272
rect 14 138 18 142
rect 62 248 66 252
rect 102 158 106 162
rect 86 148 90 152
rect 150 138 154 142
rect 54 108 58 112
rect 14 88 18 92
rect 70 78 74 82
rect 102 88 106 92
rect 126 78 130 82
rect 118 68 122 72
rect 150 68 154 72
rect 190 288 194 292
rect 214 288 218 292
rect 246 338 250 342
rect 310 338 314 342
rect 366 338 370 342
rect 262 328 266 332
rect 254 318 258 322
rect 254 268 258 272
rect 214 248 218 252
rect 206 188 210 192
rect 166 148 170 152
rect 182 128 186 132
rect 318 328 322 332
rect 366 328 370 332
rect 358 308 362 312
rect 366 308 370 312
rect 302 278 306 282
rect 382 288 386 292
rect 342 268 346 272
rect 286 258 290 262
rect 238 188 242 192
rect 270 168 274 172
rect 294 168 298 172
rect 502 848 506 852
rect 494 828 498 832
rect 486 808 490 812
rect 518 788 522 792
rect 502 758 506 762
rect 422 748 426 752
rect 454 748 458 752
rect 462 748 466 752
rect 542 868 546 872
rect 598 1088 602 1092
rect 646 1088 650 1092
rect 614 1068 618 1072
rect 630 1068 634 1072
rect 622 1058 626 1062
rect 574 1048 578 1052
rect 598 1048 602 1052
rect 566 968 570 972
rect 630 988 634 992
rect 670 1158 674 1162
rect 726 1158 730 1162
rect 726 1148 730 1152
rect 694 1138 698 1142
rect 718 1138 722 1142
rect 694 1118 698 1122
rect 702 1108 706 1112
rect 686 1088 690 1092
rect 678 1068 682 1072
rect 654 1048 658 1052
rect 662 1048 666 1052
rect 670 988 674 992
rect 646 978 650 982
rect 582 948 586 952
rect 598 948 602 952
rect 654 958 658 962
rect 598 928 602 932
rect 630 928 634 932
rect 646 928 650 932
rect 574 908 578 912
rect 606 898 610 902
rect 630 898 634 902
rect 590 868 594 872
rect 582 858 586 862
rect 550 848 554 852
rect 614 868 618 872
rect 622 858 626 862
rect 654 908 658 912
rect 646 888 650 892
rect 638 868 642 872
rect 614 798 618 802
rect 630 798 634 802
rect 622 768 626 772
rect 574 748 578 752
rect 462 738 466 742
rect 478 728 482 732
rect 470 718 474 722
rect 478 708 482 712
rect 494 718 498 722
rect 486 698 490 702
rect 510 708 514 712
rect 478 688 482 692
rect 446 678 450 682
rect 558 698 562 702
rect 534 678 538 682
rect 486 648 490 652
rect 494 638 498 642
rect 486 608 490 612
rect 454 588 458 592
rect 606 688 610 692
rect 662 898 666 902
rect 662 878 666 882
rect 686 978 690 982
rect 974 1318 978 1322
rect 926 1308 930 1312
rect 942 1268 946 1272
rect 950 1268 954 1272
rect 966 1268 970 1272
rect 902 1248 906 1252
rect 886 1218 890 1222
rect 838 1208 842 1212
rect 830 1198 834 1202
rect 878 1188 882 1192
rect 814 1168 818 1172
rect 830 1168 834 1172
rect 822 1158 826 1162
rect 806 1148 810 1152
rect 758 1138 762 1142
rect 782 1128 786 1132
rect 814 1128 818 1132
rect 774 1098 778 1102
rect 798 1098 802 1102
rect 798 1088 802 1092
rect 814 1068 818 1072
rect 798 1038 802 1042
rect 814 1028 818 1032
rect 718 988 722 992
rect 750 988 754 992
rect 734 958 738 962
rect 678 948 682 952
rect 694 948 698 952
rect 718 888 722 892
rect 710 878 714 882
rect 646 758 650 762
rect 678 858 682 862
rect 710 858 714 862
rect 670 848 674 852
rect 718 848 722 852
rect 710 818 714 822
rect 662 778 666 782
rect 710 728 714 732
rect 638 698 642 702
rect 814 958 818 962
rect 766 878 770 882
rect 782 878 786 882
rect 798 858 802 862
rect 758 838 762 842
rect 726 718 730 722
rect 758 748 762 752
rect 774 748 778 752
rect 750 738 754 742
rect 766 738 770 742
rect 798 828 802 832
rect 798 748 802 752
rect 846 1148 850 1152
rect 830 1068 834 1072
rect 886 1128 890 1132
rect 850 1103 854 1107
rect 857 1103 861 1107
rect 878 1068 882 1072
rect 838 1018 842 1022
rect 830 958 834 962
rect 850 903 854 907
rect 857 903 861 907
rect 822 898 826 902
rect 830 868 834 872
rect 814 858 818 862
rect 862 858 866 862
rect 830 848 834 852
rect 846 838 850 842
rect 822 798 826 802
rect 950 1218 954 1222
rect 926 1208 930 1212
rect 958 1208 962 1212
rect 918 1178 922 1182
rect 902 1168 906 1172
rect 910 1158 914 1162
rect 926 1148 930 1152
rect 982 1308 986 1312
rect 982 1298 986 1302
rect 990 1278 994 1282
rect 990 1218 994 1222
rect 982 1208 986 1212
rect 990 1148 994 1152
rect 1014 1268 1018 1272
rect 1014 1208 1018 1212
rect 1022 1168 1026 1172
rect 1118 1388 1122 1392
rect 1086 1368 1090 1372
rect 1118 1368 1122 1372
rect 1038 1358 1042 1362
rect 1046 1358 1050 1362
rect 1038 1338 1042 1342
rect 1054 1338 1058 1342
rect 1038 1328 1042 1332
rect 1150 1388 1154 1392
rect 1158 1388 1162 1392
rect 1174 1378 1178 1382
rect 1134 1358 1138 1362
rect 1142 1358 1146 1362
rect 1214 1498 1218 1502
rect 1246 1468 1250 1472
rect 1326 1538 1330 1542
rect 1294 1528 1298 1532
rect 1310 1488 1314 1492
rect 1262 1458 1266 1462
rect 1334 1468 1338 1472
rect 1334 1458 1338 1462
rect 1350 1458 1354 1462
rect 1222 1448 1226 1452
rect 1238 1448 1242 1452
rect 1254 1448 1258 1452
rect 1294 1448 1298 1452
rect 1214 1438 1218 1442
rect 1198 1358 1202 1362
rect 1206 1358 1210 1362
rect 1254 1438 1258 1442
rect 1230 1408 1234 1412
rect 1302 1428 1306 1432
rect 1406 1558 1410 1562
rect 1414 1558 1418 1562
rect 1366 1448 1370 1452
rect 1342 1428 1346 1432
rect 1354 1403 1358 1407
rect 1361 1403 1365 1407
rect 1318 1388 1322 1392
rect 1342 1388 1346 1392
rect 1374 1378 1378 1382
rect 1166 1348 1170 1352
rect 1222 1348 1226 1352
rect 1238 1338 1242 1342
rect 1246 1338 1250 1342
rect 1302 1338 1306 1342
rect 1118 1328 1122 1332
rect 1062 1318 1066 1322
rect 1286 1328 1290 1332
rect 1302 1328 1306 1332
rect 1070 1298 1074 1302
rect 1046 1278 1050 1282
rect 1086 1268 1090 1272
rect 1094 1268 1098 1272
rect 1054 1218 1058 1222
rect 1062 1218 1066 1222
rect 1046 1158 1050 1162
rect 1094 1198 1098 1202
rect 1270 1308 1274 1312
rect 1198 1298 1202 1302
rect 1334 1318 1338 1322
rect 1350 1318 1354 1322
rect 1310 1308 1314 1312
rect 1302 1268 1306 1272
rect 1142 1259 1146 1263
rect 1318 1268 1322 1272
rect 1398 1388 1402 1392
rect 1382 1298 1386 1302
rect 1390 1298 1394 1302
rect 1558 1968 1562 1972
rect 1686 2038 1690 2042
rect 1614 2028 1618 2032
rect 1582 1988 1586 1992
rect 1726 2048 1730 2052
rect 1694 2008 1698 2012
rect 1726 1998 1730 2002
rect 1614 1968 1618 1972
rect 1910 2288 1914 2292
rect 1934 2448 1938 2452
rect 1966 2438 1970 2442
rect 1966 2398 1970 2402
rect 1958 2358 1962 2362
rect 1966 2358 1970 2362
rect 1934 2348 1938 2352
rect 1934 2318 1938 2322
rect 2038 2518 2042 2522
rect 2014 2498 2018 2502
rect 1998 2488 2002 2492
rect 2062 2488 2066 2492
rect 1990 2468 1994 2472
rect 2014 2468 2018 2472
rect 2030 2468 2034 2472
rect 2054 2448 2058 2452
rect 2054 2418 2058 2422
rect 1982 2398 1986 2402
rect 2022 2398 2026 2402
rect 2326 2898 2330 2902
rect 2342 2938 2346 2942
rect 2350 2908 2354 2912
rect 2342 2878 2346 2882
rect 2342 2828 2346 2832
rect 2270 2738 2274 2742
rect 2278 2738 2282 2742
rect 2342 2738 2346 2742
rect 2246 2698 2250 2702
rect 2326 2688 2330 2692
rect 2262 2658 2266 2662
rect 2190 2628 2194 2632
rect 2190 2608 2194 2612
rect 2238 2608 2242 2612
rect 2142 2548 2146 2552
rect 2182 2548 2186 2552
rect 2126 2528 2130 2532
rect 2102 2518 2106 2522
rect 2094 2508 2098 2512
rect 2094 2498 2098 2502
rect 2238 2598 2242 2602
rect 2198 2568 2202 2572
rect 2254 2568 2258 2572
rect 2118 2478 2122 2482
rect 2118 2458 2122 2462
rect 2134 2458 2138 2462
rect 2158 2458 2162 2462
rect 2102 2448 2106 2452
rect 2126 2448 2130 2452
rect 2134 2438 2138 2442
rect 2142 2438 2146 2442
rect 2182 2448 2186 2452
rect 2174 2418 2178 2422
rect 2118 2408 2122 2412
rect 2158 2398 2162 2402
rect 2166 2398 2170 2402
rect 2134 2378 2138 2382
rect 2022 2358 2026 2362
rect 2070 2358 2074 2362
rect 2078 2358 2082 2362
rect 2046 2348 2050 2352
rect 2078 2348 2082 2352
rect 1974 2328 1978 2332
rect 1974 2318 1978 2322
rect 1966 2288 1970 2292
rect 1990 2288 1994 2292
rect 1910 2278 1914 2282
rect 1894 2198 1898 2202
rect 1838 2168 1842 2172
rect 1910 2168 1914 2172
rect 1846 2158 1850 2162
rect 1894 2158 1898 2162
rect 1910 2158 1914 2162
rect 1862 2148 1866 2152
rect 1886 2148 1890 2152
rect 1902 2138 1906 2142
rect 1910 2138 1914 2142
rect 1838 2128 1842 2132
rect 1798 2108 1802 2112
rect 1790 2088 1794 2092
rect 1766 2078 1770 2082
rect 1582 1948 1586 1952
rect 1606 1948 1610 1952
rect 1630 1948 1634 1952
rect 1694 1948 1698 1952
rect 1702 1948 1706 1952
rect 1470 1918 1474 1922
rect 1542 1928 1546 1932
rect 1598 1928 1602 1932
rect 1526 1898 1530 1902
rect 1550 1878 1554 1882
rect 1566 1878 1570 1882
rect 1558 1868 1562 1872
rect 1622 1938 1626 1942
rect 1654 1938 1658 1942
rect 1710 1938 1714 1942
rect 1726 1938 1730 1942
rect 1638 1928 1642 1932
rect 1702 1928 1706 1932
rect 1718 1918 1722 1922
rect 1670 1898 1674 1902
rect 1718 1888 1722 1892
rect 1614 1878 1618 1882
rect 1622 1878 1626 1882
rect 1726 1878 1730 1882
rect 1606 1868 1610 1872
rect 1526 1858 1530 1862
rect 1542 1858 1546 1862
rect 1574 1858 1578 1862
rect 1582 1858 1586 1862
rect 1462 1818 1466 1822
rect 1606 1848 1610 1852
rect 1590 1838 1594 1842
rect 1614 1818 1618 1822
rect 1558 1768 1562 1772
rect 1510 1758 1514 1762
rect 1558 1758 1562 1762
rect 1518 1698 1522 1702
rect 1462 1668 1466 1672
rect 1494 1668 1498 1672
rect 1510 1658 1514 1662
rect 1494 1648 1498 1652
rect 1486 1608 1490 1612
rect 1462 1558 1466 1562
rect 1478 1558 1482 1562
rect 1462 1538 1466 1542
rect 1454 1528 1458 1532
rect 1494 1568 1498 1572
rect 1510 1558 1514 1562
rect 1550 1748 1554 1752
rect 1542 1738 1546 1742
rect 1582 1738 1586 1742
rect 1526 1608 1530 1612
rect 1550 1598 1554 1602
rect 1574 1668 1578 1672
rect 1574 1659 1578 1663
rect 1558 1568 1562 1572
rect 1574 1568 1578 1572
rect 1582 1548 1586 1552
rect 1494 1538 1498 1542
rect 1534 1538 1538 1542
rect 1518 1528 1522 1532
rect 1478 1488 1482 1492
rect 1742 1868 1746 1872
rect 1662 1858 1666 1862
rect 1694 1848 1698 1852
rect 1718 1848 1722 1852
rect 1678 1818 1682 1822
rect 1670 1808 1674 1812
rect 1654 1748 1658 1752
rect 1630 1708 1634 1712
rect 1622 1698 1626 1702
rect 1750 1838 1754 1842
rect 1726 1768 1730 1772
rect 1734 1768 1738 1772
rect 1710 1758 1714 1762
rect 1758 1758 1762 1762
rect 1710 1748 1714 1752
rect 1774 2068 1778 2072
rect 1874 2103 1878 2107
rect 1881 2103 1885 2107
rect 1902 2098 1906 2102
rect 1862 2088 1866 2092
rect 1870 2068 1874 2072
rect 1894 2068 1898 2072
rect 1958 2268 1962 2272
rect 1934 2258 1938 2262
rect 1950 2258 1954 2262
rect 1926 2198 1930 2202
rect 2006 2268 2010 2272
rect 1974 2258 1978 2262
rect 1990 2208 1994 2212
rect 1950 2188 1954 2192
rect 1974 2188 1978 2192
rect 1990 2178 1994 2182
rect 1958 2158 1962 2162
rect 1982 2148 1986 2152
rect 1926 2138 1930 2142
rect 1958 2138 1962 2142
rect 1942 2128 1946 2132
rect 1934 2108 1938 2112
rect 1974 2108 1978 2112
rect 1982 2108 1986 2112
rect 1966 2098 1970 2102
rect 1966 2088 1970 2092
rect 1918 2078 1922 2082
rect 1926 2078 1930 2082
rect 1982 2078 1986 2082
rect 1982 2068 1986 2072
rect 1846 2058 1850 2062
rect 1830 2048 1834 2052
rect 1838 2048 1842 2052
rect 1846 2038 1850 2042
rect 1854 2038 1858 2042
rect 1814 2028 1818 2032
rect 1790 1988 1794 1992
rect 1774 1968 1778 1972
rect 1774 1898 1778 1902
rect 1774 1858 1778 1862
rect 1798 1968 1802 1972
rect 1838 1988 1842 1992
rect 1862 1988 1866 1992
rect 1830 1968 1834 1972
rect 1918 2048 1922 2052
rect 1926 2048 1930 2052
rect 1942 2048 1946 2052
rect 1982 2048 1986 2052
rect 1950 2038 1954 2042
rect 1974 2038 1978 2042
rect 1934 2028 1938 2032
rect 1902 1988 1906 1992
rect 1870 1968 1874 1972
rect 1854 1948 1858 1952
rect 1870 1948 1874 1952
rect 1790 1878 1794 1882
rect 1814 1818 1818 1822
rect 1798 1768 1802 1772
rect 1798 1748 1802 1752
rect 1678 1738 1682 1742
rect 1718 1738 1722 1742
rect 1766 1738 1770 1742
rect 1734 1718 1738 1722
rect 1686 1708 1690 1712
rect 1670 1678 1674 1682
rect 1654 1668 1658 1672
rect 1638 1658 1642 1662
rect 1622 1648 1626 1652
rect 1678 1648 1682 1652
rect 1710 1688 1714 1692
rect 1718 1688 1722 1692
rect 1718 1648 1722 1652
rect 1702 1638 1706 1642
rect 1686 1608 1690 1612
rect 1694 1608 1698 1612
rect 1678 1598 1682 1602
rect 1662 1568 1666 1572
rect 1622 1558 1626 1562
rect 1646 1558 1650 1562
rect 1558 1538 1562 1542
rect 1662 1538 1666 1542
rect 1542 1508 1546 1512
rect 1502 1468 1506 1472
rect 1446 1448 1450 1452
rect 1454 1448 1458 1452
rect 1430 1428 1434 1432
rect 1438 1428 1442 1432
rect 1462 1408 1466 1412
rect 1422 1388 1426 1392
rect 1430 1388 1434 1392
rect 1486 1388 1490 1392
rect 1510 1388 1514 1392
rect 1470 1348 1474 1352
rect 1526 1408 1530 1412
rect 1534 1398 1538 1402
rect 1422 1338 1426 1342
rect 1518 1338 1522 1342
rect 1406 1308 1410 1312
rect 1414 1308 1418 1312
rect 1358 1278 1362 1282
rect 1390 1278 1394 1282
rect 1406 1278 1410 1282
rect 1382 1268 1386 1272
rect 1166 1258 1170 1262
rect 1214 1258 1218 1262
rect 1246 1258 1250 1262
rect 1118 1228 1122 1232
rect 1102 1188 1106 1192
rect 1094 1168 1098 1172
rect 1118 1168 1122 1172
rect 1070 1158 1074 1162
rect 998 1128 1002 1132
rect 1006 1128 1010 1132
rect 1070 1138 1074 1142
rect 1102 1138 1106 1142
rect 1150 1158 1154 1162
rect 1294 1248 1298 1252
rect 1222 1168 1226 1172
rect 1062 1118 1066 1122
rect 1086 1098 1090 1102
rect 966 1078 970 1082
rect 990 1078 994 1082
rect 1006 1078 1010 1082
rect 1038 1078 1042 1082
rect 1062 1078 1066 1082
rect 1102 1078 1106 1082
rect 1014 1058 1018 1062
rect 1046 1058 1050 1062
rect 1070 1058 1074 1062
rect 1030 1048 1034 1052
rect 966 1038 970 1042
rect 998 1038 1002 1042
rect 918 1018 922 1022
rect 894 1008 898 1012
rect 950 998 954 1002
rect 1046 1028 1050 1032
rect 982 968 986 972
rect 958 958 962 962
rect 974 958 978 962
rect 902 948 906 952
rect 934 938 938 942
rect 894 928 898 932
rect 1030 958 1034 962
rect 1118 1028 1122 1032
rect 1094 988 1098 992
rect 966 948 970 952
rect 1038 948 1042 952
rect 1046 948 1050 952
rect 1062 948 1066 952
rect 958 938 962 942
rect 886 918 890 922
rect 894 918 898 922
rect 886 898 890 902
rect 878 878 882 882
rect 918 898 922 902
rect 974 918 978 922
rect 958 878 962 882
rect 934 868 938 872
rect 926 858 930 862
rect 942 858 946 862
rect 902 848 906 852
rect 918 828 922 832
rect 902 808 906 812
rect 910 808 914 812
rect 854 758 858 762
rect 870 758 874 762
rect 814 748 818 752
rect 758 728 762 732
rect 782 728 786 732
rect 670 688 674 692
rect 726 688 730 692
rect 670 668 674 672
rect 630 658 634 662
rect 646 658 650 662
rect 614 628 618 632
rect 518 608 522 612
rect 542 608 546 612
rect 582 578 586 582
rect 542 558 546 562
rect 502 548 506 552
rect 502 528 506 532
rect 542 498 546 502
rect 518 488 522 492
rect 566 518 570 522
rect 550 478 554 482
rect 494 468 498 472
rect 518 468 522 472
rect 542 468 546 472
rect 422 458 426 462
rect 526 458 530 462
rect 406 448 410 452
rect 414 378 418 382
rect 406 368 410 372
rect 406 358 410 362
rect 398 338 402 342
rect 406 288 410 292
rect 438 368 442 372
rect 454 358 458 362
rect 470 348 474 352
rect 454 338 458 342
rect 438 288 442 292
rect 446 278 450 282
rect 422 268 426 272
rect 438 268 442 272
rect 502 318 506 322
rect 486 308 490 312
rect 454 268 458 272
rect 486 268 490 272
rect 390 258 394 262
rect 330 203 334 207
rect 337 203 341 207
rect 414 248 418 252
rect 454 248 458 252
rect 174 98 178 102
rect 198 98 202 102
rect 222 98 226 102
rect 214 88 218 92
rect 302 88 306 92
rect 430 158 434 162
rect 462 158 466 162
rect 390 148 394 152
rect 406 148 410 152
rect 438 148 442 152
rect 446 138 450 142
rect 134 58 138 62
rect 166 58 170 62
rect 190 58 194 62
rect 454 118 458 122
rect 422 98 426 102
rect 446 98 450 102
rect 534 258 538 262
rect 550 448 554 452
rect 550 398 554 402
rect 590 459 594 463
rect 582 338 586 342
rect 606 278 610 282
rect 566 268 570 272
rect 662 648 666 652
rect 646 638 650 642
rect 646 618 650 622
rect 734 678 738 682
rect 758 678 762 682
rect 710 658 714 662
rect 710 648 714 652
rect 678 638 682 642
rect 662 558 666 562
rect 822 728 826 732
rect 838 728 842 732
rect 806 708 810 712
rect 830 708 834 712
rect 798 628 802 632
rect 742 608 746 612
rect 878 718 882 722
rect 850 703 854 707
rect 857 703 861 707
rect 878 688 882 692
rect 870 658 874 662
rect 838 628 842 632
rect 774 578 778 582
rect 766 568 770 572
rect 662 548 666 552
rect 646 528 650 532
rect 630 498 634 502
rect 702 518 706 522
rect 694 508 698 512
rect 686 498 690 502
rect 710 508 714 512
rect 814 558 818 562
rect 846 608 850 612
rect 854 568 858 572
rect 870 578 874 582
rect 798 548 802 552
rect 862 548 866 552
rect 790 538 794 542
rect 806 538 810 542
rect 790 518 794 522
rect 798 518 802 522
rect 742 488 746 492
rect 678 468 682 472
rect 734 468 738 472
rect 686 458 690 462
rect 678 378 682 382
rect 654 368 658 372
rect 774 478 778 482
rect 742 448 746 452
rect 750 448 754 452
rect 766 438 770 442
rect 750 388 754 392
rect 758 388 762 392
rect 726 378 730 382
rect 750 368 754 372
rect 710 338 714 342
rect 638 328 642 332
rect 646 308 650 312
rect 814 478 818 482
rect 806 388 810 392
rect 850 503 854 507
rect 857 503 861 507
rect 854 488 858 492
rect 830 438 834 442
rect 886 648 890 652
rect 902 638 906 642
rect 894 558 898 562
rect 982 888 986 892
rect 982 798 986 802
rect 934 758 938 762
rect 926 728 930 732
rect 918 558 922 562
rect 886 538 890 542
rect 886 468 890 472
rect 878 428 882 432
rect 942 718 946 722
rect 998 758 1002 762
rect 1046 898 1050 902
rect 1046 878 1050 882
rect 1118 958 1122 962
rect 1102 948 1106 952
rect 1134 948 1138 952
rect 1078 938 1082 942
rect 1070 888 1074 892
rect 1118 928 1122 932
rect 1118 878 1122 882
rect 1062 858 1066 862
rect 1094 848 1098 852
rect 1078 828 1082 832
rect 1014 778 1018 782
rect 1046 778 1050 782
rect 982 728 986 732
rect 990 728 994 732
rect 966 668 970 672
rect 1038 758 1042 762
rect 998 658 1002 662
rect 942 548 946 552
rect 1014 628 1018 632
rect 982 568 986 572
rect 974 548 978 552
rect 958 528 962 532
rect 942 498 946 502
rect 934 488 938 492
rect 910 478 914 482
rect 966 478 970 482
rect 950 458 954 462
rect 982 458 986 462
rect 942 448 946 452
rect 950 448 954 452
rect 942 438 946 442
rect 942 418 946 422
rect 958 418 962 422
rect 902 398 906 402
rect 934 398 938 402
rect 838 388 842 392
rect 798 358 802 362
rect 822 358 826 362
rect 750 288 754 292
rect 662 278 666 282
rect 686 268 690 272
rect 774 268 778 272
rect 638 248 642 252
rect 646 248 650 252
rect 598 238 602 242
rect 550 148 554 152
rect 566 148 570 152
rect 630 148 634 152
rect 542 128 546 132
rect 518 118 522 122
rect 550 118 554 122
rect 598 118 602 122
rect 606 118 610 122
rect 542 108 546 112
rect 558 78 562 82
rect 662 148 666 152
rect 910 368 914 372
rect 1054 748 1058 752
rect 1078 747 1082 751
rect 1054 718 1058 722
rect 1086 688 1090 692
rect 1118 838 1122 842
rect 1182 1098 1186 1102
rect 1222 1158 1226 1162
rect 1286 1158 1290 1162
rect 1222 1138 1226 1142
rect 1222 1068 1226 1072
rect 1190 1028 1194 1032
rect 1342 1248 1346 1252
rect 1358 1248 1362 1252
rect 1350 1228 1354 1232
rect 1354 1203 1358 1207
rect 1361 1203 1365 1207
rect 1374 1198 1378 1202
rect 1310 1188 1314 1192
rect 1326 1188 1330 1192
rect 1350 1168 1354 1172
rect 1318 1158 1322 1162
rect 1302 1148 1306 1152
rect 1334 1148 1338 1152
rect 1270 1128 1274 1132
rect 1294 1118 1298 1122
rect 1254 1108 1258 1112
rect 1278 1108 1282 1112
rect 1270 1038 1274 1042
rect 1238 998 1242 1002
rect 1318 1068 1322 1072
rect 1294 1058 1298 1062
rect 1294 1048 1298 1052
rect 1310 1048 1314 1052
rect 1286 1008 1290 1012
rect 1222 988 1226 992
rect 1238 988 1242 992
rect 1278 988 1282 992
rect 1158 968 1162 972
rect 1166 958 1170 962
rect 1174 958 1178 962
rect 1262 958 1266 962
rect 1222 938 1226 942
rect 1198 918 1202 922
rect 1198 878 1202 882
rect 1246 928 1250 932
rect 1222 898 1226 902
rect 1142 868 1146 872
rect 1214 848 1218 852
rect 1134 828 1138 832
rect 1166 828 1170 832
rect 1094 678 1098 682
rect 1046 668 1050 672
rect 1054 668 1058 672
rect 1062 658 1066 662
rect 1006 578 1010 582
rect 1022 578 1026 582
rect 1014 558 1018 562
rect 1150 758 1154 762
rect 1230 888 1234 892
rect 1246 868 1250 872
rect 1270 948 1274 952
rect 1270 888 1274 892
rect 1254 858 1258 862
rect 1262 858 1266 862
rect 1334 948 1338 952
rect 1318 938 1322 942
rect 1334 888 1338 892
rect 1326 878 1330 882
rect 1238 848 1242 852
rect 1246 848 1250 852
rect 1238 818 1242 822
rect 1190 778 1194 782
rect 1190 758 1194 762
rect 1198 758 1202 762
rect 1262 778 1266 782
rect 1230 748 1234 752
rect 1414 1268 1418 1272
rect 1398 1258 1402 1262
rect 1414 1228 1418 1232
rect 1406 1158 1410 1162
rect 1390 1148 1394 1152
rect 1406 1148 1410 1152
rect 1526 1278 1530 1282
rect 1550 1468 1554 1472
rect 1582 1518 1586 1522
rect 1598 1488 1602 1492
rect 1750 1678 1754 1682
rect 1766 1678 1770 1682
rect 1942 2008 1946 2012
rect 2006 2218 2010 2222
rect 1998 2088 2002 2092
rect 2038 2318 2042 2322
rect 2054 2268 2058 2272
rect 2022 2258 2026 2262
rect 2022 2238 2026 2242
rect 2030 2128 2034 2132
rect 2038 2068 2042 2072
rect 2070 2318 2074 2322
rect 2070 2248 2074 2252
rect 2182 2378 2186 2382
rect 2166 2368 2170 2372
rect 2126 2328 2130 2332
rect 2118 2298 2122 2302
rect 2222 2548 2226 2552
rect 2254 2548 2258 2552
rect 2286 2648 2290 2652
rect 2270 2568 2274 2572
rect 2286 2568 2290 2572
rect 2214 2538 2218 2542
rect 2206 2528 2210 2532
rect 2278 2518 2282 2522
rect 2230 2508 2234 2512
rect 2222 2458 2226 2462
rect 2214 2408 2218 2412
rect 2198 2388 2202 2392
rect 2190 2358 2194 2362
rect 2174 2338 2178 2342
rect 2150 2308 2154 2312
rect 2118 2278 2122 2282
rect 2102 2238 2106 2242
rect 2190 2308 2194 2312
rect 2174 2298 2178 2302
rect 2158 2288 2162 2292
rect 2134 2258 2138 2262
rect 2150 2248 2154 2252
rect 2102 2168 2106 2172
rect 2094 2158 2098 2162
rect 2086 2108 2090 2112
rect 2062 2058 2066 2062
rect 2078 2058 2082 2062
rect 2014 2048 2018 2052
rect 2030 2038 2034 2042
rect 2030 2028 2034 2032
rect 2006 2008 2010 2012
rect 1998 1968 2002 1972
rect 1886 1938 1890 1942
rect 1894 1938 1898 1942
rect 1974 1938 1978 1942
rect 1870 1928 1874 1932
rect 1894 1928 1898 1932
rect 1926 1928 1930 1932
rect 1950 1928 1954 1932
rect 1874 1903 1878 1907
rect 1881 1903 1885 1907
rect 1926 1898 1930 1902
rect 2070 1968 2074 1972
rect 2078 1968 2082 1972
rect 2054 1958 2058 1962
rect 2006 1948 2010 1952
rect 2022 1948 2026 1952
rect 2078 1948 2082 1952
rect 2014 1938 2018 1942
rect 2006 1928 2010 1932
rect 1862 1878 1866 1882
rect 1990 1878 1994 1882
rect 1854 1868 1858 1872
rect 1846 1858 1850 1862
rect 1838 1798 1842 1802
rect 1790 1738 1794 1742
rect 1830 1738 1834 1742
rect 1806 1688 1810 1692
rect 1830 1718 1834 1722
rect 1742 1658 1746 1662
rect 1782 1658 1786 1662
rect 1734 1608 1738 1612
rect 1726 1598 1730 1602
rect 1710 1578 1714 1582
rect 1638 1498 1642 1502
rect 1702 1498 1706 1502
rect 1574 1468 1578 1472
rect 1630 1468 1634 1472
rect 1558 1448 1562 1452
rect 1558 1428 1562 1432
rect 1566 1428 1570 1432
rect 1590 1428 1594 1432
rect 1694 1488 1698 1492
rect 1718 1568 1722 1572
rect 1734 1568 1738 1572
rect 1726 1548 1730 1552
rect 1758 1648 1762 1652
rect 1758 1608 1762 1612
rect 1814 1608 1818 1612
rect 1750 1598 1754 1602
rect 1718 1528 1722 1532
rect 1734 1528 1738 1532
rect 1750 1498 1754 1502
rect 1798 1598 1802 1602
rect 1782 1568 1786 1572
rect 1774 1558 1778 1562
rect 1766 1538 1770 1542
rect 1774 1528 1778 1532
rect 1766 1508 1770 1512
rect 1782 1508 1786 1512
rect 1758 1488 1762 1492
rect 1726 1478 1730 1482
rect 1694 1468 1698 1472
rect 1734 1468 1738 1472
rect 1750 1468 1754 1472
rect 1694 1448 1698 1452
rect 1630 1388 1634 1392
rect 1582 1358 1586 1362
rect 1606 1358 1610 1362
rect 1622 1358 1626 1362
rect 1686 1358 1690 1362
rect 1702 1348 1706 1352
rect 1566 1338 1570 1342
rect 1598 1338 1602 1342
rect 1614 1338 1618 1342
rect 1638 1338 1642 1342
rect 1654 1338 1658 1342
rect 1718 1338 1722 1342
rect 1582 1328 1586 1332
rect 1646 1328 1650 1332
rect 1702 1328 1706 1332
rect 1614 1318 1618 1322
rect 1606 1308 1610 1312
rect 1598 1298 1602 1302
rect 1678 1298 1682 1302
rect 1430 1248 1434 1252
rect 1438 1158 1442 1162
rect 1430 1148 1434 1152
rect 1366 1078 1370 1082
rect 1382 1068 1386 1072
rect 1422 1068 1426 1072
rect 1390 1058 1394 1062
rect 1354 1003 1358 1007
rect 1361 1003 1365 1007
rect 1430 1048 1434 1052
rect 1406 1038 1410 1042
rect 1430 1038 1434 1042
rect 1406 1008 1410 1012
rect 1302 838 1306 842
rect 1294 788 1298 792
rect 1286 778 1290 782
rect 1326 768 1330 772
rect 1422 988 1426 992
rect 1414 958 1418 962
rect 1430 948 1434 952
rect 1422 878 1426 882
rect 1414 858 1418 862
rect 1374 828 1378 832
rect 1354 803 1358 807
rect 1361 803 1365 807
rect 1406 798 1410 802
rect 1382 788 1386 792
rect 1422 758 1426 762
rect 1278 748 1282 752
rect 1334 748 1338 752
rect 1182 728 1186 732
rect 1206 728 1210 732
rect 1230 728 1234 732
rect 1254 728 1258 732
rect 1142 688 1146 692
rect 1230 718 1234 722
rect 1206 678 1210 682
rect 1142 668 1146 672
rect 1174 668 1178 672
rect 1198 668 1202 672
rect 1222 658 1226 662
rect 1062 588 1066 592
rect 1070 588 1074 592
rect 1238 578 1242 582
rect 1046 568 1050 572
rect 1230 558 1234 562
rect 1238 558 1242 562
rect 1030 548 1034 552
rect 1038 548 1042 552
rect 1086 548 1090 552
rect 1030 538 1034 542
rect 1110 538 1114 542
rect 1134 538 1138 542
rect 1150 538 1154 542
rect 1054 528 1058 532
rect 1022 518 1026 522
rect 1118 518 1122 522
rect 1038 468 1042 472
rect 1158 528 1162 532
rect 1230 518 1234 522
rect 1150 488 1154 492
rect 1206 478 1210 482
rect 1054 458 1058 462
rect 1126 458 1130 462
rect 1190 459 1194 463
rect 998 448 1002 452
rect 1102 448 1106 452
rect 1014 428 1018 432
rect 1062 428 1066 432
rect 1006 358 1010 362
rect 814 338 818 342
rect 926 338 930 342
rect 990 338 994 342
rect 886 318 890 322
rect 850 303 854 307
rect 857 303 861 307
rect 822 298 826 302
rect 886 278 890 282
rect 806 268 810 272
rect 822 268 826 272
rect 862 268 866 272
rect 878 268 882 272
rect 798 258 802 262
rect 822 258 826 262
rect 718 218 722 222
rect 694 168 698 172
rect 718 168 722 172
rect 838 168 842 172
rect 670 128 674 132
rect 662 78 666 82
rect 702 118 706 122
rect 734 138 738 142
rect 726 118 730 122
rect 830 118 834 122
rect 710 98 714 102
rect 686 68 690 72
rect 374 58 378 62
rect 414 58 418 62
rect 630 58 634 62
rect 678 58 682 62
rect 246 48 250 52
rect 630 48 634 52
rect 646 48 650 52
rect 850 103 854 107
rect 857 103 861 107
rect 798 78 802 82
rect 926 308 930 312
rect 918 278 922 282
rect 894 238 898 242
rect 886 158 890 162
rect 950 318 954 322
rect 990 318 994 322
rect 950 298 954 302
rect 982 298 986 302
rect 942 248 946 252
rect 1046 288 1050 292
rect 1038 268 1042 272
rect 1046 258 1050 262
rect 1022 238 1026 242
rect 1014 158 1018 162
rect 902 148 906 152
rect 1014 138 1018 142
rect 958 128 962 132
rect 950 118 954 122
rect 926 78 930 82
rect 1014 108 1018 112
rect 1006 98 1010 102
rect 966 78 970 82
rect 718 68 722 72
rect 814 68 818 72
rect 846 68 850 72
rect 878 68 882 72
rect 894 68 898 72
rect 910 68 914 72
rect 782 48 786 52
rect 1206 358 1210 362
rect 1190 348 1194 352
rect 1078 338 1082 342
rect 1118 338 1122 342
rect 1206 338 1210 342
rect 1070 298 1074 302
rect 1070 288 1074 292
rect 1126 318 1130 322
rect 1094 308 1098 312
rect 1206 298 1210 302
rect 1270 698 1274 702
rect 1270 668 1274 672
rect 1342 738 1346 742
rect 1302 728 1306 732
rect 1334 728 1338 732
rect 1286 708 1290 712
rect 1286 688 1290 692
rect 1302 558 1306 562
rect 1270 548 1274 552
rect 1286 548 1290 552
rect 1302 548 1306 552
rect 1302 528 1306 532
rect 1262 518 1266 522
rect 1294 518 1298 522
rect 1350 718 1354 722
rect 1398 708 1402 712
rect 1390 678 1394 682
rect 1374 668 1378 672
rect 1366 648 1370 652
rect 1382 648 1386 652
rect 1354 603 1358 607
rect 1361 603 1365 607
rect 1366 568 1370 572
rect 1342 558 1346 562
rect 1398 578 1402 582
rect 1398 568 1402 572
rect 1374 548 1378 552
rect 1294 508 1298 512
rect 1326 508 1330 512
rect 1342 508 1346 512
rect 1302 498 1306 502
rect 1334 498 1338 502
rect 1270 478 1274 482
rect 1302 468 1306 472
rect 1318 458 1322 462
rect 1334 458 1338 462
rect 1254 398 1258 402
rect 1294 438 1298 442
rect 1318 418 1322 422
rect 1302 388 1306 392
rect 1222 348 1226 352
rect 1214 288 1218 292
rect 1206 278 1210 282
rect 1094 268 1098 272
rect 1174 268 1178 272
rect 1078 258 1082 262
rect 1246 328 1250 332
rect 1358 488 1362 492
rect 1430 708 1434 712
rect 1430 588 1434 592
rect 1430 578 1434 582
rect 1414 468 1418 472
rect 1430 468 1434 472
rect 1406 448 1410 452
rect 1374 428 1378 432
rect 1354 403 1358 407
rect 1361 403 1365 407
rect 1342 398 1346 402
rect 1334 368 1338 372
rect 1350 368 1354 372
rect 1382 368 1386 372
rect 1414 358 1418 362
rect 1310 348 1314 352
rect 1326 348 1330 352
rect 1478 1268 1482 1272
rect 1638 1278 1642 1282
rect 1526 1258 1530 1262
rect 1558 1258 1562 1262
rect 1654 1258 1658 1262
rect 1670 1258 1674 1262
rect 1470 1248 1474 1252
rect 1486 1228 1490 1232
rect 1486 1208 1490 1212
rect 1462 1188 1466 1192
rect 1454 1168 1458 1172
rect 1494 1158 1498 1162
rect 1470 1148 1474 1152
rect 1534 1148 1538 1152
rect 1518 1098 1522 1102
rect 1454 1088 1458 1092
rect 1470 1088 1474 1092
rect 1478 1088 1482 1092
rect 1454 1068 1458 1072
rect 1526 1068 1530 1072
rect 1502 1058 1506 1062
rect 1534 1008 1538 1012
rect 1446 998 1450 1002
rect 1494 968 1498 972
rect 1454 958 1458 962
rect 1446 948 1450 952
rect 1478 938 1482 942
rect 1502 938 1506 942
rect 1486 928 1490 932
rect 1478 908 1482 912
rect 1454 898 1458 902
rect 1454 868 1458 872
rect 1462 868 1466 872
rect 1462 858 1466 862
rect 1462 838 1466 842
rect 1454 748 1458 752
rect 1574 1248 1578 1252
rect 1550 1198 1554 1202
rect 1558 1188 1562 1192
rect 1550 1118 1554 1122
rect 1614 1248 1618 1252
rect 1606 1238 1610 1242
rect 1606 1188 1610 1192
rect 1598 1178 1602 1182
rect 1590 1148 1594 1152
rect 1558 958 1562 962
rect 1606 1148 1610 1152
rect 1630 1148 1634 1152
rect 1630 1118 1634 1122
rect 1606 1068 1610 1072
rect 1718 1298 1722 1302
rect 1710 1278 1714 1282
rect 1790 1478 1794 1482
rect 1774 1468 1778 1472
rect 1798 1468 1802 1472
rect 1734 1448 1738 1452
rect 1782 1438 1786 1442
rect 1822 1458 1826 1462
rect 1774 1388 1778 1392
rect 1822 1388 1826 1392
rect 1798 1358 1802 1362
rect 1782 1348 1786 1352
rect 1758 1308 1762 1312
rect 1734 1278 1738 1282
rect 1686 1258 1690 1262
rect 1726 1248 1730 1252
rect 1726 1238 1730 1242
rect 1766 1258 1770 1262
rect 1694 1178 1698 1182
rect 1654 1158 1658 1162
rect 1678 1148 1682 1152
rect 1766 1148 1770 1152
rect 1654 1128 1658 1132
rect 1686 1078 1690 1082
rect 1614 1058 1618 1062
rect 1630 1058 1634 1062
rect 1646 1058 1650 1062
rect 1614 998 1618 1002
rect 1502 908 1506 912
rect 1542 908 1546 912
rect 1542 888 1546 892
rect 1566 868 1570 872
rect 1590 828 1594 832
rect 1518 818 1522 822
rect 1470 718 1474 722
rect 1606 818 1610 822
rect 1654 1008 1658 1012
rect 1822 1318 1826 1322
rect 1854 1588 1858 1592
rect 1838 1538 1842 1542
rect 1846 1528 1850 1532
rect 1838 1408 1842 1412
rect 1838 1318 1842 1322
rect 1838 1298 1842 1302
rect 2038 1898 2042 1902
rect 2062 1938 2066 1942
rect 2086 1928 2090 1932
rect 2086 1908 2090 1912
rect 2046 1888 2050 1892
rect 2062 1888 2066 1892
rect 2014 1878 2018 1882
rect 2030 1868 2034 1872
rect 2054 1868 2058 1872
rect 2070 1868 2074 1872
rect 1958 1858 1962 1862
rect 1942 1848 1946 1852
rect 1990 1848 1994 1852
rect 2022 1848 2026 1852
rect 2030 1848 2034 1852
rect 1934 1798 1938 1802
rect 2006 1818 2010 1822
rect 2070 1818 2074 1822
rect 2030 1808 2034 1812
rect 1974 1768 1978 1772
rect 2014 1758 2018 1762
rect 1902 1748 1906 1752
rect 1918 1748 1922 1752
rect 1966 1748 1970 1752
rect 1982 1748 1986 1752
rect 1974 1738 1978 1742
rect 1934 1728 1938 1732
rect 1874 1703 1878 1707
rect 1881 1703 1885 1707
rect 1926 1688 1930 1692
rect 1934 1688 1938 1692
rect 1950 1718 1954 1722
rect 1958 1718 1962 1722
rect 1966 1718 1970 1722
rect 1958 1698 1962 1702
rect 1974 1688 1978 1692
rect 1942 1678 1946 1682
rect 1902 1658 1906 1662
rect 1942 1658 1946 1662
rect 1894 1648 1898 1652
rect 1934 1648 1938 1652
rect 1894 1598 1898 1602
rect 1902 1588 1906 1592
rect 1958 1628 1962 1632
rect 1950 1608 1954 1612
rect 1942 1578 1946 1582
rect 1918 1568 1922 1572
rect 1966 1558 1970 1562
rect 2014 1728 2018 1732
rect 2006 1648 2010 1652
rect 1990 1638 1994 1642
rect 2006 1608 2010 1612
rect 2046 1798 2050 1802
rect 2054 1768 2058 1772
rect 2062 1758 2066 1762
rect 2038 1728 2042 1732
rect 2038 1708 2042 1712
rect 2062 1728 2066 1732
rect 2046 1698 2050 1702
rect 2038 1678 2042 1682
rect 2046 1678 2050 1682
rect 2150 2148 2154 2152
rect 2150 2078 2154 2082
rect 2222 2368 2226 2372
rect 2222 2358 2226 2362
rect 2254 2478 2258 2482
rect 2318 2648 2322 2652
rect 2486 3248 2490 3252
rect 2446 3208 2450 3212
rect 2430 3148 2434 3152
rect 2422 3068 2426 3072
rect 2454 3058 2458 3062
rect 2366 3048 2370 3052
rect 2374 3048 2378 3052
rect 2386 3003 2390 3007
rect 2393 3003 2397 3007
rect 2438 3048 2442 3052
rect 2446 3048 2450 3052
rect 2454 2988 2458 2992
rect 2430 2948 2434 2952
rect 2446 2948 2450 2952
rect 2390 2918 2394 2922
rect 2430 2868 2434 2872
rect 2366 2858 2370 2862
rect 2422 2858 2426 2862
rect 2366 2848 2370 2852
rect 2386 2803 2390 2807
rect 2393 2803 2397 2807
rect 2406 2798 2410 2802
rect 2382 2768 2386 2772
rect 2358 2698 2362 2702
rect 2422 2648 2426 2652
rect 2326 2638 2330 2642
rect 2358 2638 2362 2642
rect 2342 2628 2346 2632
rect 2310 2618 2314 2622
rect 2302 2538 2306 2542
rect 2286 2508 2290 2512
rect 2302 2498 2306 2502
rect 2238 2458 2242 2462
rect 2246 2448 2250 2452
rect 2238 2438 2242 2442
rect 2286 2448 2290 2452
rect 2270 2438 2274 2442
rect 2334 2598 2338 2602
rect 2386 2603 2390 2607
rect 2393 2603 2397 2607
rect 2470 3198 2474 3202
rect 2494 3158 2498 3162
rect 2486 3148 2490 3152
rect 2526 3248 2530 3252
rect 2534 3228 2538 3232
rect 2526 3208 2530 3212
rect 2510 3198 2514 3202
rect 2510 3178 2514 3182
rect 2518 3158 2522 3162
rect 2478 3138 2482 3142
rect 2510 3138 2514 3142
rect 2486 3128 2490 3132
rect 2558 3328 2562 3332
rect 2566 3298 2570 3302
rect 2646 3488 2650 3492
rect 2638 3478 2642 3482
rect 2638 3458 2642 3462
rect 2622 3428 2626 3432
rect 2622 3378 2626 3382
rect 2630 3358 2634 3362
rect 2614 3348 2618 3352
rect 2598 3318 2602 3322
rect 2614 3308 2618 3312
rect 2638 3338 2642 3342
rect 2638 3318 2642 3322
rect 2638 3298 2642 3302
rect 2678 3538 2682 3542
rect 2686 3478 2690 3482
rect 2678 3468 2682 3472
rect 2702 3458 2706 3462
rect 2782 3738 2786 3742
rect 2798 3738 2802 3742
rect 2790 3728 2794 3732
rect 2830 3748 2834 3752
rect 2890 3903 2894 3907
rect 2897 3903 2901 3907
rect 3054 3928 3058 3932
rect 2926 3908 2930 3912
rect 2974 3898 2978 3902
rect 2974 3888 2978 3892
rect 2878 3878 2882 3882
rect 2918 3878 2922 3882
rect 2910 3868 2914 3872
rect 2918 3858 2922 3862
rect 2974 3858 2978 3862
rect 2862 3848 2866 3852
rect 2926 3838 2930 3842
rect 2838 3738 2842 3742
rect 2814 3718 2818 3722
rect 2878 3728 2882 3732
rect 2862 3718 2866 3722
rect 2742 3698 2746 3702
rect 2846 3698 2850 3702
rect 2806 3688 2810 3692
rect 2790 3678 2794 3682
rect 2814 3678 2818 3682
rect 2838 3678 2842 3682
rect 2734 3668 2738 3672
rect 2726 3608 2730 3612
rect 2766 3648 2770 3652
rect 2774 3648 2778 3652
rect 2750 3638 2754 3642
rect 2890 3703 2894 3707
rect 2897 3703 2901 3707
rect 2846 3658 2850 3662
rect 2798 3648 2802 3652
rect 2782 3628 2786 3632
rect 2766 3608 2770 3612
rect 2742 3588 2746 3592
rect 2790 3578 2794 3582
rect 2742 3548 2746 3552
rect 2846 3648 2850 3652
rect 2854 3648 2858 3652
rect 2814 3608 2818 3612
rect 2878 3648 2882 3652
rect 2902 3648 2906 3652
rect 2862 3598 2866 3602
rect 2870 3598 2874 3602
rect 2830 3578 2834 3582
rect 2814 3568 2818 3572
rect 2846 3568 2850 3572
rect 2878 3578 2882 3582
rect 2830 3558 2834 3562
rect 2862 3558 2866 3562
rect 2822 3548 2826 3552
rect 2774 3528 2778 3532
rect 2790 3498 2794 3502
rect 2750 3488 2754 3492
rect 2670 3438 2674 3442
rect 2814 3538 2818 3542
rect 2902 3547 2906 3551
rect 2878 3538 2882 3542
rect 2854 3528 2858 3532
rect 2870 3518 2874 3522
rect 2830 3508 2834 3512
rect 2862 3508 2866 3512
rect 2814 3478 2818 3482
rect 2838 3478 2842 3482
rect 2798 3468 2802 3472
rect 3126 3908 3130 3912
rect 3094 3878 3098 3882
rect 3118 3878 3122 3882
rect 3126 3868 3130 3872
rect 3046 3858 3050 3862
rect 3070 3858 3074 3862
rect 3134 3858 3138 3862
rect 3150 3858 3154 3862
rect 3038 3838 3042 3842
rect 3086 3808 3090 3812
rect 2982 3788 2986 3792
rect 3086 3788 3090 3792
rect 3046 3768 3050 3772
rect 3022 3758 3026 3762
rect 3030 3758 3034 3762
rect 3046 3758 3050 3762
rect 2918 3748 2922 3752
rect 2950 3748 2954 3752
rect 2982 3748 2986 3752
rect 3006 3748 3010 3752
rect 2974 3728 2978 3732
rect 2966 3708 2970 3712
rect 2974 3708 2978 3712
rect 2918 3698 2922 3702
rect 2998 3728 3002 3732
rect 2982 3698 2986 3702
rect 2966 3688 2970 3692
rect 2974 3688 2978 3692
rect 2990 3678 2994 3682
rect 2966 3668 2970 3672
rect 3022 3678 3026 3682
rect 3014 3668 3018 3672
rect 2934 3658 2938 3662
rect 2942 3658 2946 3662
rect 2958 3658 2962 3662
rect 2982 3658 2986 3662
rect 2950 3648 2954 3652
rect 2974 3648 2978 3652
rect 2926 3638 2930 3642
rect 2918 3628 2922 3632
rect 3110 3708 3114 3712
rect 3038 3688 3042 3692
rect 3086 3688 3090 3692
rect 3102 3688 3106 3692
rect 3198 3918 3202 3922
rect 3214 3918 3218 3922
rect 3214 3878 3218 3882
rect 3222 3858 3226 3862
rect 3182 3848 3186 3852
rect 3182 3828 3186 3832
rect 3150 3758 3154 3762
rect 3158 3728 3162 3732
rect 3206 3788 3210 3792
rect 3174 3748 3178 3752
rect 3278 4128 3282 4132
rect 3270 4088 3274 4092
rect 3278 4088 3282 4092
rect 3302 4198 3306 4202
rect 3318 4178 3322 4182
rect 3310 4098 3314 4102
rect 3302 4078 3306 4082
rect 3262 4058 3266 4062
rect 3254 4048 3258 4052
rect 3246 4038 3250 4042
rect 3310 4038 3314 4042
rect 3302 3998 3306 4002
rect 3286 3968 3290 3972
rect 3550 4998 3554 5002
rect 3654 5008 3658 5012
rect 3542 4978 3546 4982
rect 3558 4978 3562 4982
rect 3630 4978 3634 4982
rect 3534 4968 3538 4972
rect 3558 4968 3562 4972
rect 3510 4958 3514 4962
rect 3542 4958 3546 4962
rect 3486 4947 3490 4951
rect 3502 4878 3506 4882
rect 3662 4968 3666 4972
rect 3654 4958 3658 4962
rect 3550 4948 3554 4952
rect 3614 4948 3618 4952
rect 3654 4948 3658 4952
rect 3574 4938 3578 4942
rect 3590 4938 3594 4942
rect 3566 4918 3570 4922
rect 3582 4918 3586 4922
rect 3550 4878 3554 4882
rect 3622 4918 3626 4922
rect 3598 4888 3602 4892
rect 3614 4888 3618 4892
rect 3550 4868 3554 4872
rect 3478 4838 3482 4842
rect 3502 4838 3506 4842
rect 3526 4798 3530 4802
rect 3494 4748 3498 4752
rect 3542 4748 3546 4752
rect 3446 4738 3450 4742
rect 3462 4678 3466 4682
rect 3438 4668 3442 4672
rect 3502 4708 3506 4712
rect 3486 4698 3490 4702
rect 3462 4648 3466 4652
rect 3486 4648 3490 4652
rect 3494 4648 3498 4652
rect 3454 4548 3458 4552
rect 3446 4538 3450 4542
rect 3502 4618 3506 4622
rect 3494 4578 3498 4582
rect 3478 4558 3482 4562
rect 3462 4528 3466 4532
rect 3622 4878 3626 4882
rect 3654 4918 3658 4922
rect 3710 5048 3714 5052
rect 3726 5048 3730 5052
rect 3694 5038 3698 5042
rect 3702 5038 3706 5042
rect 3718 5038 3722 5042
rect 3702 4998 3706 5002
rect 3734 5018 3738 5022
rect 3766 5008 3770 5012
rect 3694 4948 3698 4952
rect 3678 4938 3682 4942
rect 3686 4938 3690 4942
rect 3694 4938 3698 4942
rect 3670 4878 3674 4882
rect 3702 4928 3706 4932
rect 3726 4938 3730 4942
rect 3574 4848 3578 4852
rect 3598 4848 3602 4852
rect 3606 4838 3610 4842
rect 3614 4838 3618 4842
rect 3582 4798 3586 4802
rect 3630 4858 3634 4862
rect 3622 4808 3626 4812
rect 3566 4728 3570 4732
rect 3550 4708 3554 4712
rect 3574 4708 3578 4712
rect 3566 4678 3570 4682
rect 3590 4678 3594 4682
rect 3654 4838 3658 4842
rect 3678 4858 3682 4862
rect 3686 4858 3690 4862
rect 3670 4838 3674 4842
rect 3662 4808 3666 4812
rect 3678 4808 3682 4812
rect 3638 4758 3642 4762
rect 3662 4748 3666 4752
rect 3718 4848 3722 4852
rect 3702 4768 3706 4772
rect 3838 5048 3842 5052
rect 4014 5028 4018 5032
rect 3998 5018 4002 5022
rect 3838 4998 3842 5002
rect 3798 4988 3802 4992
rect 3846 4988 3850 4992
rect 3790 4958 3794 4962
rect 3782 4948 3786 4952
rect 3758 4918 3762 4922
rect 3758 4888 3762 4892
rect 3734 4878 3738 4882
rect 3742 4848 3746 4852
rect 3750 4828 3754 4832
rect 3734 4788 3738 4792
rect 3750 4778 3754 4782
rect 3678 4708 3682 4712
rect 3638 4678 3642 4682
rect 3678 4668 3682 4672
rect 3630 4658 3634 4662
rect 3534 4548 3538 4552
rect 3510 4538 3514 4542
rect 3526 4538 3530 4542
rect 3454 4518 3458 4522
rect 3494 4518 3498 4522
rect 3438 4468 3442 4472
rect 3446 4378 3450 4382
rect 3438 4358 3442 4362
rect 3422 4328 3426 4332
rect 3446 4348 3450 4352
rect 3390 4318 3394 4322
rect 3390 4258 3394 4262
rect 3462 4448 3466 4452
rect 3334 4138 3338 4142
rect 3358 4138 3362 4142
rect 3326 4128 3330 4132
rect 3350 4078 3354 4082
rect 3334 4028 3338 4032
rect 3326 3978 3330 3982
rect 3318 3948 3322 3952
rect 3286 3928 3290 3932
rect 3262 3898 3266 3902
rect 3318 3918 3322 3922
rect 3318 3898 3322 3902
rect 3278 3878 3282 3882
rect 3310 3858 3314 3862
rect 3294 3838 3298 3842
rect 3278 3808 3282 3812
rect 3262 3778 3266 3782
rect 3222 3748 3226 3752
rect 3230 3748 3234 3752
rect 3182 3728 3186 3732
rect 3270 3728 3274 3732
rect 3198 3718 3202 3722
rect 3254 3698 3258 3702
rect 3030 3668 3034 3672
rect 3046 3668 3050 3672
rect 3118 3668 3122 3672
rect 3166 3668 3170 3672
rect 3246 3668 3250 3672
rect 3270 3668 3274 3672
rect 3038 3658 3042 3662
rect 3086 3658 3090 3662
rect 3158 3658 3162 3662
rect 3054 3638 3058 3642
rect 3054 3588 3058 3592
rect 2966 3568 2970 3572
rect 3030 3568 3034 3572
rect 3054 3568 3058 3572
rect 2974 3558 2978 3562
rect 2998 3558 3002 3562
rect 3022 3548 3026 3552
rect 3046 3548 3050 3552
rect 2910 3508 2914 3512
rect 2890 3503 2894 3507
rect 2897 3503 2901 3507
rect 2750 3448 2754 3452
rect 2822 3448 2826 3452
rect 2750 3438 2754 3442
rect 2814 3438 2818 3442
rect 2846 3438 2850 3442
rect 2886 3438 2890 3442
rect 2726 3418 2730 3422
rect 2678 3398 2682 3402
rect 2710 3408 2714 3412
rect 2694 3378 2698 3382
rect 2694 3368 2698 3372
rect 2670 3358 2674 3362
rect 2742 3358 2746 3362
rect 2782 3418 2786 3422
rect 2662 3348 2666 3352
rect 2702 3348 2706 3352
rect 2726 3348 2730 3352
rect 2758 3348 2762 3352
rect 2806 3378 2810 3382
rect 2798 3358 2802 3362
rect 2654 3338 2658 3342
rect 2766 3338 2770 3342
rect 2662 3308 2666 3312
rect 2670 3288 2674 3292
rect 2678 3288 2682 3292
rect 2710 3318 2714 3322
rect 2790 3308 2794 3312
rect 2742 3298 2746 3302
rect 2678 3268 2682 3272
rect 2686 3268 2690 3272
rect 2726 3268 2730 3272
rect 2646 3228 2650 3232
rect 2606 3198 2610 3202
rect 2574 3178 2578 3182
rect 2550 3158 2554 3162
rect 2614 3158 2618 3162
rect 2566 3148 2570 3152
rect 2638 3168 2642 3172
rect 2654 3168 2658 3172
rect 2670 3218 2674 3222
rect 2670 3168 2674 3172
rect 2654 3138 2658 3142
rect 2534 3128 2538 3132
rect 2550 3118 2554 3122
rect 2478 3088 2482 3092
rect 2494 3088 2498 3092
rect 2566 3098 2570 3102
rect 2598 3098 2602 3102
rect 2662 3118 2666 3122
rect 2630 3088 2634 3092
rect 2958 3538 2962 3542
rect 2998 3518 3002 3522
rect 3118 3547 3122 3551
rect 3238 3658 3242 3662
rect 3206 3648 3210 3652
rect 3214 3648 3218 3652
rect 3190 3638 3194 3642
rect 3222 3608 3226 3612
rect 3246 3598 3250 3602
rect 3158 3588 3162 3592
rect 3174 3578 3178 3582
rect 3190 3568 3194 3572
rect 3182 3548 3186 3552
rect 3246 3548 3250 3552
rect 3038 3538 3042 3542
rect 2950 3488 2954 3492
rect 2974 3478 2978 3482
rect 3078 3478 3082 3482
rect 2966 3468 2970 3472
rect 2990 3468 2994 3472
rect 3006 3468 3010 3472
rect 3190 3538 3194 3542
rect 3158 3518 3162 3522
rect 3206 3518 3210 3522
rect 3254 3528 3258 3532
rect 3222 3518 3226 3522
rect 3214 3498 3218 3502
rect 3206 3488 3210 3492
rect 3174 3468 3178 3472
rect 3006 3458 3010 3462
rect 2950 3448 2954 3452
rect 2950 3418 2954 3422
rect 2926 3408 2930 3412
rect 2902 3348 2906 3352
rect 2862 3338 2866 3342
rect 2902 3338 2906 3342
rect 2974 3408 2978 3412
rect 2990 3328 2994 3332
rect 2966 3318 2970 3322
rect 2890 3303 2894 3307
rect 2897 3303 2901 3307
rect 2814 3298 2818 3302
rect 2870 3298 2874 3302
rect 2926 3298 2930 3302
rect 2966 3298 2970 3302
rect 2838 3288 2842 3292
rect 2870 3288 2874 3292
rect 2950 3288 2954 3292
rect 2958 3288 2962 3292
rect 2990 3278 2994 3282
rect 2702 3258 2706 3262
rect 2758 3258 2762 3262
rect 2886 3258 2890 3262
rect 2934 3258 2938 3262
rect 2942 3258 2946 3262
rect 2990 3258 2994 3262
rect 2718 3238 2722 3242
rect 2758 3248 2762 3252
rect 2750 3228 2754 3232
rect 2838 3248 2842 3252
rect 2806 3238 2810 3242
rect 2766 3198 2770 3202
rect 2726 3178 2730 3182
rect 2782 3178 2786 3182
rect 2686 3168 2690 3172
rect 2790 3158 2794 3162
rect 2790 3148 2794 3152
rect 2726 3128 2730 3132
rect 2702 3088 2706 3092
rect 2558 3078 2562 3082
rect 2678 3078 2682 3082
rect 2470 3068 2474 3072
rect 2598 3068 2602 3072
rect 2606 3068 2610 3072
rect 2630 3068 2634 3072
rect 2518 3058 2522 3062
rect 2558 3058 2562 3062
rect 2590 3058 2594 3062
rect 2614 3058 2618 3062
rect 2638 3058 2642 3062
rect 2470 3018 2474 3022
rect 2470 2998 2474 3002
rect 2534 3048 2538 3052
rect 2582 3048 2586 3052
rect 2630 3048 2634 3052
rect 2478 2968 2482 2972
rect 2502 2968 2506 2972
rect 2510 2948 2514 2952
rect 2486 2938 2490 2942
rect 2566 3008 2570 3012
rect 2566 2988 2570 2992
rect 2550 2978 2554 2982
rect 2686 2968 2690 2972
rect 2574 2958 2578 2962
rect 2646 2958 2650 2962
rect 2670 2958 2674 2962
rect 2622 2948 2626 2952
rect 2510 2918 2514 2922
rect 2478 2888 2482 2892
rect 2462 2818 2466 2822
rect 2462 2808 2466 2812
rect 2446 2738 2450 2742
rect 2510 2868 2514 2872
rect 2566 2938 2570 2942
rect 2550 2928 2554 2932
rect 2614 2938 2618 2942
rect 2654 2938 2658 2942
rect 2582 2918 2586 2922
rect 2534 2908 2538 2912
rect 2598 2898 2602 2902
rect 2574 2888 2578 2892
rect 2598 2888 2602 2892
rect 2526 2878 2530 2882
rect 2558 2878 2562 2882
rect 2518 2848 2522 2852
rect 2486 2798 2490 2802
rect 2486 2768 2490 2772
rect 2502 2768 2506 2772
rect 2782 3118 2786 3122
rect 2790 3108 2794 3112
rect 2758 3078 2762 3082
rect 2718 3048 2722 3052
rect 2782 3058 2786 3062
rect 2782 3048 2786 3052
rect 2854 3218 2858 3222
rect 2830 3208 2834 3212
rect 2814 3158 2818 3162
rect 2902 3238 2906 3242
rect 2910 3218 2914 3222
rect 2894 3188 2898 3192
rect 2838 3168 2842 3172
rect 2854 3158 2858 3162
rect 2846 3138 2850 3142
rect 2838 3128 2842 3132
rect 2902 3128 2906 3132
rect 2890 3103 2894 3107
rect 2897 3103 2901 3107
rect 2878 3098 2882 3102
rect 2878 3088 2882 3092
rect 2846 3078 2850 3082
rect 2838 3058 2842 3062
rect 2862 3058 2866 3062
rect 2886 3058 2890 3062
rect 2830 3048 2834 3052
rect 2774 3038 2778 3042
rect 2862 3038 2866 3042
rect 2830 3018 2834 3022
rect 2766 2968 2770 2972
rect 2814 2968 2818 2972
rect 2710 2958 2714 2962
rect 2702 2948 2706 2952
rect 2702 2938 2706 2942
rect 2758 2938 2762 2942
rect 2638 2908 2642 2912
rect 2678 2908 2682 2912
rect 2630 2898 2634 2902
rect 2622 2888 2626 2892
rect 2638 2878 2642 2882
rect 2542 2868 2546 2872
rect 2590 2868 2594 2872
rect 2622 2868 2626 2872
rect 2614 2858 2618 2862
rect 2662 2859 2666 2863
rect 2670 2828 2674 2832
rect 2526 2818 2530 2822
rect 2654 2778 2658 2782
rect 2558 2768 2562 2772
rect 2494 2758 2498 2762
rect 2534 2758 2538 2762
rect 2606 2758 2610 2762
rect 2510 2748 2514 2752
rect 2550 2748 2554 2752
rect 2638 2748 2642 2752
rect 2478 2718 2482 2722
rect 2510 2718 2514 2722
rect 2446 2638 2450 2642
rect 2478 2698 2482 2702
rect 2470 2648 2474 2652
rect 2518 2648 2522 2652
rect 2502 2638 2506 2642
rect 2462 2608 2466 2612
rect 2486 2608 2490 2612
rect 2398 2558 2402 2562
rect 2446 2558 2450 2562
rect 2382 2518 2386 2522
rect 2374 2478 2378 2482
rect 2350 2458 2354 2462
rect 2246 2388 2250 2392
rect 2254 2368 2258 2372
rect 2238 2358 2242 2362
rect 2262 2358 2266 2362
rect 2294 2358 2298 2362
rect 2246 2348 2250 2352
rect 2238 2338 2242 2342
rect 2230 2308 2234 2312
rect 2222 2268 2226 2272
rect 2246 2268 2250 2272
rect 2278 2338 2282 2342
rect 2294 2338 2298 2342
rect 2270 2298 2274 2302
rect 2326 2438 2330 2442
rect 2342 2398 2346 2402
rect 2286 2318 2290 2322
rect 2318 2318 2322 2322
rect 2334 2328 2338 2332
rect 2334 2298 2338 2302
rect 2278 2268 2282 2272
rect 2334 2268 2338 2272
rect 2246 2238 2250 2242
rect 2214 2218 2218 2222
rect 2238 2198 2242 2202
rect 2198 2158 2202 2162
rect 2422 2498 2426 2502
rect 2414 2448 2418 2452
rect 2374 2438 2378 2442
rect 2382 2438 2386 2442
rect 2430 2438 2434 2442
rect 2386 2403 2390 2407
rect 2393 2403 2397 2407
rect 2470 2468 2474 2472
rect 2478 2468 2482 2472
rect 2454 2458 2458 2462
rect 2462 2448 2466 2452
rect 2438 2408 2442 2412
rect 2374 2388 2378 2392
rect 2358 2378 2362 2382
rect 2358 2298 2362 2302
rect 2302 2258 2306 2262
rect 2310 2258 2314 2262
rect 2278 2198 2282 2202
rect 2262 2168 2266 2172
rect 2254 2158 2258 2162
rect 2182 2148 2186 2152
rect 2230 2148 2234 2152
rect 2278 2148 2282 2152
rect 2302 2208 2306 2212
rect 2310 2188 2314 2192
rect 2302 2158 2306 2162
rect 2358 2198 2362 2202
rect 2318 2168 2322 2172
rect 2318 2148 2322 2152
rect 2214 2098 2218 2102
rect 2166 2068 2170 2072
rect 2102 2058 2106 2062
rect 2134 2058 2138 2062
rect 2150 2058 2154 2062
rect 2110 2048 2114 2052
rect 2110 2028 2114 2032
rect 2126 2048 2130 2052
rect 2142 2038 2146 2042
rect 2134 1998 2138 2002
rect 2118 1988 2122 1992
rect 2102 1968 2106 1972
rect 2126 1968 2130 1972
rect 2110 1948 2114 1952
rect 2118 1938 2122 1942
rect 2166 2048 2170 2052
rect 2126 1928 2130 1932
rect 2142 1928 2146 1932
rect 2158 1918 2162 1922
rect 2166 1898 2170 1902
rect 2254 2138 2258 2142
rect 2262 2138 2266 2142
rect 2302 2138 2306 2142
rect 2270 2128 2274 2132
rect 2254 2108 2258 2112
rect 2238 2088 2242 2092
rect 2246 2078 2250 2082
rect 2230 2048 2234 2052
rect 2294 2118 2298 2122
rect 2310 2108 2314 2112
rect 2350 2138 2354 2142
rect 2414 2368 2418 2372
rect 2422 2358 2426 2362
rect 2430 2358 2434 2362
rect 2398 2348 2402 2352
rect 2374 2338 2378 2342
rect 2374 2308 2378 2312
rect 2374 2258 2378 2262
rect 2406 2248 2410 2252
rect 2382 2238 2386 2242
rect 2414 2228 2418 2232
rect 2374 2208 2378 2212
rect 2386 2203 2390 2207
rect 2393 2203 2397 2207
rect 2414 2098 2418 2102
rect 2446 2388 2450 2392
rect 2454 2328 2458 2332
rect 2430 2268 2434 2272
rect 2446 2268 2450 2272
rect 2438 2168 2442 2172
rect 2446 2148 2450 2152
rect 2438 2118 2442 2122
rect 2430 2108 2434 2112
rect 2438 2108 2442 2112
rect 2366 2078 2370 2082
rect 2422 2078 2426 2082
rect 2294 2068 2298 2072
rect 2326 2068 2330 2072
rect 2358 2068 2362 2072
rect 2262 2018 2266 2022
rect 2230 1968 2234 1972
rect 2246 1968 2250 1972
rect 2230 1938 2234 1942
rect 2262 1918 2266 1922
rect 2222 1898 2226 1902
rect 2174 1878 2178 1882
rect 2446 2078 2450 2082
rect 2294 2048 2298 2052
rect 2390 2028 2394 2032
rect 2318 2018 2322 2022
rect 2374 2008 2378 2012
rect 2386 2003 2390 2007
rect 2393 2003 2397 2007
rect 2342 1988 2346 1992
rect 2430 1988 2434 1992
rect 2294 1958 2298 1962
rect 2366 1948 2370 1952
rect 2414 1948 2418 1952
rect 2334 1928 2338 1932
rect 2358 1928 2362 1932
rect 2270 1888 2274 1892
rect 2334 1888 2338 1892
rect 2342 1888 2346 1892
rect 2230 1878 2234 1882
rect 2270 1878 2274 1882
rect 2118 1868 2122 1872
rect 2238 1868 2242 1872
rect 2094 1798 2098 1802
rect 2102 1778 2106 1782
rect 2190 1858 2194 1862
rect 2158 1778 2162 1782
rect 2166 1768 2170 1772
rect 2102 1698 2106 1702
rect 2086 1688 2090 1692
rect 2094 1688 2098 1692
rect 2022 1588 2026 1592
rect 1982 1578 1986 1582
rect 1926 1538 1930 1542
rect 1974 1538 1978 1542
rect 1862 1528 1866 1532
rect 1874 1503 1878 1507
rect 1881 1503 1885 1507
rect 1862 1498 1866 1502
rect 1918 1498 1922 1502
rect 1854 1478 1858 1482
rect 1966 1528 1970 1532
rect 1942 1508 1946 1512
rect 1958 1508 1962 1512
rect 1966 1488 1970 1492
rect 1894 1458 1898 1462
rect 1902 1458 1906 1462
rect 1918 1458 1922 1462
rect 1854 1438 1858 1442
rect 1838 1268 1842 1272
rect 1822 1258 1826 1262
rect 1838 1258 1842 1262
rect 1894 1398 1898 1402
rect 1862 1358 1866 1362
rect 1878 1348 1882 1352
rect 1874 1303 1878 1307
rect 1881 1303 1885 1307
rect 1862 1288 1866 1292
rect 1822 1168 1826 1172
rect 1846 1148 1850 1152
rect 1782 1118 1786 1122
rect 1822 1118 1826 1122
rect 1758 1108 1762 1112
rect 1742 1098 1746 1102
rect 1758 1098 1762 1102
rect 1798 1088 1802 1092
rect 1838 1098 1842 1102
rect 1718 1068 1722 1072
rect 1734 1068 1738 1072
rect 1734 1058 1738 1062
rect 1750 1058 1754 1062
rect 1806 1058 1810 1062
rect 1710 1038 1714 1042
rect 1670 958 1674 962
rect 1686 958 1690 962
rect 1654 948 1658 952
rect 1678 938 1682 942
rect 1638 918 1642 922
rect 1686 898 1690 902
rect 1774 978 1778 982
rect 1710 948 1714 952
rect 1742 948 1746 952
rect 1726 938 1730 942
rect 1686 878 1690 882
rect 1694 878 1698 882
rect 1654 868 1658 872
rect 1622 858 1626 862
rect 1646 858 1650 862
rect 1718 918 1722 922
rect 1726 908 1730 912
rect 1710 868 1714 872
rect 1694 858 1698 862
rect 1702 858 1706 862
rect 1734 858 1738 862
rect 1630 848 1634 852
rect 1670 848 1674 852
rect 1622 808 1626 812
rect 1614 798 1618 802
rect 1718 848 1722 852
rect 1742 848 1746 852
rect 1766 918 1770 922
rect 1758 888 1762 892
rect 1758 858 1762 862
rect 1750 838 1754 842
rect 1678 788 1682 792
rect 1694 768 1698 772
rect 1766 808 1770 812
rect 1766 788 1770 792
rect 1750 758 1754 762
rect 1526 748 1530 752
rect 1630 748 1634 752
rect 1662 748 1666 752
rect 1542 738 1546 742
rect 1518 718 1522 722
rect 1502 708 1506 712
rect 1542 688 1546 692
rect 1710 738 1714 742
rect 1606 728 1610 732
rect 1670 718 1674 722
rect 1718 718 1722 722
rect 1638 708 1642 712
rect 1614 688 1618 692
rect 1574 678 1578 682
rect 1454 658 1458 662
rect 1486 658 1490 662
rect 1678 688 1682 692
rect 1686 688 1690 692
rect 1614 668 1618 672
rect 1654 668 1658 672
rect 1566 658 1570 662
rect 1510 638 1514 642
rect 1510 628 1514 632
rect 1470 598 1474 602
rect 1486 588 1490 592
rect 1718 668 1722 672
rect 1646 658 1650 662
rect 1678 658 1682 662
rect 1622 648 1626 652
rect 1598 638 1602 642
rect 1574 608 1578 612
rect 1574 558 1578 562
rect 1502 528 1506 532
rect 1462 488 1466 492
rect 1486 478 1490 482
rect 1558 548 1562 552
rect 1550 538 1554 542
rect 1566 528 1570 532
rect 1574 488 1578 492
rect 1590 568 1594 572
rect 1750 748 1754 752
rect 1742 738 1746 742
rect 1758 738 1762 742
rect 1806 938 1810 942
rect 1806 918 1810 922
rect 1782 858 1786 862
rect 1782 808 1786 812
rect 1790 778 1794 782
rect 1782 728 1786 732
rect 1774 678 1778 682
rect 1822 868 1826 872
rect 1830 858 1834 862
rect 1806 848 1810 852
rect 1822 768 1826 772
rect 1934 1468 1938 1472
rect 1950 1468 1954 1472
rect 1974 1468 1978 1472
rect 1998 1558 2002 1562
rect 2030 1558 2034 1562
rect 2038 1548 2042 1552
rect 2006 1538 2010 1542
rect 2030 1538 2034 1542
rect 2046 1538 2050 1542
rect 1998 1528 2002 1532
rect 2038 1528 2042 1532
rect 2014 1468 2018 1472
rect 1990 1458 1994 1462
rect 1982 1418 1986 1422
rect 1958 1408 1962 1412
rect 1974 1408 1978 1412
rect 1958 1358 1962 1362
rect 1958 1348 1962 1352
rect 1942 1278 1946 1282
rect 1934 1248 1938 1252
rect 1966 1328 1970 1332
rect 1982 1298 1986 1302
rect 1974 1288 1978 1292
rect 1982 1278 1986 1282
rect 2022 1448 2026 1452
rect 2014 1438 2018 1442
rect 2046 1518 2050 1522
rect 2054 1498 2058 1502
rect 2142 1738 2146 1742
rect 2158 1728 2162 1732
rect 2174 1718 2178 1722
rect 2206 1848 2210 1852
rect 2190 1838 2194 1842
rect 2182 1688 2186 1692
rect 2118 1668 2122 1672
rect 2126 1668 2130 1672
rect 2110 1658 2114 1662
rect 2070 1648 2074 1652
rect 2086 1648 2090 1652
rect 2118 1638 2122 1642
rect 2110 1588 2114 1592
rect 2166 1588 2170 1592
rect 2134 1548 2138 1552
rect 2174 1548 2178 1552
rect 2142 1528 2146 1532
rect 2086 1518 2090 1522
rect 2134 1518 2138 1522
rect 2062 1468 2066 1472
rect 2054 1458 2058 1462
rect 2150 1508 2154 1512
rect 2126 1488 2130 1492
rect 2118 1468 2122 1472
rect 2150 1458 2154 1462
rect 2078 1438 2082 1442
rect 2102 1438 2106 1442
rect 2014 1368 2018 1372
rect 2094 1368 2098 1372
rect 2014 1348 2018 1352
rect 2038 1348 2042 1352
rect 2046 1348 2050 1352
rect 2022 1338 2026 1342
rect 1998 1318 2002 1322
rect 2014 1308 2018 1312
rect 2014 1288 2018 1292
rect 2030 1328 2034 1332
rect 2014 1258 2018 1262
rect 1958 1238 1962 1242
rect 1982 1208 1986 1212
rect 1894 1198 1898 1202
rect 1950 1198 1954 1202
rect 1878 1148 1882 1152
rect 1894 1108 1898 1112
rect 1874 1103 1878 1107
rect 1881 1103 1885 1107
rect 1934 1118 1938 1122
rect 2022 1248 2026 1252
rect 2006 1238 2010 1242
rect 2022 1228 2026 1232
rect 2126 1448 2130 1452
rect 2110 1308 2114 1312
rect 2038 1258 2042 1262
rect 2070 1248 2074 1252
rect 2070 1188 2074 1192
rect 2030 1178 2034 1182
rect 2046 1148 2050 1152
rect 2062 1148 2066 1152
rect 2014 1138 2018 1142
rect 2038 1118 2042 1122
rect 2006 1088 2010 1092
rect 2046 1098 2050 1102
rect 1958 1068 1962 1072
rect 1990 1068 1994 1072
rect 1998 1068 2002 1072
rect 1854 1058 1858 1062
rect 1910 1058 1914 1062
rect 1942 1058 1946 1062
rect 1966 1058 1970 1062
rect 1990 1058 1994 1062
rect 1886 1048 1890 1052
rect 1982 1038 1986 1042
rect 1902 978 1906 982
rect 1966 968 1970 972
rect 1966 958 1970 962
rect 2038 1048 2042 1052
rect 2030 1008 2034 1012
rect 1998 988 2002 992
rect 2102 1248 2106 1252
rect 2102 1218 2106 1222
rect 2086 1168 2090 1172
rect 2094 1158 2098 1162
rect 2142 1358 2146 1362
rect 2182 1518 2186 1522
rect 2174 1478 2178 1482
rect 2158 1418 2162 1422
rect 2230 1818 2234 1822
rect 2222 1798 2226 1802
rect 2206 1768 2210 1772
rect 2214 1728 2218 1732
rect 2230 1668 2234 1672
rect 2270 1828 2274 1832
rect 2334 1858 2338 1862
rect 2326 1828 2330 1832
rect 2310 1818 2314 1822
rect 2318 1818 2322 1822
rect 2286 1808 2290 1812
rect 2262 1708 2266 1712
rect 2254 1658 2258 1662
rect 2214 1628 2218 1632
rect 2246 1598 2250 1602
rect 2230 1588 2234 1592
rect 2230 1558 2234 1562
rect 2222 1478 2226 1482
rect 2214 1468 2218 1472
rect 2422 1908 2426 1912
rect 2414 1898 2418 1902
rect 2406 1888 2410 1892
rect 2462 2268 2466 2272
rect 2494 2538 2498 2542
rect 2510 2508 2514 2512
rect 2502 2358 2506 2362
rect 2486 2328 2490 2332
rect 2518 2328 2522 2332
rect 2494 2308 2498 2312
rect 2542 2718 2546 2722
rect 2574 2718 2578 2722
rect 2582 2718 2586 2722
rect 2606 2738 2610 2742
rect 2630 2738 2634 2742
rect 2598 2728 2602 2732
rect 2622 2728 2626 2732
rect 2598 2718 2602 2722
rect 2590 2708 2594 2712
rect 2550 2698 2554 2702
rect 2558 2698 2562 2702
rect 2582 2698 2586 2702
rect 2566 2608 2570 2612
rect 2574 2558 2578 2562
rect 2558 2548 2562 2552
rect 2590 2548 2594 2552
rect 2638 2698 2642 2702
rect 2622 2638 2626 2642
rect 2646 2638 2650 2642
rect 2678 2768 2682 2772
rect 2678 2738 2682 2742
rect 2670 2688 2674 2692
rect 2686 2678 2690 2682
rect 2678 2668 2682 2672
rect 2726 2918 2730 2922
rect 2742 2898 2746 2902
rect 2750 2778 2754 2782
rect 2774 2858 2778 2862
rect 2782 2858 2786 2862
rect 2766 2838 2770 2842
rect 2790 2778 2794 2782
rect 2838 3008 2842 3012
rect 2862 2958 2866 2962
rect 2890 2903 2894 2907
rect 2897 2903 2901 2907
rect 2854 2868 2858 2872
rect 2814 2858 2818 2862
rect 2846 2858 2850 2862
rect 2870 2858 2874 2862
rect 2854 2848 2858 2852
rect 2822 2778 2826 2782
rect 2750 2748 2754 2752
rect 2782 2768 2786 2772
rect 2806 2768 2810 2772
rect 2846 2768 2850 2772
rect 2798 2748 2802 2752
rect 2862 2758 2866 2762
rect 2878 2748 2882 2752
rect 2774 2738 2778 2742
rect 2862 2728 2866 2732
rect 2814 2718 2818 2722
rect 2742 2708 2746 2712
rect 2806 2708 2810 2712
rect 2750 2688 2754 2692
rect 2766 2678 2770 2682
rect 2702 2658 2706 2662
rect 2718 2658 2722 2662
rect 2734 2648 2738 2652
rect 2782 2648 2786 2652
rect 2766 2628 2770 2632
rect 2806 2628 2810 2632
rect 2734 2618 2738 2622
rect 2582 2538 2586 2542
rect 2622 2498 2626 2502
rect 2558 2488 2562 2492
rect 2598 2488 2602 2492
rect 2534 2478 2538 2482
rect 2574 2458 2578 2462
rect 2534 2448 2538 2452
rect 2542 2448 2546 2452
rect 2622 2448 2626 2452
rect 2558 2428 2562 2432
rect 2550 2408 2554 2412
rect 2534 2398 2538 2402
rect 2678 2598 2682 2602
rect 2654 2548 2658 2552
rect 2662 2548 2666 2552
rect 2726 2558 2730 2562
rect 2758 2558 2762 2562
rect 2702 2548 2706 2552
rect 2718 2548 2722 2552
rect 2790 2558 2794 2562
rect 2798 2548 2802 2552
rect 2782 2538 2786 2542
rect 2678 2528 2682 2532
rect 2670 2508 2674 2512
rect 2742 2528 2746 2532
rect 2734 2508 2738 2512
rect 2694 2488 2698 2492
rect 2702 2488 2706 2492
rect 2726 2478 2730 2482
rect 2694 2468 2698 2472
rect 2710 2468 2714 2472
rect 2782 2508 2786 2512
rect 2822 2618 2826 2622
rect 2798 2528 2802 2532
rect 2790 2488 2794 2492
rect 2742 2478 2746 2482
rect 2774 2478 2778 2482
rect 2806 2518 2810 2522
rect 2758 2468 2762 2472
rect 2718 2458 2722 2462
rect 2750 2458 2754 2462
rect 2686 2428 2690 2432
rect 2742 2428 2746 2432
rect 2782 2468 2786 2472
rect 2662 2408 2666 2412
rect 2750 2408 2754 2412
rect 2766 2408 2770 2412
rect 2662 2398 2666 2402
rect 2726 2398 2730 2402
rect 2566 2388 2570 2392
rect 2638 2388 2642 2392
rect 2646 2388 2650 2392
rect 2622 2378 2626 2382
rect 2614 2368 2618 2372
rect 2606 2358 2610 2362
rect 2558 2348 2562 2352
rect 2542 2328 2546 2332
rect 2574 2328 2578 2332
rect 2590 2328 2594 2332
rect 2566 2318 2570 2322
rect 2534 2308 2538 2312
rect 2526 2288 2530 2292
rect 2486 2268 2490 2272
rect 2478 2258 2482 2262
rect 2566 2268 2570 2272
rect 2550 2248 2554 2252
rect 2510 2238 2514 2242
rect 2526 2238 2530 2242
rect 2502 2228 2506 2232
rect 2494 2208 2498 2212
rect 2526 2208 2530 2212
rect 2462 2148 2466 2152
rect 2510 2148 2514 2152
rect 2470 2128 2474 2132
rect 2462 2108 2466 2112
rect 2462 2078 2466 2082
rect 2454 2058 2458 2062
rect 2486 2098 2490 2102
rect 2542 2198 2546 2202
rect 2534 2118 2538 2122
rect 2510 2048 2514 2052
rect 2494 2038 2498 2042
rect 2542 2038 2546 2042
rect 2518 2008 2522 2012
rect 2502 1988 2506 1992
rect 2454 1968 2458 1972
rect 2470 1968 2474 1972
rect 2486 1968 2490 1972
rect 2446 1958 2450 1962
rect 2438 1948 2442 1952
rect 2566 2188 2570 2192
rect 2614 2318 2618 2322
rect 2606 2308 2610 2312
rect 2630 2358 2634 2362
rect 2654 2358 2658 2362
rect 2710 2358 2714 2362
rect 2646 2348 2650 2352
rect 2854 2698 2858 2702
rect 2838 2688 2842 2692
rect 2886 2728 2890 2732
rect 2890 2703 2894 2707
rect 2897 2703 2901 2707
rect 2894 2658 2898 2662
rect 2902 2638 2906 2642
rect 2926 3078 2930 3082
rect 2926 3058 2930 3062
rect 2990 3248 2994 3252
rect 2974 3238 2978 3242
rect 2982 3198 2986 3202
rect 2958 3158 2962 3162
rect 2950 3138 2954 3142
rect 2966 3148 2970 3152
rect 2990 3158 2994 3162
rect 3038 3408 3042 3412
rect 3262 3508 3266 3512
rect 3238 3478 3242 3482
rect 3134 3458 3138 3462
rect 3206 3458 3210 3462
rect 3142 3448 3146 3452
rect 3246 3438 3250 3442
rect 3126 3418 3130 3422
rect 3182 3418 3186 3422
rect 3198 3418 3202 3422
rect 3230 3418 3234 3422
rect 3070 3368 3074 3372
rect 3102 3368 3106 3372
rect 3046 3358 3050 3362
rect 3142 3368 3146 3372
rect 3166 3358 3170 3362
rect 3006 3348 3010 3352
rect 3038 3348 3042 3352
rect 3086 3348 3090 3352
rect 3126 3348 3130 3352
rect 3046 3338 3050 3342
rect 3054 3338 3058 3342
rect 3094 3338 3098 3342
rect 3206 3328 3210 3332
rect 3086 3308 3090 3312
rect 3102 3298 3106 3302
rect 3166 3298 3170 3302
rect 3014 3288 3018 3292
rect 3062 3288 3066 3292
rect 3126 3278 3130 3282
rect 3062 3268 3066 3272
rect 3006 3198 3010 3202
rect 3046 3198 3050 3202
rect 3006 3168 3010 3172
rect 3054 3158 3058 3162
rect 2998 3148 3002 3152
rect 3118 3228 3122 3232
rect 3134 3228 3138 3232
rect 3102 3218 3106 3222
rect 3118 3198 3122 3202
rect 3126 3158 3130 3162
rect 3142 3208 3146 3212
rect 3142 3158 3146 3162
rect 3198 3158 3202 3162
rect 3182 3148 3186 3152
rect 3110 3128 3114 3132
rect 3174 3138 3178 3142
rect 3166 3118 3170 3122
rect 3070 3108 3074 3112
rect 3006 3098 3010 3102
rect 3054 3088 3058 3092
rect 3118 3088 3122 3092
rect 3022 3058 3026 3062
rect 2942 3048 2946 3052
rect 2982 3038 2986 3042
rect 3062 3068 3066 3072
rect 3094 3068 3098 3072
rect 3126 3068 3130 3072
rect 3078 3058 3082 3062
rect 3086 3048 3090 3052
rect 3094 3048 3098 3052
rect 3142 3048 3146 3052
rect 3078 3038 3082 3042
rect 3030 3028 3034 3032
rect 3046 3018 3050 3022
rect 3014 2998 3018 3002
rect 3070 3008 3074 3012
rect 2990 2958 2994 2962
rect 3030 2958 3034 2962
rect 2942 2948 2946 2952
rect 2974 2948 2978 2952
rect 2998 2938 3002 2942
rect 2990 2928 2994 2932
rect 3030 2928 3034 2932
rect 3070 2928 3074 2932
rect 2942 2858 2946 2862
rect 2942 2818 2946 2822
rect 2926 2768 2930 2772
rect 2926 2758 2930 2762
rect 2934 2758 2938 2762
rect 2918 2748 2922 2752
rect 2918 2708 2922 2712
rect 2918 2598 2922 2602
rect 2910 2558 2914 2562
rect 2846 2548 2850 2552
rect 2886 2548 2890 2552
rect 2902 2548 2906 2552
rect 2838 2538 2842 2542
rect 2926 2538 2930 2542
rect 2966 2868 2970 2872
rect 2950 2758 2954 2762
rect 2958 2758 2962 2762
rect 2950 2748 2954 2752
rect 3014 2868 3018 2872
rect 3006 2798 3010 2802
rect 3014 2778 3018 2782
rect 2966 2708 2970 2712
rect 2998 2708 3002 2712
rect 2990 2688 2994 2692
rect 2990 2668 2994 2672
rect 3054 2858 3058 2862
rect 3046 2828 3050 2832
rect 3030 2808 3034 2812
rect 3022 2768 3026 2772
rect 3038 2778 3042 2782
rect 3030 2688 3034 2692
rect 3022 2668 3026 2672
rect 2990 2658 2994 2662
rect 3006 2658 3010 2662
rect 2966 2648 2970 2652
rect 2950 2638 2954 2642
rect 2990 2618 2994 2622
rect 2974 2568 2978 2572
rect 2974 2558 2978 2562
rect 2958 2548 2962 2552
rect 2998 2568 3002 2572
rect 3022 2558 3026 2562
rect 3030 2558 3034 2562
rect 3070 2748 3074 2752
rect 3078 2658 3082 2662
rect 3062 2638 3066 2642
rect 3206 3098 3210 3102
rect 3246 3398 3250 3402
rect 3230 3368 3234 3372
rect 3254 3368 3258 3372
rect 3254 3338 3258 3342
rect 3230 3318 3234 3322
rect 3222 3268 3226 3272
rect 3238 3258 3242 3262
rect 3222 3168 3226 3172
rect 3222 3138 3226 3142
rect 3238 3168 3242 3172
rect 3214 3088 3218 3092
rect 3206 3078 3210 3082
rect 3158 3028 3162 3032
rect 3174 3028 3178 3032
rect 3102 3018 3106 3022
rect 3174 2998 3178 3002
rect 3182 2978 3186 2982
rect 3198 2978 3202 2982
rect 3158 2958 3162 2962
rect 3150 2948 3154 2952
rect 3094 2868 3098 2872
rect 3142 2888 3146 2892
rect 3134 2878 3138 2882
rect 3126 2858 3130 2862
rect 3126 2848 3130 2852
rect 3110 2808 3114 2812
rect 3102 2748 3106 2752
rect 3174 2868 3178 2872
rect 3198 2968 3202 2972
rect 3198 2958 3202 2962
rect 3254 3268 3258 3272
rect 3286 3758 3290 3762
rect 3342 3988 3346 3992
rect 3358 4008 3362 4012
rect 3374 3998 3378 4002
rect 3374 3988 3378 3992
rect 3350 3868 3354 3872
rect 3402 4203 3406 4207
rect 3409 4203 3413 4207
rect 3406 4138 3410 4142
rect 3446 4218 3450 4222
rect 3470 4168 3474 4172
rect 3542 4498 3546 4502
rect 3502 4478 3506 4482
rect 3710 4708 3714 4712
rect 3638 4638 3642 4642
rect 3686 4638 3690 4642
rect 3734 4728 3738 4732
rect 3742 4688 3746 4692
rect 3774 4918 3778 4922
rect 3862 4958 3866 4962
rect 3878 4948 3882 4952
rect 3982 4948 3986 4952
rect 3822 4928 3826 4932
rect 3822 4918 3826 4922
rect 3806 4868 3810 4872
rect 3798 4818 3802 4822
rect 3974 4908 3978 4912
rect 3922 4903 3926 4907
rect 3929 4903 3933 4907
rect 3934 4888 3938 4892
rect 3854 4858 3858 4862
rect 3838 4848 3842 4852
rect 3790 4798 3794 4802
rect 3806 4798 3810 4802
rect 3774 4758 3778 4762
rect 3766 4738 3770 4742
rect 3774 4708 3778 4712
rect 3758 4668 3762 4672
rect 3774 4658 3778 4662
rect 3742 4648 3746 4652
rect 3750 4648 3754 4652
rect 3726 4618 3730 4622
rect 3622 4588 3626 4592
rect 3726 4578 3730 4582
rect 3614 4558 3618 4562
rect 3654 4548 3658 4552
rect 3678 4548 3682 4552
rect 3710 4548 3714 4552
rect 3574 4538 3578 4542
rect 3566 4508 3570 4512
rect 3550 4488 3554 4492
rect 3582 4488 3586 4492
rect 3670 4538 3674 4542
rect 3662 4528 3666 4532
rect 3910 4838 3914 4842
rect 4006 4908 4010 4912
rect 3998 4868 4002 4872
rect 3958 4858 3962 4862
rect 3950 4838 3954 4842
rect 3926 4828 3930 4832
rect 3814 4768 3818 4772
rect 3838 4768 3842 4772
rect 3950 4768 3954 4772
rect 3846 4758 3850 4762
rect 3870 4758 3874 4762
rect 3910 4758 3914 4762
rect 3878 4748 3882 4752
rect 3854 4738 3858 4742
rect 3830 4708 3834 4712
rect 3798 4688 3802 4692
rect 3862 4678 3866 4682
rect 3862 4668 3866 4672
rect 3922 4703 3926 4707
rect 3929 4703 3933 4707
rect 3902 4698 3906 4702
rect 3886 4688 3890 4692
rect 3910 4678 3914 4682
rect 3814 4658 3818 4662
rect 3870 4658 3874 4662
rect 3790 4648 3794 4652
rect 3814 4638 3818 4642
rect 3822 4608 3826 4612
rect 3814 4598 3818 4602
rect 3806 4548 3810 4552
rect 3838 4588 3842 4592
rect 3830 4558 3834 4562
rect 3878 4558 3882 4562
rect 3734 4538 3738 4542
rect 3702 4518 3706 4522
rect 3694 4498 3698 4502
rect 3670 4488 3674 4492
rect 3686 4478 3690 4482
rect 3566 4468 3570 4472
rect 3614 4468 3618 4472
rect 3502 4428 3506 4432
rect 3494 4418 3498 4422
rect 3486 4388 3490 4392
rect 3494 4318 3498 4322
rect 3518 4358 3522 4362
rect 3542 4458 3546 4462
rect 3566 4458 3570 4462
rect 3566 4448 3570 4452
rect 3534 4438 3538 4442
rect 3614 4388 3618 4392
rect 3662 4388 3666 4392
rect 3558 4368 3562 4372
rect 3550 4358 3554 4362
rect 3622 4378 3626 4382
rect 3534 4348 3538 4352
rect 3550 4348 3554 4352
rect 3510 4328 3514 4332
rect 3486 4238 3490 4242
rect 3502 4178 3506 4182
rect 3478 4158 3482 4162
rect 3526 4308 3530 4312
rect 3542 4338 3546 4342
rect 3542 4328 3546 4332
rect 3550 4298 3554 4302
rect 3638 4338 3642 4342
rect 3630 4288 3634 4292
rect 3590 4258 3594 4262
rect 3606 4258 3610 4262
rect 3526 4248 3530 4252
rect 3558 4248 3562 4252
rect 3630 4248 3634 4252
rect 3550 4228 3554 4232
rect 3558 4228 3562 4232
rect 3614 4218 3618 4222
rect 3526 4168 3530 4172
rect 3510 4158 3514 4162
rect 3518 4158 3522 4162
rect 3478 4148 3482 4152
rect 3510 4148 3514 4152
rect 3454 4138 3458 4142
rect 3446 4128 3450 4132
rect 3470 4108 3474 4112
rect 3494 4108 3498 4112
rect 3494 4098 3498 4102
rect 3438 4088 3442 4092
rect 3454 4078 3458 4082
rect 3390 4058 3394 4062
rect 3430 4059 3434 4063
rect 3558 4138 3562 4142
rect 3542 4128 3546 4132
rect 3566 4128 3570 4132
rect 3470 4058 3474 4062
rect 3502 4058 3506 4062
rect 3422 4008 3426 4012
rect 3402 4003 3406 4007
rect 3409 4003 3413 4007
rect 3430 3978 3434 3982
rect 3430 3958 3434 3962
rect 3382 3948 3386 3952
rect 3390 3938 3394 3942
rect 3366 3898 3370 3902
rect 3374 3898 3378 3902
rect 3358 3858 3362 3862
rect 3366 3828 3370 3832
rect 3286 3738 3290 3742
rect 3326 3738 3330 3742
rect 3278 3498 3282 3502
rect 3286 3478 3290 3482
rect 3278 3458 3282 3462
rect 3334 3728 3338 3732
rect 3342 3688 3346 3692
rect 3342 3668 3346 3672
rect 3382 3888 3386 3892
rect 3406 3888 3410 3892
rect 3438 3868 3442 3872
rect 3382 3848 3386 3852
rect 3402 3803 3406 3807
rect 3409 3803 3413 3807
rect 3526 4028 3530 4032
rect 3542 4028 3546 4032
rect 3494 4018 3498 4022
rect 3550 4018 3554 4022
rect 3486 4008 3490 4012
rect 3486 3948 3490 3952
rect 3454 3918 3458 3922
rect 3502 3958 3506 3962
rect 3518 3948 3522 3952
rect 3526 3938 3530 3942
rect 3470 3928 3474 3932
rect 3494 3918 3498 3922
rect 3542 3918 3546 3922
rect 3462 3908 3466 3912
rect 3534 3888 3538 3892
rect 3526 3868 3530 3872
rect 3542 3878 3546 3882
rect 3494 3848 3498 3852
rect 3542 3848 3546 3852
rect 3494 3838 3498 3842
rect 3398 3778 3402 3782
rect 3446 3778 3450 3782
rect 3390 3748 3394 3752
rect 3366 3738 3370 3742
rect 3382 3738 3386 3742
rect 3478 3758 3482 3762
rect 3502 3798 3506 3802
rect 3526 3778 3530 3782
rect 3486 3748 3490 3752
rect 3414 3738 3418 3742
rect 3462 3738 3466 3742
rect 3454 3728 3458 3732
rect 3374 3688 3378 3692
rect 3334 3658 3338 3662
rect 3350 3658 3354 3662
rect 3366 3658 3370 3662
rect 3318 3648 3322 3652
rect 3318 3638 3322 3642
rect 3326 3588 3330 3592
rect 3326 3558 3330 3562
rect 3358 3548 3362 3552
rect 3310 3508 3314 3512
rect 3326 3459 3330 3463
rect 3302 3448 3306 3452
rect 3350 3428 3354 3432
rect 3318 3418 3322 3422
rect 3366 3418 3370 3422
rect 3294 3408 3298 3412
rect 3358 3368 3362 3372
rect 3278 3358 3282 3362
rect 3286 3348 3290 3352
rect 3334 3328 3338 3332
rect 3270 3298 3274 3302
rect 3294 3288 3298 3292
rect 3286 3268 3290 3272
rect 3318 3268 3322 3272
rect 3270 3258 3274 3262
rect 3254 3238 3258 3242
rect 3350 3348 3354 3352
rect 3422 3668 3426 3672
rect 3454 3668 3458 3672
rect 3494 3708 3498 3712
rect 3718 4488 3722 4492
rect 3774 4518 3778 4522
rect 3766 4508 3770 4512
rect 3726 4468 3730 4472
rect 3710 4458 3714 4462
rect 3734 4438 3738 4442
rect 3710 4408 3714 4412
rect 3694 4388 3698 4392
rect 3806 4538 3810 4542
rect 3790 4458 3794 4462
rect 3798 4448 3802 4452
rect 3766 4378 3770 4382
rect 3782 4378 3786 4382
rect 3686 4358 3690 4362
rect 3678 4298 3682 4302
rect 3654 4268 3658 4272
rect 3670 4238 3674 4242
rect 3614 4168 3618 4172
rect 3622 4158 3626 4162
rect 3662 4158 3666 4162
rect 3622 4108 3626 4112
rect 3606 4078 3610 4082
rect 3638 4098 3642 4102
rect 3638 4078 3642 4082
rect 3590 4048 3594 4052
rect 3598 4018 3602 4022
rect 3574 3988 3578 3992
rect 3558 3968 3562 3972
rect 3718 4348 3722 4352
rect 3774 4348 3778 4352
rect 3790 4348 3794 4352
rect 3758 4338 3762 4342
rect 3766 4338 3770 4342
rect 3822 4488 3826 4492
rect 3846 4548 3850 4552
rect 3878 4548 3882 4552
rect 3878 4508 3882 4512
rect 3846 4498 3850 4502
rect 3854 4498 3858 4502
rect 3878 4498 3882 4502
rect 3838 4478 3842 4482
rect 3854 4488 3858 4492
rect 3862 4488 3866 4492
rect 3822 4458 3826 4462
rect 3838 4448 3842 4452
rect 3870 4478 3874 4482
rect 3902 4538 3906 4542
rect 3918 4538 3922 4542
rect 3974 4818 3978 4822
rect 3990 4838 3994 4842
rect 3982 4798 3986 4802
rect 4086 5058 4090 5062
rect 4222 5058 4226 5062
rect 4310 5048 4314 5052
rect 4286 5038 4290 5042
rect 4206 5028 4210 5032
rect 4342 5028 4346 5032
rect 4142 5018 4146 5022
rect 4302 4998 4306 5002
rect 4246 4968 4250 4972
rect 4070 4958 4074 4962
rect 4230 4958 4234 4962
rect 4134 4948 4138 4952
rect 4046 4918 4050 4922
rect 4054 4918 4058 4922
rect 4022 4868 4026 4872
rect 4014 4858 4018 4862
rect 3990 4778 3994 4782
rect 3998 4778 4002 4782
rect 3998 4768 4002 4772
rect 3982 4758 3986 4762
rect 4006 4748 4010 4752
rect 3958 4738 3962 4742
rect 3990 4728 3994 4732
rect 3998 4728 4002 4732
rect 3966 4668 3970 4672
rect 3990 4668 3994 4672
rect 4022 4848 4026 4852
rect 4134 4928 4138 4932
rect 4166 4948 4170 4952
rect 4246 4948 4250 4952
rect 4142 4918 4146 4922
rect 4158 4918 4162 4922
rect 4102 4888 4106 4892
rect 4118 4878 4122 4882
rect 4054 4868 4058 4872
rect 4110 4868 4114 4872
rect 4086 4858 4090 4862
rect 4118 4858 4122 4862
rect 4142 4858 4146 4862
rect 4046 4848 4050 4852
rect 4078 4848 4082 4852
rect 4038 4808 4042 4812
rect 4046 4778 4050 4782
rect 4030 4748 4034 4752
rect 4046 4738 4050 4742
rect 4094 4848 4098 4852
rect 4102 4848 4106 4852
rect 4086 4778 4090 4782
rect 4070 4758 4074 4762
rect 4062 4708 4066 4712
rect 4014 4658 4018 4662
rect 4030 4658 4034 4662
rect 3990 4648 3994 4652
rect 3998 4628 4002 4632
rect 3942 4578 3946 4582
rect 3966 4568 3970 4572
rect 3950 4538 3954 4542
rect 3982 4528 3986 4532
rect 3894 4438 3898 4442
rect 3878 4378 3882 4382
rect 3922 4503 3926 4507
rect 3929 4503 3933 4507
rect 3942 4488 3946 4492
rect 4006 4488 4010 4492
rect 3910 4468 3914 4472
rect 3942 4368 3946 4372
rect 3838 4358 3842 4362
rect 3846 4358 3850 4362
rect 3862 4358 3866 4362
rect 3894 4358 3898 4362
rect 3902 4358 3906 4362
rect 3814 4338 3818 4342
rect 3798 4328 3802 4332
rect 3766 4308 3770 4312
rect 3822 4328 3826 4332
rect 3830 4328 3834 4332
rect 3838 4308 3842 4312
rect 3790 4298 3794 4302
rect 3806 4298 3810 4302
rect 3822 4278 3826 4282
rect 3734 4268 3738 4272
rect 3694 4258 3698 4262
rect 3710 4258 3714 4262
rect 3750 4258 3754 4262
rect 3702 4248 3706 4252
rect 3686 4128 3690 4132
rect 3726 4178 3730 4182
rect 3734 4158 3738 4162
rect 3742 4148 3746 4152
rect 3718 4088 3722 4092
rect 3710 4078 3714 4082
rect 3782 4258 3786 4262
rect 3886 4348 3890 4352
rect 3926 4348 3930 4352
rect 3854 4338 3858 4342
rect 3878 4338 3882 4342
rect 3870 4308 3874 4312
rect 3922 4303 3926 4307
rect 3929 4303 3933 4307
rect 3902 4288 3906 4292
rect 3910 4288 3914 4292
rect 4030 4648 4034 4652
rect 4038 4588 4042 4592
rect 4062 4618 4066 4622
rect 4062 4568 4066 4572
rect 4206 4938 4210 4942
rect 4190 4928 4194 4932
rect 4190 4918 4194 4922
rect 4246 4918 4250 4922
rect 4238 4898 4242 4902
rect 4206 4878 4210 4882
rect 4230 4878 4234 4882
rect 4190 4848 4194 4852
rect 4182 4818 4186 4822
rect 4126 4788 4130 4792
rect 4174 4808 4178 4812
rect 4166 4788 4170 4792
rect 4078 4738 4082 4742
rect 4094 4668 4098 4672
rect 4078 4648 4082 4652
rect 4086 4618 4090 4622
rect 4070 4558 4074 4562
rect 4134 4718 4138 4722
rect 4126 4688 4130 4692
rect 4158 4738 4162 4742
rect 4150 4728 4154 4732
rect 4142 4658 4146 4662
rect 4110 4638 4114 4642
rect 4142 4608 4146 4612
rect 4118 4598 4122 4602
rect 4102 4588 4106 4592
rect 4134 4578 4138 4582
rect 4158 4578 4162 4582
rect 4182 4768 4186 4772
rect 4190 4748 4194 4752
rect 4214 4868 4218 4872
rect 4230 4868 4234 4872
rect 4358 4978 4362 4982
rect 4358 4968 4362 4972
rect 4318 4948 4322 4952
rect 4310 4908 4314 4912
rect 4294 4898 4298 4902
rect 4286 4888 4290 4892
rect 4294 4888 4298 4892
rect 4270 4878 4274 4882
rect 4286 4878 4290 4882
rect 4326 4878 4330 4882
rect 4270 4868 4274 4872
rect 4302 4868 4306 4872
rect 4310 4858 4314 4862
rect 4222 4848 4226 4852
rect 4270 4848 4274 4852
rect 4318 4838 4322 4842
rect 4214 4718 4218 4722
rect 4230 4718 4234 4722
rect 4238 4708 4242 4712
rect 4206 4678 4210 4682
rect 4222 4678 4226 4682
rect 4166 4568 4170 4572
rect 4150 4558 4154 4562
rect 4174 4558 4178 4562
rect 4102 4538 4106 4542
rect 4230 4578 4234 4582
rect 4222 4558 4226 4562
rect 4198 4538 4202 4542
rect 4110 4528 4114 4532
rect 4134 4528 4138 4532
rect 4166 4528 4170 4532
rect 4190 4528 4194 4532
rect 4054 4518 4058 4522
rect 4206 4518 4210 4522
rect 4094 4508 4098 4512
rect 4166 4478 4170 4482
rect 4102 4468 4106 4472
rect 4022 4458 4026 4462
rect 4062 4458 4066 4462
rect 4190 4458 4194 4462
rect 4094 4448 4098 4452
rect 4102 4448 4106 4452
rect 4014 4438 4018 4442
rect 4094 4438 4098 4442
rect 3982 4418 3986 4422
rect 4006 4358 4010 4362
rect 3974 4348 3978 4352
rect 4030 4358 4034 4362
rect 4094 4378 4098 4382
rect 4086 4368 4090 4372
rect 4062 4358 4066 4362
rect 4022 4348 4026 4352
rect 4086 4348 4090 4352
rect 4014 4338 4018 4342
rect 4070 4338 4074 4342
rect 3998 4328 4002 4332
rect 3974 4288 3978 4292
rect 3878 4278 3882 4282
rect 3910 4278 3914 4282
rect 3958 4278 3962 4282
rect 3878 4268 3882 4272
rect 3790 4248 3794 4252
rect 3798 4248 3802 4252
rect 3782 4238 3786 4242
rect 3766 4188 3770 4192
rect 3774 4178 3778 4182
rect 3814 4218 3818 4222
rect 3798 4208 3802 4212
rect 3790 4158 3794 4162
rect 3806 4158 3810 4162
rect 3790 4138 3794 4142
rect 3782 4118 3786 4122
rect 3758 4108 3762 4112
rect 3790 4098 3794 4102
rect 3766 4088 3770 4092
rect 3814 4088 3818 4092
rect 3638 4058 3642 4062
rect 3710 4058 3714 4062
rect 3742 4058 3746 4062
rect 3774 4058 3778 4062
rect 3630 4038 3634 4042
rect 3646 4038 3650 4042
rect 3654 4028 3658 4032
rect 3622 3988 3626 3992
rect 3622 3968 3626 3972
rect 3606 3958 3610 3962
rect 3718 4048 3722 4052
rect 3678 4018 3682 4022
rect 3614 3948 3618 3952
rect 3638 3948 3642 3952
rect 3606 3938 3610 3942
rect 3638 3938 3642 3942
rect 3574 3918 3578 3922
rect 3582 3918 3586 3922
rect 3566 3908 3570 3912
rect 3566 3878 3570 3882
rect 3590 3898 3594 3902
rect 3614 3898 3618 3902
rect 3582 3888 3586 3892
rect 3678 3928 3682 3932
rect 3670 3898 3674 3902
rect 3646 3878 3650 3882
rect 3558 3758 3562 3762
rect 3526 3738 3530 3742
rect 3510 3728 3514 3732
rect 3502 3688 3506 3692
rect 3502 3678 3506 3682
rect 3542 3708 3546 3712
rect 3526 3698 3530 3702
rect 3518 3688 3522 3692
rect 3646 3858 3650 3862
rect 3582 3848 3586 3852
rect 3598 3818 3602 3822
rect 3694 3938 3698 3942
rect 3686 3888 3690 3892
rect 3678 3868 3682 3872
rect 3694 3868 3698 3872
rect 3726 4028 3730 4032
rect 3726 3958 3730 3962
rect 3726 3948 3730 3952
rect 3734 3938 3738 3942
rect 3726 3928 3730 3932
rect 3782 3958 3786 3962
rect 3822 4058 3826 4062
rect 3798 3988 3802 3992
rect 3750 3918 3754 3922
rect 3726 3878 3730 3882
rect 3702 3828 3706 3832
rect 3630 3788 3634 3792
rect 3662 3788 3666 3792
rect 3606 3748 3610 3752
rect 3662 3748 3666 3752
rect 3718 3848 3722 3852
rect 3742 3858 3746 3862
rect 3734 3838 3738 3842
rect 3750 3838 3754 3842
rect 3782 3828 3786 3832
rect 3710 3808 3714 3812
rect 3726 3778 3730 3782
rect 3718 3758 3722 3762
rect 3574 3688 3578 3692
rect 3550 3668 3554 3672
rect 3574 3668 3578 3672
rect 3470 3658 3474 3662
rect 3390 3648 3394 3652
rect 3558 3648 3562 3652
rect 3422 3618 3426 3622
rect 3478 3618 3482 3622
rect 3402 3603 3406 3607
rect 3409 3603 3413 3607
rect 3390 3598 3394 3602
rect 3422 3598 3426 3602
rect 3454 3588 3458 3592
rect 3430 3568 3434 3572
rect 3406 3548 3410 3552
rect 3470 3558 3474 3562
rect 3494 3558 3498 3562
rect 3502 3558 3506 3562
rect 3478 3538 3482 3542
rect 3494 3538 3498 3542
rect 3502 3538 3506 3542
rect 3446 3528 3450 3532
rect 3430 3518 3434 3522
rect 3446 3518 3450 3522
rect 3430 3488 3434 3492
rect 3398 3478 3402 3482
rect 3518 3638 3522 3642
rect 3526 3638 3530 3642
rect 3590 3648 3594 3652
rect 3606 3658 3610 3662
rect 3614 3648 3618 3652
rect 3598 3618 3602 3622
rect 3590 3598 3594 3602
rect 3542 3588 3546 3592
rect 3574 3588 3578 3592
rect 3590 3588 3594 3592
rect 3542 3558 3546 3562
rect 3534 3548 3538 3552
rect 3542 3538 3546 3542
rect 3606 3538 3610 3542
rect 3606 3498 3610 3502
rect 3542 3488 3546 3492
rect 3574 3488 3578 3492
rect 3558 3478 3562 3482
rect 3550 3468 3554 3472
rect 3566 3468 3570 3472
rect 3510 3458 3514 3462
rect 3454 3428 3458 3432
rect 3542 3458 3546 3462
rect 3558 3458 3562 3462
rect 3582 3458 3586 3462
rect 3518 3418 3522 3422
rect 3402 3403 3406 3407
rect 3409 3403 3413 3407
rect 3414 3378 3418 3382
rect 3358 3308 3362 3312
rect 3366 3288 3370 3292
rect 3342 3278 3346 3282
rect 3326 3248 3330 3252
rect 3334 3248 3338 3252
rect 3318 3178 3322 3182
rect 3286 3158 3290 3162
rect 3358 3148 3362 3152
rect 3254 3138 3258 3142
rect 3270 3078 3274 3082
rect 3302 3088 3306 3092
rect 3326 3078 3330 3082
rect 3318 3068 3322 3072
rect 3350 3068 3354 3072
rect 3246 3058 3250 3062
rect 3246 3018 3250 3022
rect 3230 2968 3234 2972
rect 3198 2938 3202 2942
rect 3206 2928 3210 2932
rect 3190 2888 3194 2892
rect 3198 2868 3202 2872
rect 3270 2998 3274 3002
rect 3222 2948 3226 2952
rect 3230 2948 3234 2952
rect 3254 2948 3258 2952
rect 3334 3058 3338 3062
rect 3382 3278 3386 3282
rect 3542 3438 3546 3442
rect 3542 3428 3546 3432
rect 3526 3388 3530 3392
rect 3486 3368 3490 3372
rect 3430 3358 3434 3362
rect 3462 3358 3466 3362
rect 3438 3348 3442 3352
rect 3446 3338 3450 3342
rect 3422 3318 3426 3322
rect 3438 3308 3442 3312
rect 3454 3288 3458 3292
rect 3550 3358 3554 3362
rect 3486 3348 3490 3352
rect 3470 3288 3474 3292
rect 3590 3408 3594 3412
rect 3598 3368 3602 3372
rect 3566 3358 3570 3362
rect 3582 3358 3586 3362
rect 3534 3338 3538 3342
rect 3558 3338 3562 3342
rect 3566 3338 3570 3342
rect 3590 3338 3594 3342
rect 3598 3328 3602 3332
rect 3526 3318 3530 3322
rect 3558 3278 3562 3282
rect 3582 3278 3586 3282
rect 3446 3268 3450 3272
rect 3502 3268 3506 3272
rect 3534 3268 3538 3272
rect 3430 3258 3434 3262
rect 3470 3258 3474 3262
rect 3558 3258 3562 3262
rect 3398 3238 3402 3242
rect 3414 3228 3418 3232
rect 3462 3238 3466 3242
rect 3422 3218 3426 3222
rect 3334 3038 3338 3042
rect 3246 2938 3250 2942
rect 3238 2928 3242 2932
rect 3286 2928 3290 2932
rect 3302 2928 3306 2932
rect 3222 2918 3226 2922
rect 3246 2908 3250 2912
rect 3238 2888 3242 2892
rect 3270 2888 3274 2892
rect 3262 2858 3266 2862
rect 3278 2858 3282 2862
rect 3302 2858 3306 2862
rect 3222 2838 3226 2842
rect 3270 2828 3274 2832
rect 3150 2748 3154 2752
rect 3166 2748 3170 2752
rect 3206 2748 3210 2752
rect 3238 2748 3242 2752
rect 3262 2748 3266 2752
rect 3174 2718 3178 2722
rect 3158 2668 3162 2672
rect 3134 2658 3138 2662
rect 3150 2638 3154 2642
rect 3126 2618 3130 2622
rect 3086 2558 3090 2562
rect 3174 2598 3178 2602
rect 3174 2568 3178 2572
rect 3006 2548 3010 2552
rect 3078 2548 3082 2552
rect 3118 2548 3122 2552
rect 3126 2548 3130 2552
rect 2982 2538 2986 2542
rect 2894 2518 2898 2522
rect 2878 2508 2882 2512
rect 2846 2498 2850 2502
rect 2890 2503 2894 2507
rect 2897 2503 2901 2507
rect 2878 2478 2882 2482
rect 2830 2468 2834 2472
rect 2846 2468 2850 2472
rect 2862 2468 2866 2472
rect 2798 2458 2802 2462
rect 2846 2448 2850 2452
rect 2838 2428 2842 2432
rect 2878 2468 2882 2472
rect 2878 2428 2882 2432
rect 2894 2428 2898 2432
rect 2798 2408 2802 2412
rect 2790 2398 2794 2402
rect 2750 2378 2754 2382
rect 2734 2368 2738 2372
rect 2790 2368 2794 2372
rect 2774 2358 2778 2362
rect 2638 2338 2642 2342
rect 2670 2338 2674 2342
rect 2686 2338 2690 2342
rect 2662 2328 2666 2332
rect 2638 2318 2642 2322
rect 2622 2308 2626 2312
rect 2662 2308 2666 2312
rect 2638 2298 2642 2302
rect 2646 2298 2650 2302
rect 2702 2328 2706 2332
rect 2630 2288 2634 2292
rect 2678 2288 2682 2292
rect 2590 2258 2594 2262
rect 2630 2248 2634 2252
rect 2574 2168 2578 2172
rect 2606 2168 2610 2172
rect 2726 2298 2730 2302
rect 2846 2368 2850 2372
rect 2830 2358 2834 2362
rect 2870 2408 2874 2412
rect 2838 2348 2842 2352
rect 2854 2348 2858 2352
rect 2918 2508 2922 2512
rect 2926 2498 2930 2502
rect 2918 2368 2922 2372
rect 2894 2348 2898 2352
rect 2814 2338 2818 2342
rect 2854 2338 2858 2342
rect 2886 2338 2890 2342
rect 2774 2298 2778 2302
rect 2822 2308 2826 2312
rect 2838 2298 2842 2302
rect 2890 2303 2894 2307
rect 2897 2303 2901 2307
rect 2990 2528 2994 2532
rect 2958 2468 2962 2472
rect 2990 2468 2994 2472
rect 2958 2458 2962 2462
rect 2974 2458 2978 2462
rect 2942 2448 2946 2452
rect 2982 2448 2986 2452
rect 2934 2408 2938 2412
rect 2934 2358 2938 2362
rect 2926 2308 2930 2312
rect 2862 2288 2866 2292
rect 2902 2288 2906 2292
rect 2742 2278 2746 2282
rect 2686 2268 2690 2272
rect 2718 2268 2722 2272
rect 2854 2268 2858 2272
rect 2886 2268 2890 2272
rect 2670 2258 2674 2262
rect 2694 2258 2698 2262
rect 2710 2258 2714 2262
rect 2734 2258 2738 2262
rect 2694 2248 2698 2252
rect 2726 2248 2730 2252
rect 2718 2228 2722 2232
rect 2742 2228 2746 2232
rect 2734 2208 2738 2212
rect 2742 2198 2746 2202
rect 2710 2178 2714 2182
rect 2566 2148 2570 2152
rect 2622 2148 2626 2152
rect 2654 2148 2658 2152
rect 2718 2148 2722 2152
rect 2614 2138 2618 2142
rect 2670 2138 2674 2142
rect 2702 2138 2706 2142
rect 2558 2128 2562 2132
rect 2558 2118 2562 2122
rect 2550 1978 2554 1982
rect 2646 2098 2650 2102
rect 2622 2078 2626 2082
rect 2574 2058 2578 2062
rect 2598 2048 2602 2052
rect 2630 2048 2634 2052
rect 2598 2028 2602 2032
rect 2574 2018 2578 2022
rect 2694 2058 2698 2062
rect 2678 2048 2682 2052
rect 2566 2008 2570 2012
rect 2582 2008 2586 2012
rect 2662 2008 2666 2012
rect 2558 1968 2562 1972
rect 2486 1948 2490 1952
rect 2518 1948 2522 1952
rect 2502 1928 2506 1932
rect 2510 1928 2514 1932
rect 2446 1898 2450 1902
rect 2470 1898 2474 1902
rect 2430 1888 2434 1892
rect 2438 1888 2442 1892
rect 2462 1888 2466 1892
rect 2366 1858 2370 1862
rect 2422 1858 2426 1862
rect 2478 1888 2482 1892
rect 2526 1928 2530 1932
rect 2550 1928 2554 1932
rect 2558 1918 2562 1922
rect 2550 1878 2554 1882
rect 2558 1878 2562 1882
rect 2486 1858 2490 1862
rect 2470 1848 2474 1852
rect 2430 1838 2434 1842
rect 2454 1838 2458 1842
rect 2366 1808 2370 1812
rect 2386 1803 2390 1807
rect 2393 1803 2397 1807
rect 2782 2258 2786 2262
rect 2822 2258 2826 2262
rect 2766 2248 2770 2252
rect 2814 2248 2818 2252
rect 2758 2208 2762 2212
rect 2830 2228 2834 2232
rect 2838 2188 2842 2192
rect 2878 2258 2882 2262
rect 2990 2428 2994 2432
rect 2982 2408 2986 2412
rect 3014 2538 3018 2542
rect 3046 2538 3050 2542
rect 3006 2528 3010 2532
rect 3030 2528 3034 2532
rect 3030 2518 3034 2522
rect 3038 2518 3042 2522
rect 3038 2498 3042 2502
rect 3070 2498 3074 2502
rect 3006 2488 3010 2492
rect 3014 2488 3018 2492
rect 3062 2488 3066 2492
rect 3110 2538 3114 2542
rect 3158 2538 3162 2542
rect 3174 2538 3178 2542
rect 3102 2528 3106 2532
rect 3150 2528 3154 2532
rect 3118 2518 3122 2522
rect 3086 2478 3090 2482
rect 3038 2468 3042 2472
rect 3030 2378 3034 2382
rect 2998 2358 3002 2362
rect 3006 2358 3010 2362
rect 2966 2338 2970 2342
rect 2974 2338 2978 2342
rect 2982 2338 2986 2342
rect 2998 2338 3002 2342
rect 3014 2338 3018 2342
rect 2950 2308 2954 2312
rect 3006 2318 3010 2322
rect 3022 2318 3026 2322
rect 3014 2308 3018 2312
rect 2966 2268 2970 2272
rect 2934 2258 2938 2262
rect 2950 2258 2954 2262
rect 2990 2258 2994 2262
rect 2870 2208 2874 2212
rect 2886 2208 2890 2212
rect 2990 2248 2994 2252
rect 3022 2248 3026 2252
rect 2934 2188 2938 2192
rect 3062 2458 3066 2462
rect 3078 2458 3082 2462
rect 3054 2438 3058 2442
rect 3054 2418 3058 2422
rect 3062 2418 3066 2422
rect 3070 2388 3074 2392
rect 3054 2348 3058 2352
rect 3038 2318 3042 2322
rect 3062 2308 3066 2312
rect 3118 2468 3122 2472
rect 3126 2448 3130 2452
rect 3166 2468 3170 2472
rect 3150 2448 3154 2452
rect 3166 2438 3170 2442
rect 3142 2428 3146 2432
rect 3150 2428 3154 2432
rect 3134 2398 3138 2402
rect 3134 2368 3138 2372
rect 3086 2358 3090 2362
rect 3110 2358 3114 2362
rect 3102 2348 3106 2352
rect 3118 2348 3122 2352
rect 3126 2348 3130 2352
rect 3126 2318 3130 2322
rect 3126 2298 3130 2302
rect 3046 2288 3050 2292
rect 3166 2348 3170 2352
rect 3198 2608 3202 2612
rect 3214 2678 3218 2682
rect 3190 2548 3194 2552
rect 3206 2558 3210 2562
rect 3238 2698 3242 2702
rect 3246 2698 3250 2702
rect 3254 2678 3258 2682
rect 3278 2798 3282 2802
rect 3302 2788 3306 2792
rect 3302 2758 3306 2762
rect 3402 3203 3406 3207
rect 3409 3203 3413 3207
rect 3438 3198 3442 3202
rect 3430 3178 3434 3182
rect 3430 3138 3434 3142
rect 3390 3098 3394 3102
rect 3454 3158 3458 3162
rect 3446 3128 3450 3132
rect 3470 3208 3474 3212
rect 3510 3178 3514 3182
rect 3550 3178 3554 3182
rect 3478 3148 3482 3152
rect 3470 3138 3474 3142
rect 3382 3068 3386 3072
rect 3414 3068 3418 3072
rect 3374 3048 3378 3052
rect 3366 3038 3370 3042
rect 3358 3008 3362 3012
rect 3414 3048 3418 3052
rect 3402 3003 3406 3007
rect 3409 3003 3413 3007
rect 3390 2988 3394 2992
rect 3438 2988 3442 2992
rect 3414 2968 3418 2972
rect 3374 2948 3378 2952
rect 3390 2948 3394 2952
rect 3350 2938 3354 2942
rect 3366 2938 3370 2942
rect 3382 2928 3386 2932
rect 3350 2888 3354 2892
rect 3318 2868 3322 2872
rect 3334 2868 3338 2872
rect 3366 2868 3370 2872
rect 3430 2938 3434 2942
rect 3454 3088 3458 3092
rect 3454 3048 3458 3052
rect 3454 3038 3458 3042
rect 3430 2858 3434 2862
rect 3318 2848 3322 2852
rect 3366 2848 3370 2852
rect 3326 2838 3330 2842
rect 3310 2678 3314 2682
rect 3318 2668 3322 2672
rect 3262 2658 3266 2662
rect 3294 2658 3298 2662
rect 3310 2638 3314 2642
rect 3350 2828 3354 2832
rect 3334 2778 3338 2782
rect 3342 2728 3346 2732
rect 3294 2568 3298 2572
rect 3246 2558 3250 2562
rect 3310 2558 3314 2562
rect 3342 2558 3346 2562
rect 3238 2548 3242 2552
rect 3214 2538 3218 2542
rect 3198 2528 3202 2532
rect 3190 2508 3194 2512
rect 3198 2508 3202 2512
rect 3190 2478 3194 2482
rect 3198 2468 3202 2472
rect 3198 2398 3202 2402
rect 3254 2538 3258 2542
rect 3310 2538 3314 2542
rect 3262 2528 3266 2532
rect 3254 2518 3258 2522
rect 3238 2508 3242 2512
rect 3230 2498 3234 2502
rect 3230 2428 3234 2432
rect 3326 2508 3330 2512
rect 3270 2498 3274 2502
rect 3478 3088 3482 3092
rect 3470 3068 3474 3072
rect 3486 3068 3490 3072
rect 3494 3018 3498 3022
rect 3470 3008 3474 3012
rect 3478 2988 3482 2992
rect 3542 3138 3546 3142
rect 3590 3138 3594 3142
rect 3518 3128 3522 3132
rect 3526 3128 3530 3132
rect 3534 3118 3538 3122
rect 3542 3078 3546 3082
rect 3582 3108 3586 3112
rect 3574 3068 3578 3072
rect 3558 2998 3562 3002
rect 3518 2968 3522 2972
rect 3510 2958 3514 2962
rect 3534 2948 3538 2952
rect 3558 2948 3562 2952
rect 3598 3078 3602 3082
rect 3726 3728 3730 3732
rect 3710 3708 3714 3712
rect 3734 3708 3738 3712
rect 3638 3668 3642 3672
rect 3654 3668 3658 3672
rect 3646 3658 3650 3662
rect 3622 3628 3626 3632
rect 3670 3628 3674 3632
rect 3638 3608 3642 3612
rect 3750 3778 3754 3782
rect 3774 3768 3778 3772
rect 3950 4218 3954 4222
rect 4054 4328 4058 4332
rect 4046 4308 4050 4312
rect 4062 4288 4066 4292
rect 4046 4278 4050 4282
rect 4030 4268 4034 4272
rect 4078 4258 4082 4262
rect 4150 4438 4154 4442
rect 4198 4438 4202 4442
rect 4158 4428 4162 4432
rect 4166 4398 4170 4402
rect 4134 4358 4138 4362
rect 4118 4348 4122 4352
rect 4150 4348 4154 4352
rect 4134 4338 4138 4342
rect 4110 4328 4114 4332
rect 4126 4328 4130 4332
rect 4102 4288 4106 4292
rect 4110 4268 4114 4272
rect 4118 4268 4122 4272
rect 4150 4268 4154 4272
rect 4246 4688 4250 4692
rect 4374 4928 4378 4932
rect 4366 4868 4370 4872
rect 4374 4858 4378 4862
rect 4334 4798 4338 4802
rect 4286 4748 4290 4752
rect 4318 4748 4322 4752
rect 4334 4748 4338 4752
rect 4358 4738 4362 4742
rect 4406 5058 4410 5062
rect 4398 5028 4402 5032
rect 4590 5058 4594 5062
rect 4574 5048 4578 5052
rect 4566 5038 4570 5042
rect 4426 5003 4430 5007
rect 4433 5003 4437 5007
rect 4422 4968 4426 4972
rect 4430 4938 4434 4942
rect 4454 4928 4458 4932
rect 4446 4898 4450 4902
rect 4406 4838 4410 4842
rect 4342 4708 4346 4712
rect 4286 4688 4290 4692
rect 4278 4648 4282 4652
rect 4270 4558 4274 4562
rect 4350 4658 4354 4662
rect 4262 4548 4266 4552
rect 4246 4528 4250 4532
rect 4238 4518 4242 4522
rect 4230 4418 4234 4422
rect 4174 4358 4178 4362
rect 4206 4358 4210 4362
rect 4254 4468 4258 4472
rect 4262 4418 4266 4422
rect 4230 4348 4234 4352
rect 4174 4338 4178 4342
rect 4206 4338 4210 4342
rect 4222 4338 4226 4342
rect 4238 4338 4242 4342
rect 4110 4248 4114 4252
rect 4094 4238 4098 4242
rect 4014 4208 4018 4212
rect 4046 4178 4050 4182
rect 4070 4178 4074 4182
rect 3982 4168 3986 4172
rect 3862 4148 3866 4152
rect 3958 4148 3962 4152
rect 4030 4148 4034 4152
rect 3922 4103 3926 4107
rect 3929 4103 3933 4107
rect 3846 4098 3850 4102
rect 3886 4078 3890 4082
rect 3902 4078 3906 4082
rect 3982 4138 3986 4142
rect 4102 4168 4106 4172
rect 4086 4148 4090 4152
rect 4206 4268 4210 4272
rect 4206 4248 4210 4252
rect 4230 4248 4234 4252
rect 4150 4228 4154 4232
rect 4134 4218 4138 4222
rect 4126 4148 4130 4152
rect 4182 4198 4186 4202
rect 4166 4178 4170 4182
rect 4198 4178 4202 4182
rect 4190 4168 4194 4172
rect 4150 4158 4154 4162
rect 4182 4158 4186 4162
rect 4158 4138 4162 4142
rect 4174 4138 4178 4142
rect 4038 4128 4042 4132
rect 4062 4128 4066 4132
rect 4062 4118 4066 4122
rect 4038 4108 4042 4112
rect 4030 4088 4034 4092
rect 4006 4078 4010 4082
rect 3990 4058 3994 4062
rect 3910 4038 3914 4042
rect 3950 4038 3954 4042
rect 3830 3968 3834 3972
rect 3910 3948 3914 3952
rect 3862 3928 3866 3932
rect 3870 3878 3874 3882
rect 4006 4038 4010 4042
rect 4062 4098 4066 4102
rect 4046 4088 4050 4092
rect 4054 4068 4058 4072
rect 4046 4058 4050 4062
rect 4054 4008 4058 4012
rect 4046 3978 4050 3982
rect 3966 3958 3970 3962
rect 3934 3948 3938 3952
rect 3950 3948 3954 3952
rect 3966 3948 3970 3952
rect 3918 3938 3922 3942
rect 3990 3938 3994 3942
rect 3958 3918 3962 3922
rect 3974 3908 3978 3912
rect 3922 3903 3926 3907
rect 3929 3903 3933 3907
rect 3942 3898 3946 3902
rect 3966 3878 3970 3882
rect 3862 3868 3866 3872
rect 3918 3868 3922 3872
rect 3854 3858 3858 3862
rect 3886 3858 3890 3862
rect 3814 3848 3818 3852
rect 3846 3838 3850 3842
rect 3806 3828 3810 3832
rect 3870 3848 3874 3852
rect 3862 3838 3866 3842
rect 3854 3798 3858 3802
rect 3854 3788 3858 3792
rect 3830 3758 3834 3762
rect 3782 3698 3786 3702
rect 3790 3688 3794 3692
rect 3838 3688 3842 3692
rect 3774 3668 3778 3672
rect 3774 3648 3778 3652
rect 3894 3778 3898 3782
rect 3910 3758 3914 3762
rect 3894 3748 3898 3752
rect 3958 3798 3962 3802
rect 3926 3778 3930 3782
rect 3950 3778 3954 3782
rect 3974 3838 3978 3842
rect 4070 4078 4074 4082
rect 4086 4068 4090 4072
rect 4110 4068 4114 4072
rect 4222 4208 4226 4212
rect 4206 4168 4210 4172
rect 4214 4158 4218 4162
rect 4230 4148 4234 4152
rect 4206 4108 4210 4112
rect 4222 4088 4226 4092
rect 4198 4068 4202 4072
rect 4230 4078 4234 4082
rect 4166 4058 4170 4062
rect 4206 4058 4210 4062
rect 4078 4048 4082 4052
rect 4086 4008 4090 4012
rect 4094 3988 4098 3992
rect 4150 4048 4154 4052
rect 4118 3968 4122 3972
rect 4110 3958 4114 3962
rect 4022 3938 4026 3942
rect 4078 3938 4082 3942
rect 4014 3928 4018 3932
rect 4062 3928 4066 3932
rect 4118 3938 4122 3942
rect 4030 3878 4034 3882
rect 4014 3828 4018 3832
rect 3998 3808 4002 3812
rect 4006 3798 4010 3802
rect 3982 3788 3986 3792
rect 3982 3778 3986 3782
rect 3990 3758 3994 3762
rect 3918 3728 3922 3732
rect 3902 3708 3906 3712
rect 3838 3658 3842 3662
rect 3782 3638 3786 3642
rect 3798 3638 3802 3642
rect 3742 3628 3746 3632
rect 3838 3648 3842 3652
rect 3822 3608 3826 3612
rect 3822 3598 3826 3602
rect 3814 3578 3818 3582
rect 3710 3558 3714 3562
rect 3726 3558 3730 3562
rect 3750 3558 3754 3562
rect 3638 3548 3642 3552
rect 3694 3548 3698 3552
rect 3774 3548 3778 3552
rect 3814 3548 3818 3552
rect 3654 3538 3658 3542
rect 3630 3498 3634 3502
rect 3622 3458 3626 3462
rect 3630 3348 3634 3352
rect 3614 3328 3618 3332
rect 3678 3528 3682 3532
rect 3670 3518 3674 3522
rect 3686 3518 3690 3522
rect 3614 3268 3618 3272
rect 3638 3308 3642 3312
rect 3662 3488 3666 3492
rect 3718 3528 3722 3532
rect 3766 3518 3770 3522
rect 3758 3478 3762 3482
rect 3774 3468 3778 3472
rect 3702 3458 3706 3462
rect 3758 3458 3762 3462
rect 3798 3458 3802 3462
rect 3774 3438 3778 3442
rect 3710 3408 3714 3412
rect 3758 3398 3762 3402
rect 3694 3358 3698 3362
rect 3734 3358 3738 3362
rect 3886 3558 3890 3562
rect 3922 3703 3926 3707
rect 3929 3703 3933 3707
rect 3950 3698 3954 3702
rect 3982 3728 3986 3732
rect 3990 3728 3994 3732
rect 4022 3758 4026 3762
rect 4062 3818 4066 3822
rect 4038 3778 4042 3782
rect 4110 3858 4114 3862
rect 4126 3858 4130 3862
rect 4118 3848 4122 3852
rect 4094 3828 4098 3832
rect 4110 3818 4114 3822
rect 4070 3748 4074 3752
rect 4030 3738 4034 3742
rect 4102 3738 4106 3742
rect 3974 3718 3978 3722
rect 3974 3708 3978 3712
rect 4006 3708 4010 3712
rect 3966 3688 3970 3692
rect 4006 3688 4010 3692
rect 3902 3638 3906 3642
rect 4038 3698 4042 3702
rect 4054 3658 4058 3662
rect 4086 3658 4090 3662
rect 3966 3638 3970 3642
rect 3974 3638 3978 3642
rect 3910 3628 3914 3632
rect 3958 3558 3962 3562
rect 3950 3548 3954 3552
rect 3862 3488 3866 3492
rect 3922 3503 3926 3507
rect 3929 3503 3933 3507
rect 3950 3478 3954 3482
rect 3822 3458 3826 3462
rect 3766 3378 3770 3382
rect 3782 3358 3786 3362
rect 3702 3348 3706 3352
rect 3678 3338 3682 3342
rect 3742 3328 3746 3332
rect 3750 3328 3754 3332
rect 3782 3328 3786 3332
rect 3718 3308 3722 3312
rect 3646 3298 3650 3302
rect 3670 3288 3674 3292
rect 3718 3288 3722 3292
rect 3694 3268 3698 3272
rect 3766 3278 3770 3282
rect 3782 3278 3786 3282
rect 3734 3268 3738 3272
rect 3686 3258 3690 3262
rect 3798 3328 3802 3332
rect 3670 3238 3674 3242
rect 3710 3238 3714 3242
rect 3686 3178 3690 3182
rect 3662 3148 3666 3152
rect 3654 3128 3658 3132
rect 3662 3098 3666 3102
rect 3630 3078 3634 3082
rect 3678 3078 3682 3082
rect 3742 3238 3746 3242
rect 3774 3238 3778 3242
rect 3790 3238 3794 3242
rect 3758 3198 3762 3202
rect 3726 3148 3730 3152
rect 3790 3148 3794 3152
rect 3814 3248 3818 3252
rect 3918 3458 3922 3462
rect 3846 3378 3850 3382
rect 3902 3398 3906 3402
rect 3830 3358 3834 3362
rect 3854 3358 3858 3362
rect 3870 3358 3874 3362
rect 3958 3358 3962 3362
rect 3990 3628 3994 3632
rect 4046 3618 4050 3622
rect 4054 3578 4058 3582
rect 3990 3568 3994 3572
rect 3998 3568 4002 3572
rect 4022 3568 4026 3572
rect 3990 3558 3994 3562
rect 4014 3558 4018 3562
rect 4030 3558 4034 3562
rect 4102 3638 4106 3642
rect 4094 3618 4098 3622
rect 4078 3608 4082 3612
rect 4150 3938 4154 3942
rect 4142 3908 4146 3912
rect 4174 4038 4178 4042
rect 4246 4328 4250 4332
rect 4246 4318 4250 4322
rect 4366 4688 4370 4692
rect 4382 4678 4386 4682
rect 4390 4658 4394 4662
rect 4422 4818 4426 4822
rect 4426 4803 4430 4807
rect 4433 4803 4437 4807
rect 4414 4768 4418 4772
rect 4454 4788 4458 4792
rect 4446 4758 4450 4762
rect 4406 4708 4410 4712
rect 4454 4738 4458 4742
rect 4430 4698 4434 4702
rect 4414 4688 4418 4692
rect 4518 5018 4522 5022
rect 4478 4998 4482 5002
rect 4494 4948 4498 4952
rect 4486 4928 4490 4932
rect 4478 4898 4482 4902
rect 4494 4868 4498 4872
rect 4494 4758 4498 4762
rect 4470 4728 4474 4732
rect 4486 4728 4490 4732
rect 4478 4718 4482 4722
rect 4462 4658 4466 4662
rect 4398 4628 4402 4632
rect 4390 4568 4394 4572
rect 4350 4518 4354 4522
rect 4294 4508 4298 4512
rect 4318 4508 4322 4512
rect 4358 4508 4362 4512
rect 4286 4488 4290 4492
rect 4350 4498 4354 4502
rect 4278 4428 4282 4432
rect 4286 4358 4290 4362
rect 4398 4488 4402 4492
rect 4478 4668 4482 4672
rect 4470 4648 4474 4652
rect 4426 4603 4430 4607
rect 4433 4603 4437 4607
rect 4526 4978 4530 4982
rect 4558 4978 4562 4982
rect 4518 4958 4522 4962
rect 4542 4958 4546 4962
rect 4606 4968 4610 4972
rect 4606 4958 4610 4962
rect 4638 4948 4642 4952
rect 4526 4898 4530 4902
rect 4542 4898 4546 4902
rect 4566 4868 4570 4872
rect 4590 4938 4594 4942
rect 4646 4908 4650 4912
rect 4566 4858 4570 4862
rect 4582 4858 4586 4862
rect 4550 4798 4554 4802
rect 4518 4758 4522 4762
rect 4534 4758 4538 4762
rect 4606 4848 4610 4852
rect 4550 4748 4554 4752
rect 4518 4728 4522 4732
rect 4526 4718 4530 4722
rect 4510 4698 4514 4702
rect 4534 4688 4538 4692
rect 4574 4738 4578 4742
rect 4630 4848 4634 4852
rect 4630 4788 4634 4792
rect 4654 4788 4658 4792
rect 4686 5038 4690 5042
rect 4694 4928 4698 4932
rect 4678 4918 4682 4922
rect 4686 4858 4690 4862
rect 4694 4848 4698 4852
rect 4686 4838 4690 4842
rect 4686 4788 4690 4792
rect 4670 4768 4674 4772
rect 4638 4758 4642 4762
rect 4614 4748 4618 4752
rect 4646 4748 4650 4752
rect 4582 4728 4586 4732
rect 4574 4718 4578 4722
rect 4630 4718 4634 4722
rect 4550 4678 4554 4682
rect 4566 4678 4570 4682
rect 4622 4688 4626 4692
rect 4758 4998 4762 5002
rect 4710 4948 4714 4952
rect 4742 4948 4746 4952
rect 4726 4868 4730 4872
rect 4710 4778 4714 4782
rect 4750 4778 4754 4782
rect 4734 4768 4738 4772
rect 4742 4758 4746 4762
rect 4702 4748 4706 4752
rect 4678 4738 4682 4742
rect 4694 4728 4698 4732
rect 4678 4698 4682 4702
rect 4518 4668 4522 4672
rect 4646 4668 4650 4672
rect 4526 4658 4530 4662
rect 4566 4648 4570 4652
rect 4526 4608 4530 4612
rect 4502 4598 4506 4602
rect 4526 4588 4530 4592
rect 4430 4558 4434 4562
rect 4486 4558 4490 4562
rect 4446 4548 4450 4552
rect 4494 4548 4498 4552
rect 4510 4548 4514 4552
rect 4462 4538 4466 4542
rect 4470 4518 4474 4522
rect 4414 4488 4418 4492
rect 4462 4488 4466 4492
rect 4438 4478 4442 4482
rect 4318 4458 4322 4462
rect 4334 4448 4338 4452
rect 4342 4398 4346 4402
rect 4382 4388 4386 4392
rect 4406 4368 4410 4372
rect 4398 4348 4402 4352
rect 4374 4338 4378 4342
rect 4390 4338 4394 4342
rect 4350 4328 4354 4332
rect 4358 4318 4362 4322
rect 4334 4288 4338 4292
rect 4302 4278 4306 4282
rect 4318 4278 4322 4282
rect 4262 4268 4266 4272
rect 4270 4268 4274 4272
rect 4278 4268 4282 4272
rect 4286 4258 4290 4262
rect 4262 4248 4266 4252
rect 4278 4248 4282 4252
rect 4262 4188 4266 4192
rect 4246 4148 4250 4152
rect 4278 4108 4282 4112
rect 4262 4068 4266 4072
rect 4294 4248 4298 4252
rect 4426 4403 4430 4407
rect 4433 4403 4437 4407
rect 4406 4308 4410 4312
rect 4374 4298 4378 4302
rect 4374 4278 4378 4282
rect 4350 4268 4354 4272
rect 4326 4258 4330 4262
rect 4302 4178 4306 4182
rect 4326 4178 4330 4182
rect 4366 4248 4370 4252
rect 4422 4318 4426 4322
rect 4446 4318 4450 4322
rect 4414 4298 4418 4302
rect 4398 4268 4402 4272
rect 4414 4268 4418 4272
rect 4502 4518 4506 4522
rect 4494 4488 4498 4492
rect 4478 4478 4482 4482
rect 4510 4468 4514 4472
rect 4550 4558 4554 4562
rect 4646 4658 4650 4662
rect 4662 4658 4666 4662
rect 4670 4648 4674 4652
rect 4654 4598 4658 4602
rect 4638 4588 4642 4592
rect 4646 4588 4650 4592
rect 4622 4558 4626 4562
rect 4534 4478 4538 4482
rect 4582 4478 4586 4482
rect 4574 4468 4578 4472
rect 4494 4458 4498 4462
rect 4518 4458 4522 4462
rect 4478 4348 4482 4352
rect 4470 4288 4474 4292
rect 4510 4328 4514 4332
rect 4518 4318 4522 4322
rect 4526 4288 4530 4292
rect 4518 4278 4522 4282
rect 4494 4268 4498 4272
rect 4406 4258 4410 4262
rect 4422 4258 4426 4262
rect 4350 4168 4354 4172
rect 4366 4168 4370 4172
rect 4350 4158 4354 4162
rect 4302 4138 4306 4142
rect 4358 4138 4362 4142
rect 4426 4203 4430 4207
rect 4433 4203 4437 4207
rect 4390 4178 4394 4182
rect 4390 4138 4394 4142
rect 4430 4138 4434 4142
rect 4310 4118 4314 4122
rect 4382 4118 4386 4122
rect 4286 4098 4290 4102
rect 4342 4108 4346 4112
rect 4374 4108 4378 4112
rect 4518 4158 4522 4162
rect 4518 4118 4522 4122
rect 4398 4108 4402 4112
rect 4494 4108 4498 4112
rect 4358 4088 4362 4092
rect 4334 4078 4338 4082
rect 4294 4068 4298 4072
rect 4326 4068 4330 4072
rect 4254 4058 4258 4062
rect 4270 4048 4274 4052
rect 4238 4038 4242 4042
rect 4182 4028 4186 4032
rect 4294 4018 4298 4022
rect 4222 3948 4226 3952
rect 4246 3998 4250 4002
rect 4254 3958 4258 3962
rect 4286 3948 4290 3952
rect 4238 3918 4242 3922
rect 4166 3908 4170 3912
rect 4230 3908 4234 3912
rect 4198 3868 4202 3872
rect 4158 3858 4162 3862
rect 4158 3828 4162 3832
rect 4222 3848 4226 3852
rect 4230 3818 4234 3822
rect 4134 3788 4138 3792
rect 4174 3788 4178 3792
rect 4134 3778 4138 3782
rect 4198 3778 4202 3782
rect 4174 3768 4178 3772
rect 4166 3728 4170 3732
rect 4134 3688 4138 3692
rect 4166 3688 4170 3692
rect 4158 3668 4162 3672
rect 4182 3718 4186 3722
rect 4206 3748 4210 3752
rect 4270 3938 4274 3942
rect 4310 3938 4314 3942
rect 4302 3928 4306 3932
rect 4334 4028 4338 4032
rect 4374 4078 4378 4082
rect 4558 4338 4562 4342
rect 4542 4308 4546 4312
rect 4606 4528 4610 4532
rect 4630 4478 4634 4482
rect 4590 4468 4594 4472
rect 4630 4448 4634 4452
rect 4630 4378 4634 4382
rect 4662 4558 4666 4562
rect 4654 4538 4658 4542
rect 4670 4518 4674 4522
rect 4670 4448 4674 4452
rect 4654 4378 4658 4382
rect 4646 4368 4650 4372
rect 4638 4358 4642 4362
rect 4654 4358 4658 4362
rect 4590 4338 4594 4342
rect 4606 4338 4610 4342
rect 4670 4338 4674 4342
rect 4622 4328 4626 4332
rect 4622 4318 4626 4322
rect 4614 4308 4618 4312
rect 4590 4278 4594 4282
rect 4590 4268 4594 4272
rect 4582 4258 4586 4262
rect 4598 4258 4602 4262
rect 4566 4248 4570 4252
rect 4558 4178 4562 4182
rect 4566 4168 4570 4172
rect 4606 4148 4610 4152
rect 4646 4298 4650 4302
rect 4638 4288 4642 4292
rect 4662 4278 4666 4282
rect 4638 4268 4642 4272
rect 4646 4228 4650 4232
rect 4646 4168 4650 4172
rect 4638 4148 4642 4152
rect 4598 4138 4602 4142
rect 4614 4138 4618 4142
rect 4630 4138 4634 4142
rect 4630 4098 4634 4102
rect 4390 4068 4394 4072
rect 4526 4068 4530 4072
rect 4614 4068 4618 4072
rect 4414 4058 4418 4062
rect 4358 4048 4362 4052
rect 4366 4048 4370 4052
rect 4382 4048 4386 4052
rect 4454 4048 4458 4052
rect 4350 3998 4354 4002
rect 4426 4003 4430 4007
rect 4433 4003 4437 4007
rect 4342 3988 4346 3992
rect 4302 3918 4306 3922
rect 4326 3918 4330 3922
rect 4270 3868 4274 3872
rect 4254 3818 4258 3822
rect 4246 3708 4250 3712
rect 4206 3698 4210 3702
rect 4230 3698 4234 3702
rect 4222 3678 4226 3682
rect 4190 3668 4194 3672
rect 4182 3658 4186 3662
rect 4206 3658 4210 3662
rect 4166 3638 4170 3642
rect 4142 3628 4146 3632
rect 4134 3608 4138 3612
rect 4126 3598 4130 3602
rect 4102 3578 4106 3582
rect 4062 3568 4066 3572
rect 4022 3548 4026 3552
rect 4062 3548 4066 3552
rect 4094 3548 4098 3552
rect 4110 3548 4114 3552
rect 3974 3528 3978 3532
rect 4022 3528 4026 3532
rect 4046 3528 4050 3532
rect 4070 3528 4074 3532
rect 3990 3518 3994 3522
rect 4022 3478 4026 3482
rect 3998 3468 4002 3472
rect 4038 3468 4042 3472
rect 4070 3468 4074 3472
rect 4014 3458 4018 3462
rect 4062 3458 4066 3462
rect 3998 3448 4002 3452
rect 3982 3408 3986 3412
rect 3982 3398 3986 3402
rect 3854 3348 3858 3352
rect 3910 3348 3914 3352
rect 3950 3348 3954 3352
rect 3830 3338 3834 3342
rect 3886 3338 3890 3342
rect 3966 3338 3970 3342
rect 3830 3328 3834 3332
rect 3886 3328 3890 3332
rect 3846 3318 3850 3322
rect 3886 3288 3890 3292
rect 3870 3268 3874 3272
rect 3806 3238 3810 3242
rect 3822 3238 3826 3242
rect 3854 3218 3858 3222
rect 3958 3328 3962 3332
rect 3942 3308 3946 3312
rect 3922 3303 3926 3307
rect 3929 3303 3933 3307
rect 3910 3288 3914 3292
rect 3990 3288 3994 3292
rect 4014 3288 4018 3292
rect 4094 3518 4098 3522
rect 4118 3498 4122 3502
rect 4126 3488 4130 3492
rect 4126 3448 4130 3452
rect 4086 3438 4090 3442
rect 4078 3418 4082 3422
rect 4062 3378 4066 3382
rect 4030 3338 4034 3342
rect 3942 3278 3946 3282
rect 4022 3278 4026 3282
rect 3990 3268 3994 3272
rect 3942 3258 3946 3262
rect 4022 3258 4026 3262
rect 3918 3248 3922 3252
rect 3894 3158 3898 3162
rect 3806 3148 3810 3152
rect 3838 3148 3842 3152
rect 3862 3148 3866 3152
rect 3854 3138 3858 3142
rect 3798 3118 3802 3122
rect 3758 3088 3762 3092
rect 3766 3088 3770 3092
rect 3718 3078 3722 3082
rect 3806 3078 3810 3082
rect 3590 3068 3594 3072
rect 3606 3068 3610 3072
rect 3662 3068 3666 3072
rect 3670 3068 3674 3072
rect 3630 3058 3634 3062
rect 3638 3058 3642 3062
rect 3694 3058 3698 3062
rect 3750 3058 3754 3062
rect 3622 3048 3626 3052
rect 3710 3048 3714 3052
rect 3718 3038 3722 3042
rect 3590 3028 3594 3032
rect 3678 3028 3682 3032
rect 3598 2998 3602 3002
rect 3478 2938 3482 2942
rect 3534 2938 3538 2942
rect 3510 2918 3514 2922
rect 3518 2888 3522 2892
rect 3494 2868 3498 2872
rect 3526 2868 3530 2872
rect 3462 2838 3466 2842
rect 3646 2948 3650 2952
rect 3630 2938 3634 2942
rect 3574 2928 3578 2932
rect 3566 2918 3570 2922
rect 3550 2898 3554 2902
rect 3542 2888 3546 2892
rect 3550 2888 3554 2892
rect 3542 2868 3546 2872
rect 3558 2868 3562 2872
rect 3590 2868 3594 2872
rect 3646 2888 3650 2892
rect 3622 2858 3626 2862
rect 3542 2848 3546 2852
rect 3574 2848 3578 2852
rect 3582 2848 3586 2852
rect 3462 2818 3466 2822
rect 3494 2818 3498 2822
rect 3534 2818 3538 2822
rect 3558 2818 3562 2822
rect 3390 2808 3394 2812
rect 3422 2808 3426 2812
rect 3402 2803 3406 2807
rect 3409 2803 3413 2807
rect 3390 2748 3394 2752
rect 3422 2748 3426 2752
rect 3358 2728 3362 2732
rect 3390 2728 3394 2732
rect 3382 2638 3386 2642
rect 3430 2638 3434 2642
rect 3398 2628 3402 2632
rect 3402 2603 3406 2607
rect 3409 2603 3413 2607
rect 3382 2568 3386 2572
rect 3374 2558 3378 2562
rect 3406 2558 3410 2562
rect 3382 2548 3386 2552
rect 3390 2548 3394 2552
rect 3406 2528 3410 2532
rect 3358 2498 3362 2502
rect 3254 2478 3258 2482
rect 3278 2478 3282 2482
rect 3294 2478 3298 2482
rect 3326 2478 3330 2482
rect 3350 2478 3354 2482
rect 3374 2478 3378 2482
rect 3270 2468 3274 2472
rect 3342 2468 3346 2472
rect 3358 2468 3362 2472
rect 3254 2448 3258 2452
rect 3246 2428 3250 2432
rect 3230 2418 3234 2422
rect 3214 2358 3218 2362
rect 3254 2408 3258 2412
rect 3254 2368 3258 2372
rect 3198 2348 3202 2352
rect 3238 2348 3242 2352
rect 3254 2348 3258 2352
rect 3158 2338 3162 2342
rect 3166 2328 3170 2332
rect 3198 2328 3202 2332
rect 3198 2318 3202 2322
rect 3182 2288 3186 2292
rect 3110 2268 3114 2272
rect 3134 2268 3138 2272
rect 3158 2268 3162 2272
rect 3206 2288 3210 2292
rect 3302 2458 3306 2462
rect 3334 2458 3338 2462
rect 3350 2458 3354 2462
rect 3294 2358 3298 2362
rect 3222 2328 3226 2332
rect 3262 2328 3266 2332
rect 3222 2298 3226 2302
rect 3214 2268 3218 2272
rect 3294 2328 3298 2332
rect 3318 2438 3322 2442
rect 3358 2388 3362 2392
rect 3318 2378 3322 2382
rect 3398 2458 3402 2462
rect 3374 2398 3378 2402
rect 3366 2378 3370 2382
rect 3350 2358 3354 2362
rect 3366 2358 3370 2362
rect 3478 2788 3482 2792
rect 3470 2758 3474 2762
rect 3494 2758 3498 2762
rect 3470 2738 3474 2742
rect 3446 2708 3450 2712
rect 3454 2678 3458 2682
rect 3454 2628 3458 2632
rect 3510 2748 3514 2752
rect 3518 2748 3522 2752
rect 3478 2708 3482 2712
rect 3542 2728 3546 2732
rect 3502 2708 3506 2712
rect 3518 2678 3522 2682
rect 3494 2668 3498 2672
rect 3518 2668 3522 2672
rect 3622 2798 3626 2802
rect 3638 2798 3642 2802
rect 3654 2778 3658 2782
rect 3566 2758 3570 2762
rect 3606 2758 3610 2762
rect 3678 2728 3682 2732
rect 3622 2698 3626 2702
rect 3598 2668 3602 2672
rect 3614 2668 3618 2672
rect 3542 2658 3546 2662
rect 3558 2658 3562 2662
rect 3590 2658 3594 2662
rect 3486 2638 3490 2642
rect 3542 2638 3546 2642
rect 3734 2998 3738 3002
rect 3846 3058 3850 3062
rect 3782 3028 3786 3032
rect 3814 3028 3818 3032
rect 3718 2988 3722 2992
rect 3742 2988 3746 2992
rect 3806 2978 3810 2982
rect 3758 2968 3762 2972
rect 3702 2958 3706 2962
rect 3694 2848 3698 2852
rect 3694 2798 3698 2802
rect 3686 2708 3690 2712
rect 3662 2688 3666 2692
rect 3686 2688 3690 2692
rect 3654 2668 3658 2672
rect 3646 2658 3650 2662
rect 3670 2658 3674 2662
rect 3502 2618 3506 2622
rect 3622 2618 3626 2622
rect 3550 2598 3554 2602
rect 3566 2598 3570 2602
rect 3582 2568 3586 2572
rect 3486 2538 3490 2542
rect 3518 2538 3522 2542
rect 3566 2538 3570 2542
rect 3598 2538 3602 2542
rect 3478 2528 3482 2532
rect 3542 2528 3546 2532
rect 3638 2538 3642 2542
rect 3678 2538 3682 2542
rect 3454 2518 3458 2522
rect 3614 2518 3618 2522
rect 3630 2518 3634 2522
rect 3446 2498 3450 2502
rect 3486 2478 3490 2482
rect 3494 2468 3498 2472
rect 3510 2468 3514 2472
rect 3542 2468 3546 2472
rect 3550 2468 3554 2472
rect 3526 2458 3530 2462
rect 3446 2418 3450 2422
rect 3438 2408 3442 2412
rect 3402 2403 3406 2407
rect 3409 2403 3413 2407
rect 3438 2398 3442 2402
rect 3422 2388 3426 2392
rect 3414 2378 3418 2382
rect 3398 2358 3402 2362
rect 3334 2348 3338 2352
rect 3350 2348 3354 2352
rect 3382 2348 3386 2352
rect 3342 2338 3346 2342
rect 3326 2328 3330 2332
rect 3310 2318 3314 2322
rect 3286 2308 3290 2312
rect 3286 2298 3290 2302
rect 3270 2288 3274 2292
rect 3278 2288 3282 2292
rect 3246 2268 3250 2272
rect 3254 2268 3258 2272
rect 3014 2218 3018 2222
rect 3030 2218 3034 2222
rect 3086 2218 3090 2222
rect 3126 2218 3130 2222
rect 3182 2218 3186 2222
rect 3046 2208 3050 2212
rect 2942 2178 2946 2182
rect 2862 2158 2866 2162
rect 2974 2158 2978 2162
rect 3054 2158 3058 2162
rect 2782 2148 2786 2152
rect 2758 2138 2762 2142
rect 2766 2138 2770 2142
rect 2758 2118 2762 2122
rect 2782 2128 2786 2132
rect 2766 2108 2770 2112
rect 2814 2098 2818 2102
rect 2750 2078 2754 2082
rect 2814 2078 2818 2082
rect 2742 2068 2746 2072
rect 2734 2058 2738 2062
rect 2822 2068 2826 2072
rect 2822 2058 2826 2062
rect 2630 1988 2634 1992
rect 2686 1988 2690 1992
rect 2710 1988 2714 1992
rect 2598 1968 2602 1972
rect 2590 1958 2594 1962
rect 2670 1958 2674 1962
rect 2694 1958 2698 1962
rect 2614 1948 2618 1952
rect 2662 1948 2666 1952
rect 2678 1938 2682 1942
rect 2614 1928 2618 1932
rect 2606 1918 2610 1922
rect 2574 1898 2578 1902
rect 2574 1888 2578 1892
rect 2606 1888 2610 1892
rect 2566 1858 2570 1862
rect 2510 1848 2514 1852
rect 2542 1848 2546 1852
rect 2566 1848 2570 1852
rect 2494 1798 2498 1802
rect 2406 1758 2410 1762
rect 2422 1758 2426 1762
rect 2590 1858 2594 1862
rect 2646 1928 2650 1932
rect 2654 1918 2658 1922
rect 2630 1888 2634 1892
rect 2678 1888 2682 1892
rect 2638 1858 2642 1862
rect 2678 1858 2682 1862
rect 2614 1848 2618 1852
rect 2670 1848 2674 1852
rect 2702 1898 2706 1902
rect 2710 1898 2714 1902
rect 2710 1858 2714 1862
rect 2582 1838 2586 1842
rect 2630 1838 2634 1842
rect 2654 1838 2658 1842
rect 2686 1838 2690 1842
rect 2702 1828 2706 1832
rect 2574 1818 2578 1822
rect 2542 1808 2546 1812
rect 2670 1808 2674 1812
rect 2622 1798 2626 1802
rect 2710 1788 2714 1792
rect 2502 1778 2506 1782
rect 2550 1778 2554 1782
rect 2598 1778 2602 1782
rect 2534 1768 2538 1772
rect 2358 1728 2362 1732
rect 2446 1728 2450 1732
rect 2646 1768 2650 1772
rect 2606 1758 2610 1762
rect 2638 1758 2642 1762
rect 2678 1758 2682 1762
rect 2598 1748 2602 1752
rect 2550 1738 2554 1742
rect 2574 1738 2578 1742
rect 2518 1718 2522 1722
rect 2590 1718 2594 1722
rect 2526 1708 2530 1712
rect 2534 1708 2538 1712
rect 2598 1708 2602 1712
rect 2494 1688 2498 1692
rect 2366 1668 2370 1672
rect 2390 1668 2394 1672
rect 2278 1658 2282 1662
rect 2294 1658 2298 1662
rect 2326 1658 2330 1662
rect 2342 1658 2346 1662
rect 2262 1638 2266 1642
rect 2278 1598 2282 1602
rect 2286 1558 2290 1562
rect 2350 1578 2354 1582
rect 2342 1548 2346 1552
rect 2254 1538 2258 1542
rect 2318 1538 2322 1542
rect 2238 1498 2242 1502
rect 2246 1498 2250 1502
rect 2238 1488 2242 1492
rect 2246 1478 2250 1482
rect 2230 1458 2234 1462
rect 2214 1428 2218 1432
rect 2238 1428 2242 1432
rect 2246 1428 2250 1432
rect 2286 1518 2290 1522
rect 2262 1508 2266 1512
rect 2318 1508 2322 1512
rect 2278 1488 2282 1492
rect 2270 1478 2274 1482
rect 2310 1478 2314 1482
rect 2302 1458 2306 1462
rect 2294 1448 2298 1452
rect 2286 1428 2290 1432
rect 2246 1418 2250 1422
rect 2254 1418 2258 1422
rect 2302 1418 2306 1422
rect 2222 1398 2226 1402
rect 2198 1378 2202 1382
rect 2166 1368 2170 1372
rect 2174 1368 2178 1372
rect 2198 1368 2202 1372
rect 2214 1368 2218 1372
rect 2198 1358 2202 1362
rect 2190 1338 2194 1342
rect 2182 1308 2186 1312
rect 2150 1298 2154 1302
rect 2190 1278 2194 1282
rect 2134 1258 2138 1262
rect 2150 1248 2154 1252
rect 2174 1248 2178 1252
rect 2182 1168 2186 1172
rect 2110 1158 2114 1162
rect 2174 1138 2178 1142
rect 2078 1118 2082 1122
rect 2150 1128 2154 1132
rect 2134 1108 2138 1112
rect 2158 1108 2162 1112
rect 2166 1098 2170 1102
rect 2094 1088 2098 1092
rect 2142 1078 2146 1082
rect 2118 1048 2122 1052
rect 2126 1038 2130 1042
rect 2126 1018 2130 1022
rect 2070 1008 2074 1012
rect 2150 1048 2154 1052
rect 2054 988 2058 992
rect 2070 988 2074 992
rect 1998 968 2002 972
rect 2006 968 2010 972
rect 2030 968 2034 972
rect 2046 968 2050 972
rect 2054 968 2058 972
rect 1974 948 1978 952
rect 1990 948 1994 952
rect 1910 938 1914 942
rect 1874 903 1878 907
rect 1881 903 1885 907
rect 1862 888 1866 892
rect 1982 928 1986 932
rect 2102 978 2106 982
rect 2094 968 2098 972
rect 2134 968 2138 972
rect 2070 958 2074 962
rect 2118 958 2122 962
rect 2022 948 2026 952
rect 2038 938 2042 942
rect 1990 898 1994 902
rect 2006 898 2010 902
rect 1918 868 1922 872
rect 1950 868 1954 872
rect 1982 868 1986 872
rect 1878 859 1882 863
rect 1958 858 1962 862
rect 1974 858 1978 862
rect 1854 818 1858 822
rect 1926 818 1930 822
rect 1886 758 1890 762
rect 1846 748 1850 752
rect 1854 748 1858 752
rect 1798 698 1802 702
rect 1790 678 1794 682
rect 1806 658 1810 662
rect 1662 648 1666 652
rect 1726 648 1730 652
rect 1702 638 1706 642
rect 1798 638 1802 642
rect 1630 628 1634 632
rect 1678 588 1682 592
rect 1718 578 1722 582
rect 1614 568 1618 572
rect 1654 568 1658 572
rect 1606 558 1610 562
rect 1598 548 1602 552
rect 1614 548 1618 552
rect 1606 538 1610 542
rect 1622 508 1626 512
rect 1566 438 1570 442
rect 1614 428 1618 432
rect 1606 408 1610 412
rect 1438 378 1442 382
rect 1510 378 1514 382
rect 1470 368 1474 372
rect 1534 358 1538 362
rect 1526 348 1530 352
rect 1542 348 1546 352
rect 1598 348 1602 352
rect 1638 558 1642 562
rect 1702 558 1706 562
rect 1686 548 1690 552
rect 1678 538 1682 542
rect 1662 518 1666 522
rect 1630 488 1634 492
rect 1654 488 1658 492
rect 1670 478 1674 482
rect 1694 478 1698 482
rect 1630 468 1634 472
rect 1766 588 1770 592
rect 1798 598 1802 602
rect 1782 578 1786 582
rect 1790 568 1794 572
rect 1790 518 1794 522
rect 1742 508 1746 512
rect 1726 498 1730 502
rect 1734 488 1738 492
rect 1742 478 1746 482
rect 1766 478 1770 482
rect 1718 468 1722 472
rect 1790 468 1794 472
rect 1662 448 1666 452
rect 1662 428 1666 432
rect 1662 418 1666 422
rect 1638 398 1642 402
rect 1622 368 1626 372
rect 1670 388 1674 392
rect 1646 348 1650 352
rect 1702 378 1706 382
rect 1702 358 1706 362
rect 1734 398 1738 402
rect 1766 398 1770 402
rect 1790 378 1794 382
rect 1790 358 1794 362
rect 1326 338 1330 342
rect 1350 338 1354 342
rect 1614 338 1618 342
rect 1278 288 1282 292
rect 1294 288 1298 292
rect 1238 268 1242 272
rect 1278 268 1282 272
rect 1310 268 1314 272
rect 1134 258 1138 262
rect 1302 258 1306 262
rect 1166 248 1170 252
rect 1214 248 1218 252
rect 1310 248 1314 252
rect 1086 238 1090 242
rect 1110 238 1114 242
rect 1102 218 1106 222
rect 1102 168 1106 172
rect 1342 328 1346 332
rect 1470 308 1474 312
rect 1438 298 1442 302
rect 1430 288 1434 292
rect 1382 278 1386 282
rect 1398 278 1402 282
rect 1334 268 1338 272
rect 1318 188 1322 192
rect 1318 178 1322 182
rect 1222 168 1226 172
rect 1278 158 1282 162
rect 1030 148 1034 152
rect 1062 148 1066 152
rect 1246 148 1250 152
rect 1038 128 1042 132
rect 1030 88 1034 92
rect 1078 138 1082 142
rect 1062 128 1066 132
rect 1078 128 1082 132
rect 1078 118 1082 122
rect 1062 98 1066 102
rect 1182 138 1186 142
rect 1118 118 1122 122
rect 1110 78 1114 82
rect 1046 68 1050 72
rect 1102 68 1106 72
rect 1238 138 1242 142
rect 1254 118 1258 122
rect 1222 108 1226 112
rect 1214 98 1218 102
rect 1206 78 1210 82
rect 1454 258 1458 262
rect 1374 248 1378 252
rect 1354 203 1358 207
rect 1361 203 1365 207
rect 1326 168 1330 172
rect 1462 168 1466 172
rect 1342 158 1346 162
rect 1478 278 1482 282
rect 1542 328 1546 332
rect 1574 328 1578 332
rect 1582 328 1586 332
rect 1510 318 1514 322
rect 1670 308 1674 312
rect 1518 298 1522 302
rect 1534 298 1538 302
rect 1622 298 1626 302
rect 1494 288 1498 292
rect 1582 288 1586 292
rect 1590 288 1594 292
rect 1486 268 1490 272
rect 1662 278 1666 282
rect 1542 268 1546 272
rect 1518 248 1522 252
rect 1494 238 1498 242
rect 1534 238 1538 242
rect 1534 168 1538 172
rect 1510 158 1514 162
rect 1470 148 1474 152
rect 1494 148 1498 152
rect 1358 138 1362 142
rect 1270 88 1274 92
rect 1310 88 1314 92
rect 1350 88 1354 92
rect 1326 68 1330 72
rect 1014 58 1018 62
rect 1022 58 1026 62
rect 1038 58 1042 62
rect 1174 58 1178 62
rect 1238 58 1242 62
rect 1262 59 1266 63
rect 894 48 898 52
rect 1190 48 1194 52
rect 1334 48 1338 52
rect 1398 128 1402 132
rect 1374 118 1378 122
rect 1582 258 1586 262
rect 1598 258 1602 262
rect 1566 228 1570 232
rect 1750 308 1754 312
rect 1726 288 1730 292
rect 1742 278 1746 282
rect 1726 268 1730 272
rect 1822 668 1826 672
rect 1862 728 1866 732
rect 1958 728 1962 732
rect 1854 708 1858 712
rect 1902 708 1906 712
rect 1846 688 1850 692
rect 1846 668 1850 672
rect 1874 703 1878 707
rect 1881 703 1885 707
rect 1958 698 1962 702
rect 1926 668 1930 672
rect 1966 668 1970 672
rect 1902 618 1906 622
rect 1910 618 1914 622
rect 1878 578 1882 582
rect 1870 558 1874 562
rect 1806 548 1810 552
rect 1830 548 1834 552
rect 1782 338 1786 342
rect 1798 328 1802 332
rect 1798 318 1802 322
rect 1774 298 1778 302
rect 1782 288 1786 292
rect 1766 278 1770 282
rect 1766 268 1770 272
rect 1838 538 1842 542
rect 1958 648 1962 652
rect 1942 608 1946 612
rect 1934 588 1938 592
rect 1910 568 1914 572
rect 1958 568 1962 572
rect 1958 558 1962 562
rect 1894 528 1898 532
rect 1926 528 1930 532
rect 1862 518 1866 522
rect 1822 498 1826 502
rect 1822 488 1826 492
rect 1874 503 1878 507
rect 1881 503 1885 507
rect 1870 478 1874 482
rect 1822 468 1826 472
rect 1926 488 1930 492
rect 1902 468 1906 472
rect 1926 458 1930 462
rect 1942 458 1946 462
rect 1862 448 1866 452
rect 1894 448 1898 452
rect 1966 508 1970 512
rect 1918 438 1922 442
rect 1950 438 1954 442
rect 1918 428 1922 432
rect 1878 408 1882 412
rect 1862 398 1866 402
rect 1854 388 1858 392
rect 1830 368 1834 372
rect 1814 358 1818 362
rect 1814 348 1818 352
rect 1822 338 1826 342
rect 1854 318 1858 322
rect 1838 288 1842 292
rect 1806 278 1810 282
rect 1742 258 1746 262
rect 1638 248 1642 252
rect 1574 218 1578 222
rect 1630 218 1634 222
rect 1670 218 1674 222
rect 1486 128 1490 132
rect 1518 128 1522 132
rect 1534 128 1538 132
rect 1486 118 1490 122
rect 1462 98 1466 102
rect 1422 88 1426 92
rect 1382 78 1386 82
rect 1582 128 1586 132
rect 1566 98 1570 102
rect 1542 68 1546 72
rect 1622 78 1626 82
rect 1694 208 1698 212
rect 1678 198 1682 202
rect 1654 148 1658 152
rect 1662 128 1666 132
rect 1646 98 1650 102
rect 1670 78 1674 82
rect 1702 178 1706 182
rect 1878 358 1882 362
rect 1982 838 1986 842
rect 1990 788 1994 792
rect 1982 778 1986 782
rect 2046 928 2050 932
rect 2054 898 2058 902
rect 2062 798 2066 802
rect 2038 768 2042 772
rect 2022 758 2026 762
rect 1998 748 2002 752
rect 1990 698 1994 702
rect 1982 558 1986 562
rect 1990 548 1994 552
rect 2030 748 2034 752
rect 2046 738 2050 742
rect 2006 718 2010 722
rect 2086 938 2090 942
rect 2110 938 2114 942
rect 2078 928 2082 932
rect 2078 888 2082 892
rect 2086 878 2090 882
rect 2182 918 2186 922
rect 2118 908 2122 912
rect 2182 908 2186 912
rect 2110 868 2114 872
rect 2086 748 2090 752
rect 2078 738 2082 742
rect 2094 738 2098 742
rect 2006 688 2010 692
rect 2070 678 2074 682
rect 2086 678 2090 682
rect 2046 658 2050 662
rect 2022 648 2026 652
rect 2038 608 2042 612
rect 2062 608 2066 612
rect 2198 1218 2202 1222
rect 2198 1148 2202 1152
rect 2198 1098 2202 1102
rect 2214 1098 2218 1102
rect 2238 1358 2242 1362
rect 2230 1338 2234 1342
rect 2238 1278 2242 1282
rect 2294 1398 2298 1402
rect 2262 1358 2266 1362
rect 2262 1338 2266 1342
rect 2286 1338 2290 1342
rect 2286 1308 2290 1312
rect 2510 1678 2514 1682
rect 2470 1658 2474 1662
rect 2478 1658 2482 1662
rect 2422 1608 2426 1612
rect 2386 1603 2390 1607
rect 2393 1603 2397 1607
rect 2398 1578 2402 1582
rect 2526 1648 2530 1652
rect 2462 1628 2466 1632
rect 2454 1588 2458 1592
rect 2462 1578 2466 1582
rect 2502 1578 2506 1582
rect 2446 1558 2450 1562
rect 2430 1548 2434 1552
rect 2406 1528 2410 1532
rect 2430 1518 2434 1522
rect 2390 1458 2394 1462
rect 2326 1448 2330 1452
rect 2342 1448 2346 1452
rect 2350 1408 2354 1412
rect 2310 1398 2314 1402
rect 2386 1403 2390 1407
rect 2393 1403 2397 1407
rect 2318 1358 2322 1362
rect 2326 1358 2330 1362
rect 2430 1488 2434 1492
rect 2430 1458 2434 1462
rect 2462 1528 2466 1532
rect 2598 1668 2602 1672
rect 2566 1568 2570 1572
rect 2494 1538 2498 1542
rect 2486 1508 2490 1512
rect 2462 1478 2466 1482
rect 2438 1438 2442 1442
rect 2446 1428 2450 1432
rect 2430 1418 2434 1422
rect 2542 1528 2546 1532
rect 2518 1518 2522 1522
rect 2742 2028 2746 2032
rect 2774 2028 2778 2032
rect 2734 1938 2738 1942
rect 2734 1908 2738 1912
rect 2806 2008 2810 2012
rect 2846 2048 2850 2052
rect 2846 2028 2850 2032
rect 2750 1968 2754 1972
rect 2790 1968 2794 1972
rect 2822 1978 2826 1982
rect 2782 1958 2786 1962
rect 2798 1958 2802 1962
rect 2806 1958 2810 1962
rect 2782 1948 2786 1952
rect 2814 1948 2818 1952
rect 2798 1928 2802 1932
rect 2814 1928 2818 1932
rect 2766 1918 2770 1922
rect 2782 1918 2786 1922
rect 2790 1888 2794 1892
rect 2750 1858 2754 1862
rect 2774 1848 2778 1852
rect 2766 1838 2770 1842
rect 2742 1788 2746 1792
rect 2766 1778 2770 1782
rect 2726 1758 2730 1762
rect 2838 1968 2842 1972
rect 3006 2148 3010 2152
rect 3214 2208 3218 2212
rect 3142 2178 3146 2182
rect 3150 2178 3154 2182
rect 3222 2178 3226 2182
rect 3126 2138 3130 2142
rect 2966 2118 2970 2122
rect 2918 2108 2922 2112
rect 2890 2103 2894 2107
rect 2897 2103 2901 2107
rect 3022 2108 3026 2112
rect 2958 2098 2962 2102
rect 2966 2088 2970 2092
rect 3046 2088 3050 2092
rect 2902 2078 2906 2082
rect 2870 2068 2874 2072
rect 2878 2068 2882 2072
rect 2926 2068 2930 2072
rect 3078 2118 3082 2122
rect 3118 2108 3122 2112
rect 3102 2088 3106 2092
rect 3102 2078 3106 2082
rect 2918 2058 2922 2062
rect 3246 2188 3250 2192
rect 3238 2158 3242 2162
rect 3238 2148 3242 2152
rect 3214 2138 3218 2142
rect 3182 2128 3186 2132
rect 3214 2128 3218 2132
rect 3174 2118 3178 2122
rect 3182 2108 3186 2112
rect 3166 2098 3170 2102
rect 3206 2088 3210 2092
rect 3190 2078 3194 2082
rect 3238 2118 3242 2122
rect 3222 2108 3226 2112
rect 3118 2058 3122 2062
rect 3166 2058 3170 2062
rect 3214 2058 3218 2062
rect 2926 2048 2930 2052
rect 2950 2048 2954 2052
rect 2958 2038 2962 2042
rect 2854 1998 2858 2002
rect 3134 2048 3138 2052
rect 3086 2038 3090 2042
rect 3150 2008 3154 2012
rect 3102 1998 3106 2002
rect 2934 1968 2938 1972
rect 3070 1968 3074 1972
rect 2918 1958 2922 1962
rect 3054 1958 3058 1962
rect 3078 1958 3082 1962
rect 3094 1958 3098 1962
rect 2934 1948 2938 1952
rect 2894 1938 2898 1942
rect 2846 1878 2850 1882
rect 2806 1868 2810 1872
rect 2822 1868 2826 1872
rect 2814 1858 2818 1862
rect 2902 1928 2906 1932
rect 2862 1908 2866 1912
rect 2870 1908 2874 1912
rect 2890 1903 2894 1907
rect 2897 1903 2901 1907
rect 3030 1948 3034 1952
rect 3062 1948 3066 1952
rect 2966 1938 2970 1942
rect 2918 1898 2922 1902
rect 2870 1878 2874 1882
rect 2974 1898 2978 1902
rect 2870 1848 2874 1852
rect 2878 1848 2882 1852
rect 2830 1838 2834 1842
rect 2854 1838 2858 1842
rect 2846 1828 2850 1832
rect 2814 1808 2818 1812
rect 2782 1758 2786 1762
rect 2942 1838 2946 1842
rect 2902 1788 2906 1792
rect 2966 1788 2970 1792
rect 3126 1988 3130 1992
rect 3158 1958 3162 1962
rect 3118 1948 3122 1952
rect 3070 1938 3074 1942
rect 3038 1878 3042 1882
rect 3046 1878 3050 1882
rect 2982 1868 2986 1872
rect 3030 1868 3034 1872
rect 2982 1858 2986 1862
rect 3022 1858 3026 1862
rect 2830 1768 2834 1772
rect 2974 1768 2978 1772
rect 2838 1758 2842 1762
rect 2862 1758 2866 1762
rect 2630 1738 2634 1742
rect 2742 1738 2746 1742
rect 2766 1738 2770 1742
rect 2614 1708 2618 1712
rect 2654 1688 2658 1692
rect 2694 1688 2698 1692
rect 2750 1678 2754 1682
rect 2622 1668 2626 1672
rect 2670 1668 2674 1672
rect 2726 1668 2730 1672
rect 2638 1658 2642 1662
rect 2654 1658 2658 1662
rect 2686 1658 2690 1662
rect 2646 1648 2650 1652
rect 2614 1628 2618 1632
rect 2630 1628 2634 1632
rect 2606 1588 2610 1592
rect 2582 1578 2586 1582
rect 2630 1578 2634 1582
rect 2590 1558 2594 1562
rect 2574 1538 2578 1542
rect 2574 1518 2578 1522
rect 2550 1508 2554 1512
rect 2494 1468 2498 1472
rect 2526 1468 2530 1472
rect 2542 1468 2546 1472
rect 2558 1468 2562 1472
rect 2462 1458 2466 1462
rect 2462 1398 2466 1402
rect 2454 1388 2458 1392
rect 2550 1458 2554 1462
rect 2510 1448 2514 1452
rect 2502 1408 2506 1412
rect 2550 1398 2554 1402
rect 2518 1378 2522 1382
rect 2542 1378 2546 1382
rect 2494 1368 2498 1372
rect 2478 1358 2482 1362
rect 2614 1528 2618 1532
rect 2598 1518 2602 1522
rect 2590 1488 2594 1492
rect 2598 1459 2602 1463
rect 2598 1448 2602 1452
rect 2566 1378 2570 1382
rect 2574 1378 2578 1382
rect 2590 1378 2594 1382
rect 2558 1368 2562 1372
rect 2422 1348 2426 1352
rect 2510 1348 2514 1352
rect 2526 1348 2530 1352
rect 2550 1348 2554 1352
rect 2334 1338 2338 1342
rect 2326 1328 2330 1332
rect 2310 1298 2314 1302
rect 2406 1338 2410 1342
rect 2342 1328 2346 1332
rect 2462 1328 2466 1332
rect 2462 1318 2466 1322
rect 2398 1298 2402 1302
rect 2406 1298 2410 1302
rect 2334 1288 2338 1292
rect 2446 1288 2450 1292
rect 2422 1278 2426 1282
rect 2446 1278 2450 1282
rect 2302 1258 2306 1262
rect 2382 1258 2386 1262
rect 2254 1248 2258 1252
rect 2238 1238 2242 1242
rect 2270 1248 2274 1252
rect 2326 1248 2330 1252
rect 2302 1238 2306 1242
rect 2342 1238 2346 1242
rect 2262 1208 2266 1212
rect 2326 1228 2330 1232
rect 2342 1218 2346 1222
rect 2326 1188 2330 1192
rect 2278 1168 2282 1172
rect 2302 1158 2306 1162
rect 2238 1148 2242 1152
rect 2270 1148 2274 1152
rect 2386 1203 2390 1207
rect 2393 1203 2397 1207
rect 2374 1188 2378 1192
rect 2366 1158 2370 1162
rect 2246 1128 2250 1132
rect 2270 1098 2274 1102
rect 2270 1058 2274 1062
rect 2214 1048 2218 1052
rect 2198 978 2202 982
rect 2246 948 2250 952
rect 2270 948 2274 952
rect 2262 938 2266 942
rect 2254 928 2258 932
rect 2270 928 2274 932
rect 2230 908 2234 912
rect 2222 878 2226 882
rect 2270 878 2274 882
rect 2214 868 2218 872
rect 2142 818 2146 822
rect 2134 798 2138 802
rect 2118 768 2122 772
rect 2126 768 2130 772
rect 2110 738 2114 742
rect 2102 648 2106 652
rect 2078 638 2082 642
rect 2110 638 2114 642
rect 2102 618 2106 622
rect 2070 578 2074 582
rect 2022 568 2026 572
rect 2046 558 2050 562
rect 2078 568 2082 572
rect 2094 568 2098 572
rect 2014 528 2018 532
rect 1998 518 2002 522
rect 2014 518 2018 522
rect 2022 498 2026 502
rect 2030 488 2034 492
rect 1990 478 1994 482
rect 2014 478 2018 482
rect 2006 468 2010 472
rect 1966 458 1970 462
rect 2022 458 2026 462
rect 1982 448 1986 452
rect 1958 408 1962 412
rect 1950 378 1954 382
rect 1926 358 1930 362
rect 1894 348 1898 352
rect 1910 348 1914 352
rect 1974 368 1978 372
rect 1934 338 1938 342
rect 1966 338 1970 342
rect 1870 328 1874 332
rect 1874 303 1878 307
rect 1881 303 1885 307
rect 1806 248 1810 252
rect 1830 238 1834 242
rect 1790 208 1794 212
rect 1742 168 1746 172
rect 1918 308 1922 312
rect 2094 558 2098 562
rect 2174 828 2178 832
rect 2158 768 2162 772
rect 2158 758 2162 762
rect 2270 868 2274 872
rect 2214 858 2218 862
rect 2190 848 2194 852
rect 2214 848 2218 852
rect 2238 848 2242 852
rect 2174 698 2178 702
rect 2182 698 2186 702
rect 2166 688 2170 692
rect 2142 668 2146 672
rect 2126 638 2130 642
rect 2134 558 2138 562
rect 2222 838 2226 842
rect 2286 1128 2290 1132
rect 2342 1098 2346 1102
rect 2326 1088 2330 1092
rect 2334 1068 2338 1072
rect 2574 1348 2578 1352
rect 2502 1338 2506 1342
rect 2494 1318 2498 1322
rect 2486 1308 2490 1312
rect 2454 1248 2458 1252
rect 2486 1258 2490 1262
rect 2478 1248 2482 1252
rect 2446 1208 2450 1212
rect 2462 1208 2466 1212
rect 2422 1198 2426 1202
rect 2414 1148 2418 1152
rect 2382 1098 2386 1102
rect 2494 1188 2498 1192
rect 2454 1168 2458 1172
rect 2486 1158 2490 1162
rect 2470 1148 2474 1152
rect 2454 1138 2458 1142
rect 2446 1088 2450 1092
rect 2430 1068 2434 1072
rect 2350 1058 2354 1062
rect 2326 1038 2330 1042
rect 2414 1058 2418 1062
rect 2382 1048 2386 1052
rect 2422 1048 2426 1052
rect 2462 1048 2466 1052
rect 2358 1038 2362 1042
rect 2334 958 2338 962
rect 2294 948 2298 952
rect 2326 938 2330 942
rect 2334 938 2338 942
rect 2386 1003 2390 1007
rect 2393 1003 2397 1007
rect 2430 958 2434 962
rect 2374 948 2378 952
rect 2542 1328 2546 1332
rect 2558 1328 2562 1332
rect 2526 1288 2530 1292
rect 2582 1318 2586 1322
rect 2614 1368 2618 1372
rect 2614 1348 2618 1352
rect 2678 1568 2682 1572
rect 2646 1548 2650 1552
rect 2774 1638 2778 1642
rect 2774 1598 2778 1602
rect 2750 1588 2754 1592
rect 2654 1508 2658 1512
rect 2654 1468 2658 1472
rect 2710 1528 2714 1532
rect 2710 1518 2714 1522
rect 2726 1518 2730 1522
rect 2742 1518 2746 1522
rect 2694 1488 2698 1492
rect 2702 1478 2706 1482
rect 2726 1478 2730 1482
rect 2694 1468 2698 1472
rect 2686 1418 2690 1422
rect 2670 1398 2674 1402
rect 2670 1338 2674 1342
rect 2614 1318 2618 1322
rect 2638 1318 2642 1322
rect 2806 1728 2810 1732
rect 2790 1718 2794 1722
rect 2918 1748 2922 1752
rect 2990 1758 2994 1762
rect 2830 1738 2834 1742
rect 2926 1738 2930 1742
rect 2958 1738 2962 1742
rect 2890 1703 2894 1707
rect 2897 1703 2901 1707
rect 2814 1698 2818 1702
rect 2814 1688 2818 1692
rect 2934 1688 2938 1692
rect 2806 1668 2810 1672
rect 2830 1678 2834 1682
rect 2854 1678 2858 1682
rect 2886 1678 2890 1682
rect 2814 1638 2818 1642
rect 2878 1668 2882 1672
rect 2838 1658 2842 1662
rect 2854 1658 2858 1662
rect 2902 1658 2906 1662
rect 2862 1628 2866 1632
rect 2846 1608 2850 1612
rect 2910 1598 2914 1602
rect 2878 1588 2882 1592
rect 2902 1588 2906 1592
rect 2822 1568 2826 1572
rect 2846 1568 2850 1572
rect 2782 1548 2786 1552
rect 2854 1548 2858 1552
rect 2790 1538 2794 1542
rect 2790 1518 2794 1522
rect 2822 1528 2826 1532
rect 2870 1528 2874 1532
rect 2902 1528 2906 1532
rect 2806 1498 2810 1502
rect 2750 1458 2754 1462
rect 2774 1458 2778 1462
rect 2766 1438 2770 1442
rect 2806 1438 2810 1442
rect 2766 1398 2770 1402
rect 2742 1388 2746 1392
rect 2734 1348 2738 1352
rect 2726 1338 2730 1342
rect 2734 1328 2738 1332
rect 2734 1298 2738 1302
rect 2702 1278 2706 1282
rect 2798 1348 2802 1352
rect 2782 1318 2786 1322
rect 2694 1268 2698 1272
rect 2526 1258 2530 1262
rect 2550 1258 2554 1262
rect 2566 1258 2570 1262
rect 2798 1278 2802 1282
rect 2890 1503 2894 1507
rect 2897 1503 2901 1507
rect 3006 1838 3010 1842
rect 3022 1838 3026 1842
rect 3006 1778 3010 1782
rect 3006 1748 3010 1752
rect 2982 1718 2986 1722
rect 2998 1718 3002 1722
rect 2974 1668 2978 1672
rect 2942 1578 2946 1582
rect 2958 1578 2962 1582
rect 2934 1568 2938 1572
rect 2926 1548 2930 1552
rect 2934 1548 2938 1552
rect 3062 1908 3066 1912
rect 3110 1928 3114 1932
rect 3094 1918 3098 1922
rect 3150 1928 3154 1932
rect 3142 1918 3146 1922
rect 3102 1888 3106 1892
rect 3158 1888 3162 1892
rect 3134 1878 3138 1882
rect 3038 1848 3042 1852
rect 3038 1838 3042 1842
rect 3078 1858 3082 1862
rect 3094 1858 3098 1862
rect 3070 1818 3074 1822
rect 3054 1798 3058 1802
rect 3078 1798 3082 1802
rect 3070 1788 3074 1792
rect 3038 1768 3042 1772
rect 3046 1748 3050 1752
rect 3062 1748 3066 1752
rect 3022 1718 3026 1722
rect 2990 1608 2994 1612
rect 2982 1548 2986 1552
rect 3046 1728 3050 1732
rect 3030 1698 3034 1702
rect 3038 1698 3042 1702
rect 3006 1638 3010 1642
rect 3014 1598 3018 1602
rect 3070 1688 3074 1692
rect 3070 1668 3074 1672
rect 3102 1778 3106 1782
rect 3086 1738 3090 1742
rect 3110 1728 3114 1732
rect 3150 1868 3154 1872
rect 3206 2048 3210 2052
rect 3246 2098 3250 2102
rect 3270 2248 3274 2252
rect 3270 2218 3274 2222
rect 3262 2188 3266 2192
rect 3254 2088 3258 2092
rect 3238 2058 3242 2062
rect 3254 2048 3258 2052
rect 3174 2038 3178 2042
rect 3198 2018 3202 2022
rect 3182 1958 3186 1962
rect 3190 1958 3194 1962
rect 3198 1938 3202 1942
rect 3182 1898 3186 1902
rect 3238 1988 3242 1992
rect 3350 2308 3354 2312
rect 3374 2308 3378 2312
rect 3334 2288 3338 2292
rect 3310 2268 3314 2272
rect 3326 2238 3330 2242
rect 3302 2208 3306 2212
rect 3398 2328 3402 2332
rect 3398 2298 3402 2302
rect 3406 2298 3410 2302
rect 3422 2358 3426 2362
rect 3502 2448 3506 2452
rect 3510 2438 3514 2442
rect 3518 2418 3522 2422
rect 3478 2398 3482 2402
rect 3494 2368 3498 2372
rect 3510 2368 3514 2372
rect 3614 2508 3618 2512
rect 3606 2478 3610 2482
rect 3582 2468 3586 2472
rect 3558 2438 3562 2442
rect 3526 2398 3530 2402
rect 3526 2368 3530 2372
rect 3542 2368 3546 2372
rect 3430 2348 3434 2352
rect 3446 2348 3450 2352
rect 3462 2348 3466 2352
rect 3518 2348 3522 2352
rect 3550 2348 3554 2352
rect 3526 2338 3530 2342
rect 3478 2318 3482 2322
rect 3494 2318 3498 2322
rect 3526 2318 3530 2322
rect 3430 2308 3434 2312
rect 3446 2308 3450 2312
rect 3502 2308 3506 2312
rect 3382 2288 3386 2292
rect 3462 2288 3466 2292
rect 3478 2288 3482 2292
rect 3494 2288 3498 2292
rect 3422 2266 3426 2270
rect 3446 2268 3450 2272
rect 3478 2268 3482 2272
rect 3494 2268 3498 2272
rect 3382 2248 3386 2252
rect 3402 2203 3406 2207
rect 3409 2203 3413 2207
rect 3534 2278 3538 2282
rect 3510 2268 3514 2272
rect 3518 2268 3522 2272
rect 3622 2458 3626 2462
rect 3678 2528 3682 2532
rect 3654 2498 3658 2502
rect 3654 2468 3658 2472
rect 3646 2448 3650 2452
rect 3598 2438 3602 2442
rect 3582 2428 3586 2432
rect 3582 2408 3586 2412
rect 3606 2408 3610 2412
rect 3590 2378 3594 2382
rect 3574 2358 3578 2362
rect 3566 2288 3570 2292
rect 3598 2278 3602 2282
rect 3582 2268 3586 2272
rect 3590 2268 3594 2272
rect 3550 2248 3554 2252
rect 3558 2248 3562 2252
rect 3470 2218 3474 2222
rect 3550 2238 3554 2242
rect 3526 2208 3530 2212
rect 3438 2198 3442 2202
rect 3438 2178 3442 2182
rect 3278 2168 3282 2172
rect 3390 2168 3394 2172
rect 3470 2168 3474 2172
rect 3534 2168 3538 2172
rect 3302 2158 3306 2162
rect 3358 2158 3362 2162
rect 3382 2158 3386 2162
rect 3318 2148 3322 2152
rect 3278 2138 3282 2142
rect 3294 2138 3298 2142
rect 3350 2138 3354 2142
rect 3358 2098 3362 2102
rect 3286 2088 3290 2092
rect 3350 2088 3354 2092
rect 3326 2058 3330 2062
rect 3278 2008 3282 2012
rect 3262 1968 3266 1972
rect 3222 1958 3226 1962
rect 3270 1938 3274 1942
rect 3294 2048 3298 2052
rect 3294 1998 3298 2002
rect 3366 2088 3370 2092
rect 3342 2058 3346 2062
rect 3542 2148 3546 2152
rect 3494 2138 3498 2142
rect 3398 2108 3402 2112
rect 3454 2098 3458 2102
rect 3390 2088 3394 2092
rect 3518 2078 3522 2082
rect 3574 2218 3578 2222
rect 3582 2218 3586 2222
rect 3598 2168 3602 2172
rect 3414 2068 3418 2072
rect 3462 2068 3466 2072
rect 3406 2058 3410 2062
rect 3454 2058 3458 2062
rect 3478 2058 3482 2062
rect 3550 2058 3554 2062
rect 3382 2048 3386 2052
rect 3374 2038 3378 2042
rect 3334 2018 3338 2022
rect 3402 2003 3406 2007
rect 3409 2003 3413 2007
rect 3318 1978 3322 1982
rect 3438 1978 3442 1982
rect 3430 1968 3434 1972
rect 3286 1928 3290 1932
rect 3230 1908 3234 1912
rect 3278 1908 3282 1912
rect 3438 1948 3442 1952
rect 3366 1938 3370 1942
rect 3422 1938 3426 1942
rect 3446 1938 3450 1942
rect 3462 1928 3466 1932
rect 3310 1918 3314 1922
rect 3294 1898 3298 1902
rect 3262 1888 3266 1892
rect 3294 1888 3298 1892
rect 3510 2048 3514 2052
rect 3502 2028 3506 2032
rect 3398 1918 3402 1922
rect 3470 1918 3474 1922
rect 3494 1918 3498 1922
rect 3454 1908 3458 1912
rect 3366 1878 3370 1882
rect 3190 1868 3194 1872
rect 3166 1858 3170 1862
rect 3222 1858 3226 1862
rect 3238 1858 3242 1862
rect 3262 1868 3266 1872
rect 3326 1868 3330 1872
rect 3270 1858 3274 1862
rect 3126 1818 3130 1822
rect 3142 1818 3146 1822
rect 3126 1808 3130 1812
rect 3142 1758 3146 1762
rect 3182 1848 3186 1852
rect 3214 1848 3218 1852
rect 3182 1818 3186 1822
rect 3238 1798 3242 1802
rect 3198 1788 3202 1792
rect 3182 1758 3186 1762
rect 3126 1748 3130 1752
rect 3134 1738 3138 1742
rect 3174 1738 3178 1742
rect 3158 1698 3162 1702
rect 3118 1688 3122 1692
rect 3150 1688 3154 1692
rect 3094 1678 3098 1682
rect 3126 1678 3130 1682
rect 3142 1678 3146 1682
rect 3086 1668 3090 1672
rect 3238 1738 3242 1742
rect 3254 1738 3258 1742
rect 3206 1718 3210 1722
rect 3222 1688 3226 1692
rect 3174 1668 3178 1672
rect 3214 1668 3218 1672
rect 3046 1658 3050 1662
rect 3078 1658 3082 1662
rect 3142 1658 3146 1662
rect 3038 1648 3042 1652
rect 3102 1648 3106 1652
rect 3190 1648 3194 1652
rect 3054 1638 3058 1642
rect 3118 1588 3122 1592
rect 3022 1578 3026 1582
rect 3078 1578 3082 1582
rect 3110 1578 3114 1582
rect 3046 1568 3050 1572
rect 3070 1568 3074 1572
rect 2974 1538 2978 1542
rect 2990 1538 2994 1542
rect 2990 1528 2994 1532
rect 2934 1518 2938 1522
rect 2934 1508 2938 1512
rect 2886 1458 2890 1462
rect 2894 1448 2898 1452
rect 2862 1438 2866 1442
rect 2878 1438 2882 1442
rect 2878 1428 2882 1432
rect 2878 1408 2882 1412
rect 2870 1308 2874 1312
rect 2894 1328 2898 1332
rect 2950 1468 2954 1472
rect 2942 1448 2946 1452
rect 2926 1418 2930 1422
rect 2918 1318 2922 1322
rect 2890 1303 2894 1307
rect 2897 1303 2901 1307
rect 2798 1268 2802 1272
rect 2830 1268 2834 1272
rect 2854 1268 2858 1272
rect 2646 1258 2650 1262
rect 2718 1258 2722 1262
rect 2734 1258 2738 1262
rect 2758 1258 2762 1262
rect 2766 1258 2770 1262
rect 2854 1258 2858 1262
rect 2870 1258 2874 1262
rect 2910 1258 2914 1262
rect 2598 1248 2602 1252
rect 2710 1248 2714 1252
rect 2566 1218 2570 1222
rect 2542 1188 2546 1192
rect 2670 1188 2674 1192
rect 2590 1178 2594 1182
rect 2550 1168 2554 1172
rect 2518 1148 2522 1152
rect 2566 1158 2570 1162
rect 2582 1148 2586 1152
rect 2606 1138 2610 1142
rect 2654 1138 2658 1142
rect 2502 1098 2506 1102
rect 2518 1078 2522 1082
rect 2526 1078 2530 1082
rect 2494 1068 2498 1072
rect 2478 948 2482 952
rect 2358 918 2362 922
rect 2302 908 2306 912
rect 2350 908 2354 912
rect 2358 898 2362 902
rect 2350 868 2354 872
rect 2286 838 2290 842
rect 2326 838 2330 842
rect 2214 768 2218 772
rect 2278 758 2282 762
rect 2342 828 2346 832
rect 2294 798 2298 802
rect 2238 748 2242 752
rect 2246 748 2250 752
rect 2254 748 2258 752
rect 2302 768 2306 772
rect 2446 938 2450 942
rect 2462 938 2466 942
rect 2406 928 2410 932
rect 2430 878 2434 882
rect 2446 868 2450 872
rect 2382 858 2386 862
rect 2398 858 2402 862
rect 2390 838 2394 842
rect 2422 818 2426 822
rect 2414 808 2418 812
rect 2386 803 2390 807
rect 2393 803 2397 807
rect 2398 778 2402 782
rect 2326 758 2330 762
rect 2310 748 2314 752
rect 2334 748 2338 752
rect 2262 738 2266 742
rect 2270 738 2274 742
rect 2278 738 2282 742
rect 2294 738 2298 742
rect 2230 688 2234 692
rect 2190 678 2194 682
rect 2222 668 2226 672
rect 2214 658 2218 662
rect 2262 698 2266 702
rect 2278 678 2282 682
rect 2254 668 2258 672
rect 2270 658 2274 662
rect 2206 638 2210 642
rect 2238 638 2242 642
rect 2246 638 2250 642
rect 2222 628 2226 632
rect 2510 948 2514 952
rect 2470 878 2474 882
rect 2454 848 2458 852
rect 2430 768 2434 772
rect 2446 758 2450 762
rect 2414 748 2418 752
rect 2358 738 2362 742
rect 2358 718 2362 722
rect 2366 678 2370 682
rect 2342 658 2346 662
rect 2182 558 2186 562
rect 2238 558 2242 562
rect 2278 558 2282 562
rect 2150 538 2154 542
rect 2166 538 2170 542
rect 2102 528 2106 532
rect 2046 518 2050 522
rect 2086 518 2090 522
rect 2110 518 2114 522
rect 2038 398 2042 402
rect 2038 378 2042 382
rect 2038 338 2042 342
rect 2102 508 2106 512
rect 2166 508 2170 512
rect 2054 478 2058 482
rect 2070 478 2074 482
rect 2054 468 2058 472
rect 2070 468 2074 472
rect 2086 448 2090 452
rect 2070 438 2074 442
rect 2070 418 2074 422
rect 2086 368 2090 372
rect 2150 498 2154 502
rect 2110 478 2114 482
rect 2134 458 2138 462
rect 2142 448 2146 452
rect 2118 428 2122 432
rect 2142 428 2146 432
rect 2102 418 2106 422
rect 2054 338 2058 342
rect 2094 338 2098 342
rect 1998 328 2002 332
rect 2030 328 2034 332
rect 2046 328 2050 332
rect 2062 328 2066 332
rect 2022 318 2026 322
rect 2094 318 2098 322
rect 2118 348 2122 352
rect 2134 348 2138 352
rect 1998 298 2002 302
rect 2102 298 2106 302
rect 2126 308 2130 312
rect 2126 298 2130 302
rect 2286 538 2290 542
rect 2262 518 2266 522
rect 2182 498 2186 502
rect 2174 488 2178 492
rect 2342 648 2346 652
rect 2302 568 2306 572
rect 2398 718 2402 722
rect 2438 698 2442 702
rect 2462 838 2466 842
rect 2438 678 2442 682
rect 2414 668 2418 672
rect 2454 668 2458 672
rect 2406 648 2410 652
rect 2406 638 2410 642
rect 2382 618 2386 622
rect 2386 603 2390 607
rect 2393 603 2397 607
rect 2430 598 2434 602
rect 2446 588 2450 592
rect 2390 558 2394 562
rect 2438 558 2442 562
rect 2302 538 2306 542
rect 2334 538 2338 542
rect 2366 538 2370 542
rect 2358 528 2362 532
rect 2318 518 2322 522
rect 2294 508 2298 512
rect 2318 508 2322 512
rect 2278 498 2282 502
rect 2310 488 2314 492
rect 2294 468 2298 472
rect 2158 458 2162 462
rect 2238 459 2242 463
rect 2166 408 2170 412
rect 2174 408 2178 412
rect 2206 408 2210 412
rect 2158 338 2162 342
rect 2150 298 2154 302
rect 2174 368 2178 372
rect 2214 368 2218 372
rect 2246 368 2250 372
rect 2182 358 2186 362
rect 2278 448 2282 452
rect 2286 438 2290 442
rect 2262 358 2266 362
rect 2310 358 2314 362
rect 2214 348 2218 352
rect 2286 348 2290 352
rect 2230 338 2234 342
rect 2262 338 2266 342
rect 2214 328 2218 332
rect 2246 328 2250 332
rect 2190 318 2194 322
rect 2182 298 2186 302
rect 2158 288 2162 292
rect 2166 278 2170 282
rect 1966 268 1970 272
rect 1982 268 1986 272
rect 2014 268 2018 272
rect 2110 268 2114 272
rect 1910 218 1914 222
rect 1886 208 1890 212
rect 1830 158 1834 162
rect 1894 168 1898 172
rect 1686 148 1690 152
rect 1766 147 1770 151
rect 1814 148 1818 152
rect 1854 148 1858 152
rect 1910 148 1914 152
rect 2006 258 2010 262
rect 2062 248 2066 252
rect 2062 218 2066 222
rect 2030 208 2034 212
rect 1982 198 1986 202
rect 1974 188 1978 192
rect 1998 188 2002 192
rect 2062 188 2066 192
rect 1974 168 1978 172
rect 2046 168 2050 172
rect 1942 158 1946 162
rect 2038 158 2042 162
rect 2022 148 2026 152
rect 1822 138 1826 142
rect 2030 138 2034 142
rect 1790 128 1794 132
rect 1686 118 1690 122
rect 1710 108 1714 112
rect 1806 108 1810 112
rect 1874 103 1878 107
rect 1881 103 1885 107
rect 1862 88 1866 92
rect 1646 68 1650 72
rect 1678 68 1682 72
rect 1750 68 1754 72
rect 1814 68 1818 72
rect 1398 58 1402 62
rect 1414 58 1418 62
rect 1630 58 1634 62
rect 1926 128 1930 132
rect 1910 88 1914 92
rect 1950 118 1954 122
rect 2014 108 2018 112
rect 2006 98 2010 102
rect 1974 78 1978 82
rect 2270 328 2274 332
rect 2230 278 2234 282
rect 2222 268 2226 272
rect 2102 208 2106 212
rect 2110 208 2114 212
rect 2094 168 2098 172
rect 2102 158 2106 162
rect 2174 248 2178 252
rect 2230 258 2234 262
rect 2214 248 2218 252
rect 2198 168 2202 172
rect 2310 338 2314 342
rect 2302 278 2306 282
rect 2254 258 2258 262
rect 2278 258 2282 262
rect 2246 248 2250 252
rect 2270 178 2274 182
rect 2326 468 2330 472
rect 2366 478 2370 482
rect 2430 528 2434 532
rect 2414 468 2418 472
rect 2334 458 2338 462
rect 2358 458 2362 462
rect 2334 448 2338 452
rect 2342 368 2346 372
rect 2358 358 2362 362
rect 2422 458 2426 462
rect 2422 448 2426 452
rect 2398 438 2402 442
rect 2430 438 2434 442
rect 2386 403 2390 407
rect 2393 403 2397 407
rect 2398 368 2402 372
rect 2382 358 2386 362
rect 2430 358 2434 362
rect 2374 348 2378 352
rect 2318 328 2322 332
rect 2318 258 2322 262
rect 2310 158 2314 162
rect 2086 148 2090 152
rect 2118 148 2122 152
rect 2238 148 2242 152
rect 2262 148 2266 152
rect 2286 148 2290 152
rect 2134 138 2138 142
rect 2190 138 2194 142
rect 2078 128 2082 132
rect 2062 108 2066 112
rect 2054 78 2058 82
rect 2150 98 2154 102
rect 2094 88 2098 92
rect 2110 88 2114 92
rect 2118 68 2122 72
rect 2142 68 2146 72
rect 2334 208 2338 212
rect 2366 178 2370 182
rect 2406 338 2410 342
rect 2382 318 2386 322
rect 2446 528 2450 532
rect 2518 938 2522 942
rect 2534 1058 2538 1062
rect 2662 1088 2666 1092
rect 2558 1078 2562 1082
rect 2574 1078 2578 1082
rect 2646 1078 2650 1082
rect 2654 1068 2658 1072
rect 2726 1168 2730 1172
rect 2726 1148 2730 1152
rect 2742 1138 2746 1142
rect 2710 1078 2714 1082
rect 2734 1068 2738 1072
rect 2750 1068 2754 1072
rect 2606 1058 2610 1062
rect 2678 1058 2682 1062
rect 2686 1058 2690 1062
rect 2718 1058 2722 1062
rect 2558 1048 2562 1052
rect 2670 1038 2674 1042
rect 2734 1038 2738 1042
rect 2782 1208 2786 1212
rect 2766 1168 2770 1172
rect 2846 1178 2850 1182
rect 2830 1168 2834 1172
rect 2806 1148 2810 1152
rect 2790 1128 2794 1132
rect 2774 1098 2778 1102
rect 2958 1398 2962 1402
rect 3030 1528 3034 1532
rect 3070 1528 3074 1532
rect 3046 1518 3050 1522
rect 3086 1548 3090 1552
rect 3126 1548 3130 1552
rect 3094 1538 3098 1542
rect 3086 1528 3090 1532
rect 3014 1508 3018 1512
rect 3078 1508 3082 1512
rect 2990 1498 2994 1502
rect 3030 1498 3034 1502
rect 2998 1478 3002 1482
rect 3014 1448 3018 1452
rect 2998 1438 3002 1442
rect 3110 1498 3114 1502
rect 3270 1668 3274 1672
rect 3254 1648 3258 1652
rect 3270 1648 3274 1652
rect 3198 1638 3202 1642
rect 3214 1638 3218 1642
rect 3230 1638 3234 1642
rect 3230 1628 3234 1632
rect 3222 1568 3226 1572
rect 3318 1758 3322 1762
rect 3374 1758 3378 1762
rect 3294 1748 3298 1752
rect 3326 1748 3330 1752
rect 3342 1748 3346 1752
rect 3526 2008 3530 2012
rect 3542 1978 3546 1982
rect 3614 2368 3618 2372
rect 3646 2368 3650 2372
rect 3630 2358 3634 2362
rect 3638 2348 3642 2352
rect 3622 2318 3626 2322
rect 3766 2958 3770 2962
rect 3798 2958 3802 2962
rect 3718 2948 3722 2952
rect 3742 2948 3746 2952
rect 3734 2888 3738 2892
rect 3782 2878 3786 2882
rect 3782 2868 3786 2872
rect 3910 3178 3914 3182
rect 3870 3068 3874 3072
rect 3910 3118 3914 3122
rect 3886 3078 3890 3082
rect 3886 3068 3890 3072
rect 3902 3068 3906 3072
rect 3894 3048 3898 3052
rect 3886 3038 3890 3042
rect 3878 3018 3882 3022
rect 3922 3103 3926 3107
rect 3929 3103 3933 3107
rect 3934 3088 3938 3092
rect 3862 2918 3866 2922
rect 3838 2908 3842 2912
rect 3854 2888 3858 2892
rect 3902 2878 3906 2882
rect 3750 2858 3754 2862
rect 3798 2858 3802 2862
rect 3830 2858 3834 2862
rect 3846 2858 3850 2862
rect 3782 2838 3786 2842
rect 3790 2818 3794 2822
rect 3846 2848 3850 2852
rect 3710 2758 3714 2762
rect 3766 2758 3770 2762
rect 3798 2758 3802 2762
rect 3806 2758 3810 2762
rect 3750 2728 3754 2732
rect 3806 2728 3810 2732
rect 3742 2708 3746 2712
rect 3718 2688 3722 2692
rect 3734 2668 3738 2672
rect 3702 2608 3706 2612
rect 3822 2698 3826 2702
rect 3750 2668 3754 2672
rect 3790 2668 3794 2672
rect 3814 2668 3818 2672
rect 3830 2678 3834 2682
rect 3926 2988 3930 2992
rect 3926 2958 3930 2962
rect 3990 3238 3994 3242
rect 4022 3238 4026 3242
rect 3958 3158 3962 3162
rect 3982 3098 3986 3102
rect 4110 3378 4114 3382
rect 4094 3368 4098 3372
rect 4110 3368 4114 3372
rect 4094 3348 4098 3352
rect 4078 3338 4082 3342
rect 4038 3328 4042 3332
rect 4046 3328 4050 3332
rect 4190 3578 4194 3582
rect 4182 3568 4186 3572
rect 4158 3558 4162 3562
rect 4302 3878 4306 3882
rect 4310 3878 4314 3882
rect 4334 3898 4338 3902
rect 4350 3958 4354 3962
rect 4374 3958 4378 3962
rect 4342 3858 4346 3862
rect 4294 3848 4298 3852
rect 4318 3848 4322 3852
rect 4278 3828 4282 3832
rect 4270 3758 4274 3762
rect 4262 3678 4266 3682
rect 4326 3758 4330 3762
rect 4342 3798 4346 3802
rect 4310 3728 4314 3732
rect 4334 3728 4338 3732
rect 4326 3718 4330 3722
rect 4318 3678 4322 3682
rect 4302 3668 4306 3672
rect 4326 3668 4330 3672
rect 4566 4058 4570 4062
rect 4486 4048 4490 4052
rect 4518 3968 4522 3972
rect 4486 3958 4490 3962
rect 4478 3948 4482 3952
rect 4502 3948 4506 3952
rect 4518 3948 4522 3952
rect 4446 3938 4450 3942
rect 4446 3908 4450 3912
rect 4398 3898 4402 3902
rect 4414 3878 4418 3882
rect 4422 3878 4426 3882
rect 4390 3858 4394 3862
rect 4430 3858 4434 3862
rect 4366 3848 4370 3852
rect 4382 3848 4386 3852
rect 4374 3828 4378 3832
rect 4358 3798 4362 3802
rect 4358 3758 4362 3762
rect 4374 3738 4378 3742
rect 4358 3718 4362 3722
rect 4426 3803 4430 3807
rect 4433 3803 4437 3807
rect 4398 3768 4402 3772
rect 4406 3758 4410 3762
rect 4550 3928 4554 3932
rect 4542 3908 4546 3912
rect 4502 3898 4506 3902
rect 4534 3898 4538 3902
rect 4494 3878 4498 3882
rect 4510 3878 4514 3882
rect 4686 4688 4690 4692
rect 4726 4718 4730 4722
rect 4742 4718 4746 4722
rect 4710 4698 4714 4702
rect 4718 4688 4722 4692
rect 4710 4658 4714 4662
rect 4694 4648 4698 4652
rect 4702 4648 4706 4652
rect 4718 4588 4722 4592
rect 4686 4558 4690 4562
rect 4734 4558 4738 4562
rect 4782 5058 4786 5062
rect 4782 5028 4786 5032
rect 4806 4968 4810 4972
rect 4806 4958 4810 4962
rect 4782 4948 4786 4952
rect 4798 4948 4802 4952
rect 4822 4948 4826 4952
rect 4790 4868 4794 4872
rect 4998 5058 5002 5062
rect 5022 5058 5026 5062
rect 5054 5058 5058 5062
rect 4902 5048 4906 5052
rect 4926 5048 4930 5052
rect 4982 5048 4986 5052
rect 5014 5048 5018 5052
rect 4966 5018 4970 5022
rect 4870 4958 4874 4962
rect 4918 4948 4922 4952
rect 4974 4948 4978 4952
rect 4862 4938 4866 4942
rect 4838 4908 4842 4912
rect 4966 4938 4970 4942
rect 4894 4918 4898 4922
rect 4938 4903 4942 4907
rect 4945 4903 4949 4907
rect 4974 4888 4978 4892
rect 4878 4878 4882 4882
rect 4974 4878 4978 4882
rect 4806 4868 4810 4872
rect 4894 4848 4898 4852
rect 4974 4848 4978 4852
rect 4798 4778 4802 4782
rect 4806 4758 4810 4762
rect 4774 4738 4778 4742
rect 4774 4718 4778 4722
rect 4758 4708 4762 4712
rect 4854 4688 4858 4692
rect 4910 4738 4914 4742
rect 5006 4968 5010 4972
rect 5014 4928 5018 4932
rect 5006 4918 5010 4922
rect 5022 4918 5026 4922
rect 4990 4818 4994 4822
rect 5038 4958 5042 4962
rect 5022 4888 5026 4892
rect 5030 4888 5034 4892
rect 5006 4868 5010 4872
rect 5014 4868 5018 4872
rect 4998 4808 5002 4812
rect 5014 4808 5018 4812
rect 5006 4778 5010 4782
rect 4998 4768 5002 4772
rect 5006 4768 5010 4772
rect 5030 4758 5034 4762
rect 4966 4728 4970 4732
rect 4990 4728 4994 4732
rect 4918 4718 4922 4722
rect 4938 4703 4942 4707
rect 4945 4703 4949 4707
rect 4902 4688 4906 4692
rect 4758 4668 4762 4672
rect 4966 4668 4970 4672
rect 4774 4658 4778 4662
rect 4862 4658 4866 4662
rect 4894 4658 4898 4662
rect 4694 4548 4698 4552
rect 4726 4548 4730 4552
rect 4758 4548 4762 4552
rect 4702 4538 4706 4542
rect 4726 4538 4730 4542
rect 4758 4538 4762 4542
rect 4702 4528 4706 4532
rect 4686 4508 4690 4512
rect 4686 4498 4690 4502
rect 4694 4488 4698 4492
rect 4726 4518 4730 4522
rect 4750 4518 4754 4522
rect 4782 4648 4786 4652
rect 4886 4648 4890 4652
rect 4902 4638 4906 4642
rect 4846 4618 4850 4622
rect 4814 4608 4818 4612
rect 4806 4578 4810 4582
rect 4990 4718 4994 4722
rect 4998 4698 5002 4702
rect 4982 4678 4986 4682
rect 4982 4648 4986 4652
rect 4974 4598 4978 4602
rect 4854 4568 4858 4572
rect 4838 4558 4842 4562
rect 4830 4548 4834 4552
rect 4774 4538 4778 4542
rect 4790 4538 4794 4542
rect 4718 4498 4722 4502
rect 4742 4508 4746 4512
rect 4790 4508 4794 4512
rect 4790 4498 4794 4502
rect 4974 4558 4978 4562
rect 4990 4558 4994 4562
rect 4846 4548 4850 4552
rect 4814 4478 4818 4482
rect 4758 4468 4762 4472
rect 4806 4458 4810 4462
rect 4862 4538 4866 4542
rect 4910 4538 4914 4542
rect 4862 4518 4866 4522
rect 4878 4518 4882 4522
rect 4854 4488 4858 4492
rect 4822 4458 4826 4462
rect 4862 4458 4866 4462
rect 4726 4448 4730 4452
rect 4830 4448 4834 4452
rect 4974 4518 4978 4522
rect 4938 4503 4942 4507
rect 4945 4503 4949 4507
rect 4902 4488 4906 4492
rect 4894 4468 4898 4472
rect 4942 4478 4946 4482
rect 4926 4468 4930 4472
rect 4902 4458 4906 4462
rect 4870 4408 4874 4412
rect 4846 4398 4850 4402
rect 4702 4388 4706 4392
rect 4766 4388 4770 4392
rect 4798 4388 4802 4392
rect 4782 4368 4786 4372
rect 4766 4348 4770 4352
rect 4694 4338 4698 4342
rect 4710 4338 4714 4342
rect 4726 4338 4730 4342
rect 4750 4338 4754 4342
rect 4774 4328 4778 4332
rect 4742 4278 4746 4282
rect 4758 4278 4762 4282
rect 4702 4258 4706 4262
rect 4710 4158 4714 4162
rect 4702 4148 4706 4152
rect 4710 4148 4714 4152
rect 4678 4138 4682 4142
rect 4694 4138 4698 4142
rect 4710 4128 4714 4132
rect 4854 4358 4858 4362
rect 4878 4358 4882 4362
rect 4894 4358 4898 4362
rect 4806 4348 4810 4352
rect 4830 4348 4834 4352
rect 4806 4338 4810 4342
rect 4790 4318 4794 4322
rect 4886 4348 4890 4352
rect 4870 4308 4874 4312
rect 4870 4288 4874 4292
rect 5086 4958 5090 4962
rect 5078 4938 5082 4942
rect 5046 4898 5050 4902
rect 5046 4848 5050 4852
rect 5062 4868 5066 4872
rect 5078 4868 5082 4872
rect 5086 4858 5090 4862
rect 5094 4848 5098 4852
rect 5054 4838 5058 4842
rect 5078 4838 5082 4842
rect 5054 4798 5058 4802
rect 5046 4768 5050 4772
rect 5046 4748 5050 4752
rect 5070 4738 5074 4742
rect 5046 4718 5050 4722
rect 5022 4698 5026 4702
rect 5038 4698 5042 4702
rect 5022 4678 5026 4682
rect 5046 4678 5050 4682
rect 5062 4658 5066 4662
rect 5142 5018 5146 5022
rect 5150 4928 5154 4932
rect 5174 4918 5178 4922
rect 5166 4888 5170 4892
rect 5166 4878 5170 4882
rect 5134 4778 5138 4782
rect 5102 4768 5106 4772
rect 5086 4698 5090 4702
rect 5134 4738 5138 4742
rect 5118 4728 5122 4732
rect 5086 4668 5090 4672
rect 5150 4808 5154 4812
rect 5142 4708 5146 4712
rect 5158 4748 5162 4752
rect 5166 4738 5170 4742
rect 5246 5058 5250 5062
rect 5302 5048 5306 5052
rect 5230 4908 5234 4912
rect 5302 4948 5306 4952
rect 5246 4878 5250 4882
rect 5254 4878 5258 4882
rect 5246 4868 5250 4872
rect 5238 4858 5242 4862
rect 5278 4858 5282 4862
rect 5262 4848 5266 4852
rect 5222 4838 5226 4842
rect 5302 4848 5306 4852
rect 5286 4818 5290 4822
rect 5238 4788 5242 4792
rect 5262 4788 5266 4792
rect 5190 4768 5194 4772
rect 5238 4748 5242 4752
rect 5222 4728 5226 4732
rect 5182 4718 5186 4722
rect 5166 4688 5170 4692
rect 5198 4668 5202 4672
rect 5246 4668 5250 4672
rect 5038 4648 5042 4652
rect 5078 4648 5082 4652
rect 5054 4638 5058 4642
rect 5054 4618 5058 4622
rect 5038 4538 5042 4542
rect 5014 4528 5018 4532
rect 5022 4528 5026 4532
rect 5006 4508 5010 4512
rect 4998 4498 5002 4502
rect 4982 4478 4986 4482
rect 4998 4478 5002 4482
rect 5030 4518 5034 4522
rect 5014 4468 5018 4472
rect 4958 4438 4962 4442
rect 4982 4438 4986 4442
rect 5014 4448 5018 4452
rect 5022 4448 5026 4452
rect 5014 4418 5018 4422
rect 4918 4348 4922 4352
rect 4910 4338 4914 4342
rect 5006 4338 5010 4342
rect 4938 4303 4942 4307
rect 4945 4303 4949 4307
rect 4958 4288 4962 4292
rect 4982 4278 4986 4282
rect 4758 4258 4762 4262
rect 4790 4258 4794 4262
rect 4814 4258 4818 4262
rect 4846 4258 4850 4262
rect 4774 4228 4778 4232
rect 4766 4198 4770 4202
rect 4742 4178 4746 4182
rect 4734 4168 4738 4172
rect 4798 4248 4802 4252
rect 4782 4188 4786 4192
rect 4758 4148 4762 4152
rect 4790 4148 4794 4152
rect 4926 4248 4930 4252
rect 4846 4188 4850 4192
rect 4734 4138 4738 4142
rect 4742 4128 4746 4132
rect 4710 4118 4714 4122
rect 4726 4118 4730 4122
rect 4654 4098 4658 4102
rect 4726 4098 4730 4102
rect 4710 4078 4714 4082
rect 4670 4058 4674 4062
rect 4654 3988 4658 3992
rect 4726 3958 4730 3962
rect 4614 3948 4618 3952
rect 4646 3928 4650 3932
rect 4622 3908 4626 3912
rect 4550 3868 4554 3872
rect 4574 3868 4578 3872
rect 4606 3868 4610 3872
rect 4454 3858 4458 3862
rect 4486 3858 4490 3862
rect 4526 3848 4530 3852
rect 4494 3828 4498 3832
rect 4510 3788 4514 3792
rect 4542 3768 4546 3772
rect 4406 3748 4410 3752
rect 4462 3748 4466 3752
rect 4494 3748 4498 3752
rect 4542 3738 4546 3742
rect 4390 3728 4394 3732
rect 4414 3718 4418 3722
rect 4502 3718 4506 3722
rect 4366 3688 4370 3692
rect 4414 3698 4418 3702
rect 4406 3688 4410 3692
rect 4630 3768 4634 3772
rect 4614 3758 4618 3762
rect 4622 3758 4626 3762
rect 4622 3748 4626 3752
rect 4574 3738 4578 3742
rect 4446 3688 4450 3692
rect 4534 3688 4538 3692
rect 4542 3678 4546 3682
rect 4358 3668 4362 3672
rect 4246 3658 4250 3662
rect 4310 3658 4314 3662
rect 4246 3648 4250 3652
rect 4254 3638 4258 3642
rect 4342 3658 4346 3662
rect 4350 3658 4354 3662
rect 4390 3658 4394 3662
rect 4278 3648 4282 3652
rect 4270 3628 4274 3632
rect 4310 3588 4314 3592
rect 4222 3558 4226 3562
rect 4174 3548 4178 3552
rect 4190 3548 4194 3552
rect 4222 3548 4226 3552
rect 4158 3528 4162 3532
rect 4142 3498 4146 3502
rect 4174 3478 4178 3482
rect 4214 3528 4218 3532
rect 4214 3508 4218 3512
rect 4206 3488 4210 3492
rect 4238 3488 4242 3492
rect 4142 3458 4146 3462
rect 4190 3428 4194 3432
rect 4126 3348 4130 3352
rect 4102 3318 4106 3322
rect 4094 3298 4098 3302
rect 4078 3278 4082 3282
rect 4038 3268 4042 3272
rect 4126 3268 4130 3272
rect 4046 3258 4050 3262
rect 4078 3258 4082 3262
rect 4054 3238 4058 3242
rect 4030 3198 4034 3202
rect 3998 3168 4002 3172
rect 3982 3068 3986 3072
rect 4046 3158 4050 3162
rect 4030 3148 4034 3152
rect 4014 3128 4018 3132
rect 4030 3088 4034 3092
rect 4046 3088 4050 3092
rect 4038 3068 4042 3072
rect 3958 3058 3962 3062
rect 4030 3058 4034 3062
rect 3998 3038 4002 3042
rect 4110 3188 4114 3192
rect 4102 3158 4106 3162
rect 4086 3148 4090 3152
rect 4134 3228 4138 3232
rect 4166 3338 4170 3342
rect 4182 3288 4186 3292
rect 4182 3228 4186 3232
rect 4150 3198 4154 3202
rect 4142 3188 4146 3192
rect 4142 3168 4146 3172
rect 4166 3188 4170 3192
rect 4134 3148 4138 3152
rect 4158 3148 4162 3152
rect 4118 3138 4122 3142
rect 4070 3128 4074 3132
rect 4062 3118 4066 3122
rect 4134 3088 4138 3092
rect 4294 3508 4298 3512
rect 4326 3558 4330 3562
rect 4350 3548 4354 3552
rect 4398 3568 4402 3572
rect 4446 3648 4450 3652
rect 4426 3603 4430 3607
rect 4433 3603 4437 3607
rect 4590 3688 4594 3692
rect 4750 4098 4754 4102
rect 4822 4108 4826 4112
rect 4806 4078 4810 4082
rect 4894 4158 4898 4162
rect 4870 4148 4874 4152
rect 4854 4138 4858 4142
rect 4878 4138 4882 4142
rect 4894 4138 4898 4142
rect 4910 4138 4914 4142
rect 4838 4128 4842 4132
rect 4902 4128 4906 4132
rect 4938 4103 4942 4107
rect 4945 4103 4949 4107
rect 4966 4088 4970 4092
rect 4918 4078 4922 4082
rect 4886 4058 4890 4062
rect 4854 4038 4858 4042
rect 4830 4028 4834 4032
rect 4958 4028 4962 4032
rect 4742 4018 4746 4022
rect 4846 4008 4850 4012
rect 4822 3988 4826 3992
rect 4750 3968 4754 3972
rect 4790 3968 4794 3972
rect 4742 3948 4746 3952
rect 4734 3938 4738 3942
rect 4726 3918 4730 3922
rect 4678 3828 4682 3832
rect 4734 3828 4738 3832
rect 4654 3768 4658 3772
rect 4702 3768 4706 3772
rect 4662 3738 4666 3742
rect 4646 3728 4650 3732
rect 4678 3728 4682 3732
rect 4726 3758 4730 3762
rect 4662 3688 4666 3692
rect 4678 3688 4682 3692
rect 4710 3688 4714 3692
rect 4566 3658 4570 3662
rect 4630 3658 4634 3662
rect 4478 3648 4482 3652
rect 4606 3648 4610 3652
rect 4358 3538 4362 3542
rect 4366 3538 4370 3542
rect 4382 3538 4386 3542
rect 4334 3528 4338 3532
rect 4390 3528 4394 3532
rect 4342 3518 4346 3522
rect 4398 3518 4402 3522
rect 4318 3508 4322 3512
rect 4334 3488 4338 3492
rect 4414 3538 4418 3542
rect 4406 3488 4410 3492
rect 4662 3648 4666 3652
rect 4646 3628 4650 3632
rect 4462 3608 4466 3612
rect 4630 3598 4634 3602
rect 4614 3588 4618 3592
rect 4558 3578 4562 3582
rect 4566 3568 4570 3572
rect 4494 3558 4498 3562
rect 4510 3558 4514 3562
rect 4526 3558 4530 3562
rect 4478 3548 4482 3552
rect 4534 3548 4538 3552
rect 4270 3478 4274 3482
rect 4366 3478 4370 3482
rect 4454 3478 4458 3482
rect 4246 3468 4250 3472
rect 4230 3448 4234 3452
rect 4214 3438 4218 3442
rect 4214 3428 4218 3432
rect 4198 3308 4202 3312
rect 4198 3288 4202 3292
rect 4278 3468 4282 3472
rect 4238 3348 4242 3352
rect 4254 3348 4258 3352
rect 4246 3338 4250 3342
rect 4214 3278 4218 3282
rect 4230 3268 4234 3272
rect 4326 3418 4330 3422
rect 4302 3388 4306 3392
rect 4310 3358 4314 3362
rect 4302 3338 4306 3342
rect 4278 3328 4282 3332
rect 4270 3308 4274 3312
rect 4294 3308 4298 3312
rect 4286 3278 4290 3282
rect 4426 3403 4430 3407
rect 4433 3403 4437 3407
rect 4406 3378 4410 3382
rect 4390 3368 4394 3372
rect 4366 3348 4370 3352
rect 4358 3328 4362 3332
rect 4398 3328 4402 3332
rect 4350 3318 4354 3322
rect 4334 3288 4338 3292
rect 4206 3258 4210 3262
rect 4262 3248 4266 3252
rect 4270 3238 4274 3242
rect 4254 3208 4258 3212
rect 4190 3158 4194 3162
rect 4182 3148 4186 3152
rect 4182 3128 4186 3132
rect 4166 3068 4170 3072
rect 4238 3098 4242 3102
rect 4198 3058 4202 3062
rect 4230 3058 4234 3062
rect 4102 3048 4106 3052
rect 4174 3048 4178 3052
rect 4086 3038 4090 3042
rect 4006 3028 4010 3032
rect 4054 3028 4058 3032
rect 4062 3018 4066 3022
rect 3974 2958 3978 2962
rect 3942 2948 3946 2952
rect 3934 2928 3938 2932
rect 3922 2903 3926 2907
rect 3929 2903 3933 2907
rect 3910 2868 3914 2872
rect 3910 2778 3914 2782
rect 3958 2938 3962 2942
rect 3982 2948 3986 2952
rect 3958 2928 3962 2932
rect 3982 2928 3986 2932
rect 4006 2968 4010 2972
rect 4022 2958 4026 2962
rect 4054 2958 4058 2962
rect 4134 3028 4138 3032
rect 4158 2958 4162 2962
rect 4022 2938 4026 2942
rect 4078 2938 4082 2942
rect 3966 2898 3970 2902
rect 3998 2898 4002 2902
rect 3958 2758 3962 2762
rect 3894 2748 3898 2752
rect 3950 2748 3954 2752
rect 3830 2658 3834 2662
rect 3750 2648 3754 2652
rect 3750 2608 3754 2612
rect 3750 2568 3754 2572
rect 3702 2538 3706 2542
rect 3734 2538 3738 2542
rect 3750 2528 3754 2532
rect 3790 2568 3794 2572
rect 3782 2548 3786 2552
rect 3774 2528 3778 2532
rect 3766 2508 3770 2512
rect 3718 2488 3722 2492
rect 3742 2488 3746 2492
rect 3710 2478 3714 2482
rect 3686 2468 3690 2472
rect 3702 2468 3706 2472
rect 3750 2448 3754 2452
rect 3782 2448 3786 2452
rect 3734 2438 3738 2442
rect 3662 2428 3666 2432
rect 3694 2428 3698 2432
rect 3742 2428 3746 2432
rect 3726 2418 3730 2422
rect 3662 2398 3666 2402
rect 3662 2338 3666 2342
rect 3638 2308 3642 2312
rect 3614 2288 3618 2292
rect 3622 2268 3626 2272
rect 3614 2248 3618 2252
rect 3670 2298 3674 2302
rect 3638 2238 3642 2242
rect 3646 2218 3650 2222
rect 3654 2218 3658 2222
rect 3630 2168 3634 2172
rect 3614 2108 3618 2112
rect 3614 2098 3618 2102
rect 3662 2198 3666 2202
rect 3686 2408 3690 2412
rect 3694 2388 3698 2392
rect 3742 2398 3746 2402
rect 3742 2388 3746 2392
rect 3734 2378 3738 2382
rect 3758 2378 3762 2382
rect 3766 2378 3770 2382
rect 3686 2348 3690 2352
rect 3694 2348 3698 2352
rect 3750 2348 3754 2352
rect 3750 2318 3754 2322
rect 4030 2928 4034 2932
rect 4110 2928 4114 2932
rect 4022 2888 4026 2892
rect 3990 2878 3994 2882
rect 3998 2868 4002 2872
rect 3982 2858 3986 2862
rect 4014 2858 4018 2862
rect 4038 2858 4042 2862
rect 4054 2898 4058 2902
rect 4126 2898 4130 2902
rect 4118 2888 4122 2892
rect 4094 2878 4098 2882
rect 4030 2848 4034 2852
rect 4046 2848 4050 2852
rect 3998 2838 4002 2842
rect 3990 2798 3994 2802
rect 3878 2728 3882 2732
rect 3942 2728 3946 2732
rect 3902 2718 3906 2722
rect 3922 2703 3926 2707
rect 3929 2703 3933 2707
rect 3950 2688 3954 2692
rect 3894 2678 3898 2682
rect 3950 2678 3954 2682
rect 3886 2668 3890 2672
rect 3862 2658 3866 2662
rect 3870 2658 3874 2662
rect 3854 2648 3858 2652
rect 3862 2588 3866 2592
rect 3846 2558 3850 2562
rect 3878 2638 3882 2642
rect 3814 2548 3818 2552
rect 3806 2538 3810 2542
rect 3870 2538 3874 2542
rect 3878 2538 3882 2542
rect 3854 2528 3858 2532
rect 3870 2528 3874 2532
rect 3822 2518 3826 2522
rect 3814 2508 3818 2512
rect 3790 2378 3794 2382
rect 3806 2378 3810 2382
rect 3790 2368 3794 2372
rect 3814 2358 3818 2362
rect 3814 2328 3818 2332
rect 3774 2308 3778 2312
rect 3814 2298 3818 2302
rect 3734 2288 3738 2292
rect 3774 2288 3778 2292
rect 3718 2268 3722 2272
rect 3750 2278 3754 2282
rect 3782 2278 3786 2282
rect 3782 2258 3786 2262
rect 3710 2238 3714 2242
rect 3718 2198 3722 2202
rect 3766 2188 3770 2192
rect 3774 2178 3778 2182
rect 3702 2138 3706 2142
rect 3710 2118 3714 2122
rect 3734 2108 3738 2112
rect 3830 2508 3834 2512
rect 3830 2468 3834 2472
rect 3838 2358 3842 2362
rect 3830 2318 3834 2322
rect 3870 2498 3874 2502
rect 3862 2428 3866 2432
rect 3934 2668 3938 2672
rect 3902 2508 3906 2512
rect 3894 2478 3898 2482
rect 3894 2458 3898 2462
rect 3886 2438 3890 2442
rect 3862 2368 3866 2372
rect 3878 2368 3882 2372
rect 3854 2298 3858 2302
rect 3878 2358 3882 2362
rect 3870 2348 3874 2352
rect 3974 2728 3978 2732
rect 3966 2678 3970 2682
rect 3958 2668 3962 2672
rect 3974 2668 3978 2672
rect 3966 2568 3970 2572
rect 3974 2548 3978 2552
rect 3958 2538 3962 2542
rect 3926 2528 3930 2532
rect 3974 2528 3978 2532
rect 3922 2503 3926 2507
rect 3929 2503 3933 2507
rect 3934 2468 3938 2472
rect 3918 2448 3922 2452
rect 3894 2398 3898 2402
rect 3910 2398 3914 2402
rect 3918 2378 3922 2382
rect 3966 2368 3970 2372
rect 3958 2358 3962 2362
rect 3958 2348 3962 2352
rect 3886 2298 3890 2302
rect 3862 2288 3866 2292
rect 3878 2268 3882 2272
rect 3838 2248 3842 2252
rect 3894 2268 3898 2272
rect 3846 2238 3850 2242
rect 3862 2198 3866 2202
rect 3822 2178 3826 2182
rect 3950 2338 3954 2342
rect 3926 2328 3930 2332
rect 3922 2303 3926 2307
rect 3929 2303 3933 2307
rect 3910 2298 3914 2302
rect 3918 2268 3922 2272
rect 3870 2188 3874 2192
rect 3910 2188 3914 2192
rect 3838 2158 3842 2162
rect 3790 2138 3794 2142
rect 3798 2108 3802 2112
rect 3678 2088 3682 2092
rect 3726 2088 3730 2092
rect 3622 2078 3626 2082
rect 3678 2078 3682 2082
rect 3606 2058 3610 2062
rect 3646 2058 3650 2062
rect 3614 2038 3618 2042
rect 3582 1968 3586 1972
rect 3542 1938 3546 1942
rect 3582 1938 3586 1942
rect 3550 1918 3554 1922
rect 3526 1898 3530 1902
rect 3518 1868 3522 1872
rect 3526 1868 3530 1872
rect 3534 1858 3538 1862
rect 3486 1848 3490 1852
rect 3502 1848 3506 1852
rect 3438 1838 3442 1842
rect 3390 1828 3394 1832
rect 3502 1838 3506 1842
rect 3454 1818 3458 1822
rect 3402 1803 3406 1807
rect 3409 1803 3413 1807
rect 3526 1828 3530 1832
rect 3518 1778 3522 1782
rect 3494 1758 3498 1762
rect 3382 1748 3386 1752
rect 3438 1748 3442 1752
rect 3510 1748 3514 1752
rect 3390 1738 3394 1742
rect 3294 1728 3298 1732
rect 3342 1728 3346 1732
rect 3358 1728 3362 1732
rect 3302 1688 3306 1692
rect 3414 1708 3418 1712
rect 3358 1688 3362 1692
rect 3334 1668 3338 1672
rect 3342 1668 3346 1672
rect 3334 1658 3338 1662
rect 3462 1688 3466 1692
rect 3558 1898 3562 1902
rect 3606 1938 3610 1942
rect 3638 2048 3642 2052
rect 3654 2038 3658 2042
rect 3630 1978 3634 1982
rect 3638 1948 3642 1952
rect 3630 1928 3634 1932
rect 3614 1888 3618 1892
rect 3598 1878 3602 1882
rect 3582 1868 3586 1872
rect 3622 1868 3626 1872
rect 3598 1858 3602 1862
rect 3542 1748 3546 1752
rect 3566 1748 3570 1752
rect 3534 1738 3538 1742
rect 3518 1728 3522 1732
rect 3542 1728 3546 1732
rect 3470 1678 3474 1682
rect 3486 1678 3490 1682
rect 3446 1668 3450 1672
rect 3390 1658 3394 1662
rect 3398 1658 3402 1662
rect 3422 1658 3426 1662
rect 3478 1658 3482 1662
rect 3350 1648 3354 1652
rect 3374 1648 3378 1652
rect 3366 1608 3370 1612
rect 3254 1558 3258 1562
rect 3278 1558 3282 1562
rect 3238 1548 3242 1552
rect 3342 1548 3346 1552
rect 3150 1538 3154 1542
rect 3190 1508 3194 1512
rect 3150 1498 3154 1502
rect 3070 1458 3074 1462
rect 3118 1458 3122 1462
rect 3102 1448 3106 1452
rect 3078 1428 3082 1432
rect 3070 1378 3074 1382
rect 2958 1368 2962 1372
rect 2974 1368 2978 1372
rect 3054 1368 3058 1372
rect 3006 1348 3010 1352
rect 3054 1348 3058 1352
rect 3166 1448 3170 1452
rect 3134 1438 3138 1442
rect 3126 1398 3130 1402
rect 3118 1388 3122 1392
rect 3174 1388 3178 1392
rect 3158 1368 3162 1372
rect 3174 1368 3178 1372
rect 3150 1358 3154 1362
rect 3134 1348 3138 1352
rect 2966 1338 2970 1342
rect 3038 1338 3042 1342
rect 3062 1338 3066 1342
rect 2990 1328 2994 1332
rect 3070 1308 3074 1312
rect 3078 1298 3082 1302
rect 2966 1288 2970 1292
rect 2958 1278 2962 1282
rect 2942 1258 2946 1262
rect 2982 1258 2986 1262
rect 3142 1338 3146 1342
rect 3102 1298 3106 1302
rect 3150 1318 3154 1322
rect 3118 1288 3122 1292
rect 3150 1268 3154 1272
rect 3206 1498 3210 1502
rect 3254 1538 3258 1542
rect 3286 1538 3290 1542
rect 3302 1538 3306 1542
rect 3350 1538 3354 1542
rect 3262 1528 3266 1532
rect 3342 1528 3346 1532
rect 3230 1518 3234 1522
rect 3254 1498 3258 1502
rect 3222 1408 3226 1412
rect 3206 1338 3210 1342
rect 3182 1288 3186 1292
rect 3230 1318 3234 1322
rect 3238 1288 3242 1292
rect 3270 1508 3274 1512
rect 3294 1498 3298 1502
rect 3326 1508 3330 1512
rect 3310 1488 3314 1492
rect 3278 1478 3282 1482
rect 3402 1603 3406 1607
rect 3409 1603 3413 1607
rect 3502 1598 3506 1602
rect 3382 1578 3386 1582
rect 3374 1568 3378 1572
rect 3478 1558 3482 1562
rect 3430 1528 3434 1532
rect 3390 1518 3394 1522
rect 3382 1498 3386 1502
rect 3350 1458 3354 1462
rect 3310 1438 3314 1442
rect 3366 1438 3370 1442
rect 3270 1358 3274 1362
rect 3294 1358 3298 1362
rect 3270 1338 3274 1342
rect 3302 1328 3306 1332
rect 3214 1268 3218 1272
rect 3222 1268 3226 1272
rect 3246 1268 3250 1272
rect 3006 1258 3010 1262
rect 3078 1258 3082 1262
rect 3086 1258 3090 1262
rect 3094 1258 3098 1262
rect 3158 1258 3162 1262
rect 2926 1248 2930 1252
rect 2942 1248 2946 1252
rect 2950 1238 2954 1242
rect 2878 1218 2882 1222
rect 2870 1188 2874 1192
rect 2926 1198 2930 1202
rect 2862 1158 2866 1162
rect 2846 1148 2850 1152
rect 2822 1138 2826 1142
rect 2894 1138 2898 1142
rect 2910 1138 2914 1142
rect 2806 1128 2810 1132
rect 2846 1128 2850 1132
rect 2798 1088 2802 1092
rect 2774 1078 2778 1082
rect 2782 1078 2786 1082
rect 2814 1078 2818 1082
rect 2782 1058 2786 1062
rect 2774 1038 2778 1042
rect 2550 1028 2554 1032
rect 2606 1028 2610 1032
rect 2590 968 2594 972
rect 2838 1028 2842 1032
rect 2806 1018 2810 1022
rect 2758 1008 2762 1012
rect 2670 978 2674 982
rect 2718 978 2722 982
rect 2630 968 2634 972
rect 2558 958 2562 962
rect 2606 958 2610 962
rect 2510 878 2514 882
rect 2526 868 2530 872
rect 2694 968 2698 972
rect 2638 958 2642 962
rect 2662 958 2666 962
rect 2654 948 2658 952
rect 2598 938 2602 942
rect 2654 938 2658 942
rect 2606 918 2610 922
rect 2638 918 2642 922
rect 2590 868 2594 872
rect 2550 838 2554 842
rect 2582 808 2586 812
rect 2606 848 2610 852
rect 2614 848 2618 852
rect 2630 848 2634 852
rect 2598 828 2602 832
rect 2598 808 2602 812
rect 2590 768 2594 772
rect 2486 728 2490 732
rect 2486 718 2490 722
rect 2486 678 2490 682
rect 2510 678 2514 682
rect 2654 828 2658 832
rect 2646 808 2650 812
rect 2630 788 2634 792
rect 2614 758 2618 762
rect 2638 768 2642 772
rect 2646 748 2650 752
rect 2630 738 2634 742
rect 2606 718 2610 722
rect 2590 698 2594 702
rect 2574 668 2578 672
rect 2478 658 2482 662
rect 2494 658 2498 662
rect 2502 628 2506 632
rect 2510 598 2514 602
rect 2502 588 2506 592
rect 2486 558 2490 562
rect 2566 547 2570 551
rect 2558 538 2562 542
rect 2510 528 2514 532
rect 2502 508 2506 512
rect 2470 488 2474 492
rect 2574 508 2578 512
rect 2574 478 2578 482
rect 2534 468 2538 472
rect 2518 458 2522 462
rect 2446 448 2450 452
rect 2462 448 2466 452
rect 2470 438 2474 442
rect 2470 428 2474 432
rect 2462 358 2466 362
rect 2446 348 2450 352
rect 2454 338 2458 342
rect 2422 308 2426 312
rect 2438 308 2442 312
rect 2478 298 2482 302
rect 2454 288 2458 292
rect 2422 268 2426 272
rect 2386 203 2390 207
rect 2393 203 2397 207
rect 2398 168 2402 172
rect 2334 148 2338 152
rect 2358 148 2362 152
rect 2486 278 2490 282
rect 2470 268 2474 272
rect 2558 438 2562 442
rect 2566 438 2570 442
rect 2606 678 2610 682
rect 2678 948 2682 952
rect 2742 958 2746 962
rect 2710 948 2714 952
rect 2830 978 2834 982
rect 2782 958 2786 962
rect 2806 958 2810 962
rect 2702 938 2706 942
rect 2750 938 2754 942
rect 2710 918 2714 922
rect 2726 898 2730 902
rect 2702 878 2706 882
rect 2718 858 2722 862
rect 2758 918 2762 922
rect 2782 938 2786 942
rect 2774 878 2778 882
rect 2742 818 2746 822
rect 2862 1118 2866 1122
rect 2870 1118 2874 1122
rect 2854 958 2858 962
rect 2846 928 2850 932
rect 2838 898 2842 902
rect 2854 878 2858 882
rect 2798 868 2802 872
rect 2814 868 2818 872
rect 2814 858 2818 862
rect 2814 828 2818 832
rect 2830 828 2834 832
rect 2822 798 2826 802
rect 2838 758 2842 762
rect 2890 1103 2894 1107
rect 2897 1103 2901 1107
rect 2870 1098 2874 1102
rect 2886 1088 2890 1092
rect 2878 1068 2882 1072
rect 2910 1058 2914 1062
rect 3054 1248 3058 1252
rect 3078 1228 3082 1232
rect 2958 1218 2962 1222
rect 3030 1218 3034 1222
rect 3014 1208 3018 1212
rect 2990 1158 2994 1162
rect 3070 1188 3074 1192
rect 3046 1168 3050 1172
rect 3150 1208 3154 1212
rect 3126 1188 3130 1192
rect 3078 1158 3082 1162
rect 3102 1158 3106 1162
rect 2958 1148 2962 1152
rect 2982 1148 2986 1152
rect 3006 1148 3010 1152
rect 3022 1148 3026 1152
rect 3134 1148 3138 1152
rect 2950 1118 2954 1122
rect 2966 1088 2970 1092
rect 3014 1138 3018 1142
rect 3046 1138 3050 1142
rect 2934 1058 2938 1062
rect 2918 968 2922 972
rect 2910 958 2914 962
rect 2910 948 2914 952
rect 2870 938 2874 942
rect 2902 938 2906 942
rect 2894 928 2898 932
rect 2890 903 2894 907
rect 2897 903 2901 907
rect 2862 868 2866 872
rect 2942 1028 2946 1032
rect 2966 1028 2970 1032
rect 2958 968 2962 972
rect 2926 888 2930 892
rect 2934 888 2938 892
rect 2974 938 2978 942
rect 3022 1118 3026 1122
rect 3038 1068 3042 1072
rect 3022 1058 3026 1062
rect 3006 1028 3010 1032
rect 3022 1028 3026 1032
rect 2990 1018 2994 1022
rect 3086 1118 3090 1122
rect 3094 1108 3098 1112
rect 3070 1088 3074 1092
rect 3054 958 3058 962
rect 3086 1058 3090 1062
rect 3294 1318 3298 1322
rect 3286 1298 3290 1302
rect 3278 1258 3282 1262
rect 3270 1248 3274 1252
rect 3294 1248 3298 1252
rect 3262 1238 3266 1242
rect 3294 1218 3298 1222
rect 3214 1208 3218 1212
rect 3230 1198 3234 1202
rect 3246 1178 3250 1182
rect 3278 1158 3282 1162
rect 3166 1148 3170 1152
rect 3254 1148 3258 1152
rect 3270 1148 3274 1152
rect 3286 1148 3290 1152
rect 3158 1138 3162 1142
rect 3174 1128 3178 1132
rect 3270 1128 3274 1132
rect 3134 1118 3138 1122
rect 3286 1118 3290 1122
rect 3158 1108 3162 1112
rect 3206 1108 3210 1112
rect 3230 1108 3234 1112
rect 3150 1088 3154 1092
rect 3270 1088 3274 1092
rect 3134 1078 3138 1082
rect 3262 1078 3266 1082
rect 3206 1068 3210 1072
rect 3246 1068 3250 1072
rect 3254 1068 3258 1072
rect 3262 1058 3266 1062
rect 3366 1398 3370 1402
rect 3326 1378 3330 1382
rect 3358 1358 3362 1362
rect 3430 1488 3434 1492
rect 3470 1498 3474 1502
rect 3582 1738 3586 1742
rect 3646 1908 3650 1912
rect 3638 1878 3642 1882
rect 3758 2078 3762 2082
rect 3702 2058 3706 2062
rect 3718 2058 3722 2062
rect 3742 2058 3746 2062
rect 3790 2058 3794 2062
rect 3686 2048 3690 2052
rect 3694 2028 3698 2032
rect 3718 1948 3722 1952
rect 3670 1928 3674 1932
rect 3678 1918 3682 1922
rect 3670 1898 3674 1902
rect 3702 1908 3706 1912
rect 3686 1898 3690 1902
rect 3654 1868 3658 1872
rect 3678 1878 3682 1882
rect 3686 1878 3690 1882
rect 3694 1868 3698 1872
rect 3646 1858 3650 1862
rect 3670 1848 3674 1852
rect 3678 1848 3682 1852
rect 3670 1828 3674 1832
rect 3630 1758 3634 1762
rect 3606 1728 3610 1732
rect 3614 1688 3618 1692
rect 3654 1748 3658 1752
rect 3670 1738 3674 1742
rect 3638 1698 3642 1702
rect 3558 1668 3562 1672
rect 3630 1678 3634 1682
rect 3662 1678 3666 1682
rect 3646 1668 3650 1672
rect 3550 1658 3554 1662
rect 3646 1658 3650 1662
rect 3670 1658 3674 1662
rect 3574 1618 3578 1622
rect 3566 1558 3570 1562
rect 3542 1548 3546 1552
rect 3486 1538 3490 1542
rect 3486 1508 3490 1512
rect 3486 1488 3490 1492
rect 3478 1468 3482 1472
rect 3470 1458 3474 1462
rect 3438 1448 3442 1452
rect 3438 1428 3442 1432
rect 3402 1403 3406 1407
rect 3409 1403 3413 1407
rect 3390 1388 3394 1392
rect 3374 1358 3378 1362
rect 3398 1368 3402 1372
rect 3406 1358 3410 1362
rect 3422 1358 3426 1362
rect 3454 1358 3458 1362
rect 3334 1338 3338 1342
rect 3366 1338 3370 1342
rect 3374 1338 3378 1342
rect 3318 1328 3322 1332
rect 3318 1288 3322 1292
rect 3334 1248 3338 1252
rect 3310 1208 3314 1212
rect 3382 1268 3386 1272
rect 3366 1208 3370 1212
rect 3310 1158 3314 1162
rect 3350 1158 3354 1162
rect 3358 1158 3362 1162
rect 3438 1328 3442 1332
rect 3526 1538 3530 1542
rect 3534 1528 3538 1532
rect 3558 1508 3562 1512
rect 3526 1498 3530 1502
rect 3510 1468 3514 1472
rect 3542 1448 3546 1452
rect 3502 1378 3506 1382
rect 3670 1648 3674 1652
rect 3710 1858 3714 1862
rect 3726 1947 3730 1951
rect 3782 1998 3786 2002
rect 3774 1948 3778 1952
rect 3750 1878 3754 1882
rect 3726 1868 3730 1872
rect 3734 1868 3738 1872
rect 3694 1808 3698 1812
rect 3694 1758 3698 1762
rect 3734 1818 3738 1822
rect 3750 1738 3754 1742
rect 3718 1688 3722 1692
rect 3710 1668 3714 1672
rect 3742 1668 3746 1672
rect 3750 1668 3754 1672
rect 3702 1658 3706 1662
rect 3678 1638 3682 1642
rect 3622 1588 3626 1592
rect 3646 1558 3650 1562
rect 3590 1538 3594 1542
rect 3574 1528 3578 1532
rect 3622 1538 3626 1542
rect 3606 1528 3610 1532
rect 3582 1448 3586 1452
rect 3646 1518 3650 1522
rect 3638 1498 3642 1502
rect 3830 2148 3834 2152
rect 3862 2148 3866 2152
rect 3838 2138 3842 2142
rect 3822 2118 3826 2122
rect 3814 2108 3818 2112
rect 3806 2088 3810 2092
rect 3822 2078 3826 2082
rect 3942 2268 3946 2272
rect 4022 2768 4026 2772
rect 4038 2768 4042 2772
rect 4022 2748 4026 2752
rect 4062 2768 4066 2772
rect 4046 2758 4050 2762
rect 4086 2758 4090 2762
rect 4046 2748 4050 2752
rect 4094 2748 4098 2752
rect 4078 2728 4082 2732
rect 4094 2718 4098 2722
rect 4062 2708 4066 2712
rect 3998 2698 4002 2702
rect 4038 2678 4042 2682
rect 4014 2668 4018 2672
rect 3998 2648 4002 2652
rect 4022 2618 4026 2622
rect 4222 3008 4226 3012
rect 4198 2998 4202 3002
rect 4214 2968 4218 2972
rect 4206 2948 4210 2952
rect 4198 2938 4202 2942
rect 4174 2928 4178 2932
rect 4190 2898 4194 2902
rect 4158 2888 4162 2892
rect 4174 2888 4178 2892
rect 4174 2878 4178 2882
rect 4166 2868 4170 2872
rect 4174 2858 4178 2862
rect 4126 2798 4130 2802
rect 4118 2788 4122 2792
rect 4110 2758 4114 2762
rect 4126 2768 4130 2772
rect 4166 2798 4170 2802
rect 4174 2758 4178 2762
rect 4198 2788 4202 2792
rect 4230 2888 4234 2892
rect 4222 2868 4226 2872
rect 4238 2848 4242 2852
rect 4230 2768 4234 2772
rect 4198 2758 4202 2762
rect 4182 2748 4186 2752
rect 4142 2698 4146 2702
rect 4118 2688 4122 2692
rect 4134 2688 4138 2692
rect 4102 2648 4106 2652
rect 4062 2638 4066 2642
rect 4062 2628 4066 2632
rect 4102 2618 4106 2622
rect 4110 2588 4114 2592
rect 4070 2548 4074 2552
rect 4062 2498 4066 2502
rect 4054 2468 4058 2472
rect 4006 2458 4010 2462
rect 4030 2458 4034 2462
rect 3982 2448 3986 2452
rect 4006 2448 4010 2452
rect 4094 2508 4098 2512
rect 4150 2678 4154 2682
rect 4198 2678 4202 2682
rect 4134 2668 4138 2672
rect 4214 2668 4218 2672
rect 4302 3228 4306 3232
rect 4286 3158 4290 3162
rect 4286 3148 4290 3152
rect 4262 3128 4266 3132
rect 4270 3098 4274 3102
rect 4262 3078 4266 3082
rect 4318 3248 4322 3252
rect 4342 3268 4346 3272
rect 4358 3288 4362 3292
rect 4358 3268 4362 3272
rect 4478 3528 4482 3532
rect 4470 3498 4474 3502
rect 4494 3518 4498 3522
rect 4510 3508 4514 3512
rect 4518 3498 4522 3502
rect 4494 3458 4498 3462
rect 4470 3398 4474 3402
rect 4486 3368 4490 3372
rect 4550 3548 4554 3552
rect 4582 3558 4586 3562
rect 4598 3558 4602 3562
rect 4686 3638 4690 3642
rect 4646 3578 4650 3582
rect 4686 3558 4690 3562
rect 4606 3548 4610 3552
rect 4654 3548 4658 3552
rect 4614 3538 4618 3542
rect 4638 3538 4642 3542
rect 4574 3518 4578 3522
rect 4590 3498 4594 3502
rect 4582 3478 4586 3482
rect 4606 3458 4610 3462
rect 4598 3438 4602 3442
rect 4502 3378 4506 3382
rect 4518 3378 4522 3382
rect 4542 3378 4546 3382
rect 4566 3378 4570 3382
rect 4494 3358 4498 3362
rect 4614 3368 4618 3372
rect 4566 3348 4570 3352
rect 4502 3338 4506 3342
rect 4550 3338 4554 3342
rect 4590 3338 4594 3342
rect 4486 3308 4490 3312
rect 4478 3298 4482 3302
rect 4478 3288 4482 3292
rect 4462 3268 4466 3272
rect 4486 3268 4490 3272
rect 4414 3258 4418 3262
rect 4406 3248 4410 3252
rect 4398 3228 4402 3232
rect 4426 3203 4430 3207
rect 4433 3203 4437 3207
rect 4358 3198 4362 3202
rect 4374 3188 4378 3192
rect 4382 3188 4386 3192
rect 4350 3168 4354 3172
rect 4358 3168 4362 3172
rect 4334 3158 4338 3162
rect 4342 3158 4346 3162
rect 4438 3158 4442 3162
rect 4422 3148 4426 3152
rect 4430 3148 4434 3152
rect 4478 3258 4482 3262
rect 4518 3288 4522 3292
rect 4526 3288 4530 3292
rect 4542 3278 4546 3282
rect 4510 3258 4514 3262
rect 4470 3228 4474 3232
rect 4470 3218 4474 3222
rect 4462 3208 4466 3212
rect 4494 3198 4498 3202
rect 4582 3328 4586 3332
rect 4582 3278 4586 3282
rect 4534 3258 4538 3262
rect 4574 3258 4578 3262
rect 4542 3248 4546 3252
rect 4566 3248 4570 3252
rect 4590 3268 4594 3272
rect 4646 3498 4650 3502
rect 4630 3438 4634 3442
rect 4638 3348 4642 3352
rect 4806 3958 4810 3962
rect 4822 3958 4826 3962
rect 4806 3948 4810 3952
rect 4790 3918 4794 3922
rect 4870 3978 4874 3982
rect 4854 3958 4858 3962
rect 4910 3958 4914 3962
rect 5078 4548 5082 4552
rect 5038 4378 5042 4382
rect 5046 4368 5050 4372
rect 5030 4358 5034 4362
rect 5030 4348 5034 4352
rect 5046 4328 5050 4332
rect 5078 4488 5082 4492
rect 5062 4478 5066 4482
rect 5062 4368 5066 4372
rect 5062 4358 5066 4362
rect 5054 4278 5058 4282
rect 5070 4318 5074 4322
rect 4990 4268 4994 4272
rect 5006 4268 5010 4272
rect 5022 4268 5026 4272
rect 5062 4268 5066 4272
rect 5014 4258 5018 4262
rect 5054 4258 5058 4262
rect 5022 4228 5026 4232
rect 5046 4238 5050 4242
rect 5030 4208 5034 4212
rect 4990 4148 4994 4152
rect 5070 4168 5074 4172
rect 5078 4148 5082 4152
rect 5046 4118 5050 4122
rect 5046 4078 5050 4082
rect 5006 4068 5010 4072
rect 5046 4058 5050 4062
rect 5014 4048 5018 4052
rect 5054 4038 5058 4042
rect 5078 4028 5082 4032
rect 5102 4658 5106 4662
rect 5134 4658 5138 4662
rect 5094 4598 5098 4602
rect 5094 4528 5098 4532
rect 5142 4648 5146 4652
rect 5118 4638 5122 4642
rect 5142 4578 5146 4582
rect 5118 4568 5122 4572
rect 5190 4588 5194 4592
rect 5190 4568 5194 4572
rect 5150 4558 5154 4562
rect 5158 4558 5162 4562
rect 5190 4558 5194 4562
rect 5206 4558 5210 4562
rect 5118 4538 5122 4542
rect 5134 4548 5138 4552
rect 5142 4538 5146 4542
rect 5166 4538 5170 4542
rect 5182 4538 5186 4542
rect 5166 4528 5170 4532
rect 5190 4528 5194 4532
rect 5134 4518 5138 4522
rect 5126 4508 5130 4512
rect 5166 4508 5170 4512
rect 5110 4488 5114 4492
rect 5126 4488 5130 4492
rect 5102 4478 5106 4482
rect 5214 4528 5218 4532
rect 5254 4518 5258 4522
rect 5206 4488 5210 4492
rect 5150 4478 5154 4482
rect 5198 4478 5202 4482
rect 5118 4468 5122 4472
rect 5118 4458 5122 4462
rect 5102 4448 5106 4452
rect 5158 4468 5162 4472
rect 5182 4468 5186 4472
rect 5254 4468 5258 4472
rect 5166 4458 5170 4462
rect 5190 4458 5194 4462
rect 5230 4448 5234 4452
rect 5110 4338 5114 4342
rect 5134 4418 5138 4422
rect 5206 4418 5210 4422
rect 5142 4358 5146 4362
rect 5174 4348 5178 4352
rect 5246 4348 5250 4352
rect 5198 4328 5202 4332
rect 5174 4308 5178 4312
rect 5174 4298 5178 4302
rect 5150 4288 5154 4292
rect 5142 4278 5146 4282
rect 5166 4268 5170 4272
rect 5110 4258 5114 4262
rect 5126 4258 5130 4262
rect 5110 4218 5114 4222
rect 5118 4218 5122 4222
rect 5110 4188 5114 4192
rect 5110 4178 5114 4182
rect 5110 4128 5114 4132
rect 4998 3968 5002 3972
rect 4894 3948 4898 3952
rect 4910 3948 4914 3952
rect 4950 3948 4954 3952
rect 4846 3928 4850 3932
rect 4918 3928 4922 3932
rect 4958 3928 4962 3932
rect 4894 3908 4898 3912
rect 4894 3878 4898 3882
rect 4918 3878 4922 3882
rect 4938 3903 4942 3907
rect 4945 3903 4949 3907
rect 4838 3868 4842 3872
rect 4862 3868 4866 3872
rect 4750 3858 4754 3862
rect 4750 3828 4754 3832
rect 4742 3768 4746 3772
rect 4790 3858 4794 3862
rect 4846 3858 4850 3862
rect 4894 3858 4898 3862
rect 4870 3848 4874 3852
rect 4886 3848 4890 3852
rect 4822 3808 4826 3812
rect 4790 3788 4794 3792
rect 4822 3788 4826 3792
rect 4798 3768 4802 3772
rect 4838 3758 4842 3762
rect 4766 3748 4770 3752
rect 4750 3738 4754 3742
rect 4766 3668 4770 3672
rect 4734 3548 4738 3552
rect 4734 3538 4738 3542
rect 4702 3508 4706 3512
rect 4678 3488 4682 3492
rect 4694 3488 4698 3492
rect 4710 3488 4714 3492
rect 4654 3468 4658 3472
rect 4718 3468 4722 3472
rect 4694 3458 4698 3462
rect 4726 3458 4730 3462
rect 4662 3428 4666 3432
rect 4686 3438 4690 3442
rect 4654 3368 4658 3372
rect 4662 3358 4666 3362
rect 4742 3498 4746 3502
rect 4734 3378 4738 3382
rect 4718 3358 4722 3362
rect 4774 3648 4778 3652
rect 4862 3818 4866 3822
rect 4910 3808 4914 3812
rect 4854 3788 4858 3792
rect 4910 3768 4914 3772
rect 4958 3798 4962 3802
rect 4942 3768 4946 3772
rect 4926 3758 4930 3762
rect 4902 3748 4906 3752
rect 4918 3748 4922 3752
rect 4838 3738 4842 3742
rect 4862 3738 4866 3742
rect 4846 3728 4850 3732
rect 4862 3728 4866 3732
rect 4918 3728 4922 3732
rect 4790 3718 4794 3722
rect 4838 3688 4842 3692
rect 4830 3658 4834 3662
rect 4854 3658 4858 3662
rect 4878 3658 4882 3662
rect 4938 3703 4942 3707
rect 4945 3703 4949 3707
rect 4958 3668 4962 3672
rect 4814 3638 4818 3642
rect 4782 3608 4786 3612
rect 4790 3548 4794 3552
rect 4814 3538 4818 3542
rect 4766 3478 4770 3482
rect 4846 3508 4850 3512
rect 4814 3468 4818 3472
rect 4846 3468 4850 3472
rect 4766 3458 4770 3462
rect 4798 3458 4802 3462
rect 4766 3448 4770 3452
rect 4758 3368 4762 3372
rect 4742 3348 4746 3352
rect 4758 3348 4762 3352
rect 4782 3348 4786 3352
rect 4798 3348 4802 3352
rect 4630 3318 4634 3322
rect 4646 3308 4650 3312
rect 4638 3268 4642 3272
rect 4598 3258 4602 3262
rect 4614 3258 4618 3262
rect 4598 3248 4602 3252
rect 4598 3238 4602 3242
rect 4526 3198 4530 3202
rect 4582 3198 4586 3202
rect 4598 3198 4602 3202
rect 4518 3178 4522 3182
rect 4494 3168 4498 3172
rect 4518 3148 4522 3152
rect 4550 3178 4554 3182
rect 4582 3178 4586 3182
rect 4542 3168 4546 3172
rect 4558 3168 4562 3172
rect 4534 3158 4538 3162
rect 4582 3148 4586 3152
rect 4590 3148 4594 3152
rect 4350 3138 4354 3142
rect 4446 3138 4450 3142
rect 4590 3138 4594 3142
rect 4334 3118 4338 3122
rect 4310 3098 4314 3102
rect 4310 3068 4314 3072
rect 4302 3058 4306 3062
rect 4262 3048 4266 3052
rect 4294 3048 4298 3052
rect 4310 3028 4314 3032
rect 4326 3028 4330 3032
rect 4318 2988 4322 2992
rect 4278 2928 4282 2932
rect 4318 2918 4322 2922
rect 4302 2908 4306 2912
rect 4318 2898 4322 2902
rect 4294 2878 4298 2882
rect 4366 3128 4370 3132
rect 4382 3128 4386 3132
rect 4398 3128 4402 3132
rect 4406 3128 4410 3132
rect 4470 3128 4474 3132
rect 4518 3128 4522 3132
rect 4566 3128 4570 3132
rect 4366 3118 4370 3122
rect 4422 3118 4426 3122
rect 4350 3038 4354 3042
rect 4334 2958 4338 2962
rect 4358 2958 4362 2962
rect 4478 3108 4482 3112
rect 4518 3108 4522 3112
rect 4502 3098 4506 3102
rect 4438 3088 4442 3092
rect 4494 3088 4498 3092
rect 4478 3058 4482 3062
rect 4526 3078 4530 3082
rect 4414 3048 4418 3052
rect 4462 3048 4466 3052
rect 4422 3028 4426 3032
rect 4382 3018 4386 3022
rect 4374 2968 4378 2972
rect 4334 2888 4338 2892
rect 4326 2868 4330 2872
rect 4334 2868 4338 2872
rect 4310 2858 4314 2862
rect 4334 2858 4338 2862
rect 4278 2818 4282 2822
rect 4230 2728 4234 2732
rect 4238 2718 4242 2722
rect 4166 2658 4170 2662
rect 4190 2648 4194 2652
rect 4174 2638 4178 2642
rect 4158 2628 4162 2632
rect 4150 2598 4154 2602
rect 4182 2588 4186 2592
rect 4174 2558 4178 2562
rect 4126 2548 4130 2552
rect 4158 2548 4162 2552
rect 4206 2608 4210 2612
rect 4230 2588 4234 2592
rect 4262 2718 4266 2722
rect 4270 2708 4274 2712
rect 4374 2918 4378 2922
rect 4350 2808 4354 2812
rect 4334 2768 4338 2772
rect 4302 2758 4306 2762
rect 4310 2748 4314 2752
rect 4334 2738 4338 2742
rect 4286 2728 4290 2732
rect 4310 2728 4314 2732
rect 4326 2718 4330 2722
rect 4278 2698 4282 2702
rect 4326 2698 4330 2702
rect 4278 2678 4282 2682
rect 4262 2668 4266 2672
rect 4390 3008 4394 3012
rect 4426 3003 4430 3007
rect 4433 3003 4437 3007
rect 4454 2988 4458 2992
rect 4398 2958 4402 2962
rect 4414 2958 4418 2962
rect 4382 2738 4386 2742
rect 4374 2728 4378 2732
rect 4382 2718 4386 2722
rect 4406 2928 4410 2932
rect 4414 2928 4418 2932
rect 4446 2928 4450 2932
rect 4430 2918 4434 2922
rect 4414 2908 4418 2912
rect 4398 2858 4402 2862
rect 4426 2803 4430 2807
rect 4433 2803 4437 2807
rect 4414 2748 4418 2752
rect 4438 2748 4442 2752
rect 4414 2718 4418 2722
rect 4398 2688 4402 2692
rect 4390 2678 4394 2682
rect 4342 2668 4346 2672
rect 4374 2668 4378 2672
rect 4406 2678 4410 2682
rect 4310 2658 4314 2662
rect 4350 2658 4354 2662
rect 4262 2648 4266 2652
rect 4334 2648 4338 2652
rect 4390 2648 4394 2652
rect 4302 2628 4306 2632
rect 4318 2628 4322 2632
rect 4318 2598 4322 2602
rect 4254 2578 4258 2582
rect 4270 2578 4274 2582
rect 4310 2578 4314 2582
rect 4342 2578 4346 2582
rect 4382 2578 4386 2582
rect 4150 2538 4154 2542
rect 4174 2538 4178 2542
rect 4126 2528 4130 2532
rect 4158 2518 4162 2522
rect 4142 2498 4146 2502
rect 4102 2478 4106 2482
rect 4126 2478 4130 2482
rect 4126 2468 4130 2472
rect 4078 2458 4082 2462
rect 4086 2458 4090 2462
rect 4110 2458 4114 2462
rect 4054 2448 4058 2452
rect 4062 2428 4066 2432
rect 4046 2418 4050 2422
rect 4022 2368 4026 2372
rect 3990 2358 3994 2362
rect 4014 2358 4018 2362
rect 4038 2358 4042 2362
rect 3974 2348 3978 2352
rect 3990 2348 3994 2352
rect 3998 2348 4002 2352
rect 3982 2338 3986 2342
rect 3982 2308 3986 2312
rect 3974 2298 3978 2302
rect 3982 2258 3986 2262
rect 3950 2248 3954 2252
rect 3974 2198 3978 2202
rect 3974 2188 3978 2192
rect 3926 2178 3930 2182
rect 3934 2178 3938 2182
rect 3950 2168 3954 2172
rect 3958 2168 3962 2172
rect 3886 2148 3890 2152
rect 3910 2148 3914 2152
rect 3886 2138 3890 2142
rect 3886 2108 3890 2112
rect 3922 2103 3926 2107
rect 3929 2103 3933 2107
rect 3910 2098 3914 2102
rect 3902 2068 3906 2072
rect 3838 2058 3842 2062
rect 3846 2038 3850 2042
rect 3822 2028 3826 2032
rect 3878 2038 3882 2042
rect 3870 2018 3874 2022
rect 3902 1968 3906 1972
rect 3798 1918 3802 1922
rect 3950 1978 3954 1982
rect 3870 1928 3874 1932
rect 3878 1928 3882 1932
rect 3862 1918 3866 1922
rect 3806 1908 3810 1912
rect 3862 1908 3866 1912
rect 3814 1868 3818 1872
rect 3774 1848 3778 1852
rect 3790 1848 3794 1852
rect 3806 1858 3810 1862
rect 3830 1848 3834 1852
rect 3830 1808 3834 1812
rect 3870 1858 3874 1862
rect 3886 1918 3890 1922
rect 3942 1908 3946 1912
rect 3922 1903 3926 1907
rect 3929 1903 3933 1907
rect 3950 1898 3954 1902
rect 3990 2248 3994 2252
rect 3998 2248 4002 2252
rect 4094 2428 4098 2432
rect 4078 2388 4082 2392
rect 4054 2378 4058 2382
rect 4102 2418 4106 2422
rect 4134 2438 4138 2442
rect 4118 2418 4122 2422
rect 4038 2348 4042 2352
rect 4046 2348 4050 2352
rect 4030 2338 4034 2342
rect 4182 2528 4186 2532
rect 4166 2398 4170 2402
rect 4150 2388 4154 2392
rect 4126 2358 4130 2362
rect 4118 2348 4122 2352
rect 4110 2338 4114 2342
rect 4022 2308 4026 2312
rect 4022 2258 4026 2262
rect 4022 2248 4026 2252
rect 4006 2238 4010 2242
rect 4014 2238 4018 2242
rect 3990 2208 3994 2212
rect 3998 2208 4002 2212
rect 4014 2198 4018 2202
rect 3966 2138 3970 2142
rect 3982 2138 3986 2142
rect 4006 2118 4010 2122
rect 4014 2118 4018 2122
rect 3966 2098 3970 2102
rect 4070 2328 4074 2332
rect 4038 2248 4042 2252
rect 4078 2318 4082 2322
rect 4070 2288 4074 2292
rect 4078 2288 4082 2292
rect 4078 2268 4082 2272
rect 4086 2258 4090 2262
rect 4054 2188 4058 2192
rect 4086 2188 4090 2192
rect 4046 2148 4050 2152
rect 4062 2138 4066 2142
rect 4030 2118 4034 2122
rect 4030 2078 4034 2082
rect 4054 2078 4058 2082
rect 4046 2068 4050 2072
rect 4006 2058 4010 2062
rect 4022 2058 4026 2062
rect 4062 2058 4066 2062
rect 4046 2048 4050 2052
rect 3982 2038 3986 2042
rect 4030 2028 4034 2032
rect 3998 2008 4002 2012
rect 3982 1978 3986 1982
rect 3998 1958 4002 1962
rect 4014 1958 4018 1962
rect 4006 1928 4010 1932
rect 3966 1908 3970 1912
rect 3966 1878 3970 1882
rect 3926 1868 3930 1872
rect 3958 1868 3962 1872
rect 4014 1868 4018 1872
rect 3918 1858 3922 1862
rect 3878 1848 3882 1852
rect 3846 1838 3850 1842
rect 3870 1838 3874 1842
rect 3862 1828 3866 1832
rect 3838 1758 3842 1762
rect 3910 1818 3914 1822
rect 3878 1798 3882 1802
rect 3838 1748 3842 1752
rect 3870 1748 3874 1752
rect 3838 1738 3842 1742
rect 3798 1678 3802 1682
rect 3830 1658 3834 1662
rect 3766 1648 3770 1652
rect 3830 1648 3834 1652
rect 3758 1628 3762 1632
rect 3782 1578 3786 1582
rect 3694 1558 3698 1562
rect 3734 1558 3738 1562
rect 3678 1548 3682 1552
rect 3670 1538 3674 1542
rect 3702 1538 3706 1542
rect 3718 1538 3722 1542
rect 3694 1518 3698 1522
rect 3654 1488 3658 1492
rect 3638 1478 3642 1482
rect 3662 1478 3666 1482
rect 3646 1468 3650 1472
rect 3630 1458 3634 1462
rect 3622 1438 3626 1442
rect 3566 1428 3570 1432
rect 3590 1428 3594 1432
rect 3598 1358 3602 1362
rect 3638 1358 3642 1362
rect 3654 1458 3658 1462
rect 3678 1448 3682 1452
rect 3686 1428 3690 1432
rect 3654 1358 3658 1362
rect 3606 1348 3610 1352
rect 3630 1348 3634 1352
rect 3662 1348 3666 1352
rect 3750 1528 3754 1532
rect 3870 1698 3874 1702
rect 3854 1678 3858 1682
rect 3854 1628 3858 1632
rect 3846 1578 3850 1582
rect 3830 1568 3834 1572
rect 3854 1568 3858 1572
rect 3838 1558 3842 1562
rect 3790 1548 3794 1552
rect 3846 1538 3850 1542
rect 3822 1528 3826 1532
rect 3902 1748 3906 1752
rect 3950 1858 3954 1862
rect 3982 1858 3986 1862
rect 4022 1858 4026 1862
rect 3990 1848 3994 1852
rect 3990 1818 3994 1822
rect 3974 1778 3978 1782
rect 4006 1788 4010 1792
rect 3990 1768 3994 1772
rect 4006 1758 4010 1762
rect 3942 1748 3946 1752
rect 4038 1978 4042 1982
rect 4078 1988 4082 1992
rect 4102 2198 4106 2202
rect 4166 2378 4170 2382
rect 4294 2538 4298 2542
rect 4350 2538 4354 2542
rect 4278 2528 4282 2532
rect 4326 2528 4330 2532
rect 4350 2528 4354 2532
rect 4382 2528 4386 2532
rect 4198 2498 4202 2502
rect 4190 2458 4194 2462
rect 4190 2358 4194 2362
rect 4150 2348 4154 2352
rect 4174 2348 4178 2352
rect 4246 2468 4250 2472
rect 4254 2448 4258 2452
rect 4326 2498 4330 2502
rect 4326 2478 4330 2482
rect 4278 2468 4282 2472
rect 4286 2458 4290 2462
rect 4294 2458 4298 2462
rect 4318 2458 4322 2462
rect 4302 2448 4306 2452
rect 4310 2448 4314 2452
rect 4262 2428 4266 2432
rect 4262 2408 4266 2412
rect 4294 2388 4298 2392
rect 4254 2378 4258 2382
rect 4206 2368 4210 2372
rect 4198 2328 4202 2332
rect 4190 2318 4194 2322
rect 4134 2278 4138 2282
rect 4150 2268 4154 2272
rect 4134 2248 4138 2252
rect 4118 2148 4122 2152
rect 4102 2078 4106 2082
rect 4286 2348 4290 2352
rect 4222 2328 4226 2332
rect 4286 2328 4290 2332
rect 4270 2318 4274 2322
rect 4262 2298 4266 2302
rect 4230 2288 4234 2292
rect 4246 2288 4250 2292
rect 4238 2278 4242 2282
rect 4166 2258 4170 2262
rect 4174 2238 4178 2242
rect 4198 2208 4202 2212
rect 4254 2258 4258 2262
rect 4278 2258 4282 2262
rect 4286 2238 4290 2242
rect 4262 2208 4266 2212
rect 4310 2398 4314 2402
rect 4310 2358 4314 2362
rect 4366 2498 4370 2502
rect 4358 2478 4362 2482
rect 4358 2468 4362 2472
rect 4358 2438 4362 2442
rect 4342 2388 4346 2392
rect 4350 2378 4354 2382
rect 4310 2348 4314 2352
rect 4318 2278 4322 2282
rect 4310 2268 4314 2272
rect 4342 2298 4346 2302
rect 4374 2488 4378 2492
rect 4382 2478 4386 2482
rect 4374 2458 4378 2462
rect 4398 2558 4402 2562
rect 4398 2548 4402 2552
rect 4398 2538 4402 2542
rect 4374 2438 4378 2442
rect 4366 2358 4370 2362
rect 4446 2728 4450 2732
rect 4510 3038 4514 3042
rect 4494 3028 4498 3032
rect 4470 2978 4474 2982
rect 4470 2968 4474 2972
rect 4486 2968 4490 2972
rect 4462 2818 4466 2822
rect 4478 2958 4482 2962
rect 4486 2928 4490 2932
rect 4478 2918 4482 2922
rect 4518 3008 4522 3012
rect 4510 2958 4514 2962
rect 4502 2938 4506 2942
rect 4518 2938 4522 2942
rect 4526 2938 4530 2942
rect 4518 2928 4522 2932
rect 4726 3338 4730 3342
rect 4686 3328 4690 3332
rect 4710 3328 4714 3332
rect 4742 3328 4746 3332
rect 4710 3308 4714 3312
rect 4654 3298 4658 3302
rect 4662 3248 4666 3252
rect 4646 3228 4650 3232
rect 4734 3259 4738 3263
rect 4798 3338 4802 3342
rect 4830 3408 4834 3412
rect 4830 3348 4834 3352
rect 4798 3328 4802 3332
rect 4814 3328 4818 3332
rect 4830 3328 4834 3332
rect 4838 3328 4842 3332
rect 4790 3298 4794 3302
rect 4814 3298 4818 3302
rect 4790 3268 4794 3272
rect 4830 3268 4834 3272
rect 4838 3258 4842 3262
rect 4910 3648 4914 3652
rect 4886 3628 4890 3632
rect 4926 3628 4930 3632
rect 4862 3548 4866 3552
rect 4870 3448 4874 3452
rect 4926 3538 4930 3542
rect 4910 3518 4914 3522
rect 4910 3508 4914 3512
rect 4886 3388 4890 3392
rect 4878 3368 4882 3372
rect 4870 3348 4874 3352
rect 4910 3398 4914 3402
rect 4894 3358 4898 3362
rect 4870 3318 4874 3322
rect 4886 3328 4890 3332
rect 4870 3268 4874 3272
rect 4902 3278 4906 3282
rect 4942 3528 4946 3532
rect 4938 3503 4942 3507
rect 4945 3503 4949 3507
rect 4926 3488 4930 3492
rect 4950 3468 4954 3472
rect 4942 3358 4946 3362
rect 4990 3958 4994 3962
rect 5014 3958 5018 3962
rect 4990 3948 4994 3952
rect 5006 3948 5010 3952
rect 5014 3948 5018 3952
rect 4998 3938 5002 3942
rect 4990 3928 4994 3932
rect 4998 3898 5002 3902
rect 4990 3888 4994 3892
rect 4982 3858 4986 3862
rect 4998 3828 5002 3832
rect 4974 3798 4978 3802
rect 4990 3778 4994 3782
rect 4998 3778 5002 3782
rect 4990 3748 4994 3752
rect 4982 3738 4986 3742
rect 4974 3728 4978 3732
rect 4974 3718 4978 3722
rect 4990 3688 4994 3692
rect 4990 3648 4994 3652
rect 4982 3608 4986 3612
rect 5054 3947 5058 3951
rect 5038 3888 5042 3892
rect 5030 3858 5034 3862
rect 5094 4008 5098 4012
rect 5110 3998 5114 4002
rect 5102 3968 5106 3972
rect 5190 4298 5194 4302
rect 5238 4298 5242 4302
rect 5198 4288 5202 4292
rect 5182 4258 5186 4262
rect 5182 4228 5186 4232
rect 5166 4218 5170 4222
rect 5134 4178 5138 4182
rect 5150 4158 5154 4162
rect 5198 4268 5202 4272
rect 5278 4318 5282 4322
rect 5206 4238 5210 4242
rect 5190 4208 5194 4212
rect 5198 4198 5202 4202
rect 5190 4168 5194 4172
rect 5158 4148 5162 4152
rect 5174 4148 5178 4152
rect 5150 4138 5154 4142
rect 5198 4118 5202 4122
rect 5198 4108 5202 4112
rect 5134 4088 5138 4092
rect 5166 4088 5170 4092
rect 5182 4088 5186 4092
rect 5190 4078 5194 4082
rect 5166 4058 5170 4062
rect 5150 4038 5154 4042
rect 5134 4028 5138 4032
rect 5126 3988 5130 3992
rect 5118 3958 5122 3962
rect 5182 4018 5186 4022
rect 5190 4018 5194 4022
rect 5142 3958 5146 3962
rect 5174 3958 5178 3962
rect 5158 3948 5162 3952
rect 5190 4008 5194 4012
rect 5078 3938 5082 3942
rect 5150 3938 5154 3942
rect 5166 3938 5170 3942
rect 5190 3938 5194 3942
rect 5014 3798 5018 3802
rect 5054 3788 5058 3792
rect 5118 3898 5122 3902
rect 5142 3888 5146 3892
rect 5118 3868 5122 3872
rect 5174 3888 5178 3892
rect 5174 3878 5178 3882
rect 5150 3858 5154 3862
rect 5174 3858 5178 3862
rect 5190 3858 5194 3862
rect 5166 3848 5170 3852
rect 5134 3838 5138 3842
rect 5126 3808 5130 3812
rect 5110 3798 5114 3802
rect 5054 3778 5058 3782
rect 5094 3778 5098 3782
rect 5110 3778 5114 3782
rect 5078 3768 5082 3772
rect 5038 3728 5042 3732
rect 5014 3718 5018 3722
rect 5118 3768 5122 3772
rect 5110 3758 5114 3762
rect 5102 3688 5106 3692
rect 5006 3588 5010 3592
rect 5006 3568 5010 3572
rect 5030 3658 5034 3662
rect 5038 3648 5042 3652
rect 5078 3648 5082 3652
rect 5030 3638 5034 3642
rect 5054 3628 5058 3632
rect 4974 3548 4978 3552
rect 5022 3548 5026 3552
rect 4974 3528 4978 3532
rect 4974 3498 4978 3502
rect 5006 3528 5010 3532
rect 5038 3528 5042 3532
rect 5046 3518 5050 3522
rect 4990 3488 4994 3492
rect 5030 3488 5034 3492
rect 5038 3478 5042 3482
rect 5014 3468 5018 3472
rect 4982 3448 4986 3452
rect 4966 3418 4970 3422
rect 5022 3448 5026 3452
rect 5014 3408 5018 3412
rect 5006 3378 5010 3382
rect 4990 3368 4994 3372
rect 4966 3348 4970 3352
rect 4950 3328 4954 3332
rect 4966 3328 4970 3332
rect 4934 3318 4938 3322
rect 4938 3303 4942 3307
rect 4945 3303 4949 3307
rect 4982 3308 4986 3312
rect 4998 3308 5002 3312
rect 4966 3288 4970 3292
rect 4950 3278 4954 3282
rect 4942 3268 4946 3272
rect 4918 3258 4922 3262
rect 4934 3258 4938 3262
rect 4846 3248 4850 3252
rect 4862 3248 4866 3252
rect 4782 3228 4786 3232
rect 4806 3188 4810 3192
rect 4686 3178 4690 3182
rect 4806 3178 4810 3182
rect 4694 3158 4698 3162
rect 4726 3158 4730 3162
rect 4638 3148 4642 3152
rect 4646 3128 4650 3132
rect 4646 3118 4650 3122
rect 4814 3158 4818 3162
rect 4758 3148 4762 3152
rect 4854 3168 4858 3172
rect 4894 3158 4898 3162
rect 4862 3148 4866 3152
rect 4886 3148 4890 3152
rect 4726 3138 4730 3142
rect 4750 3138 4754 3142
rect 4790 3138 4794 3142
rect 4670 3088 4674 3092
rect 4598 3058 4602 3062
rect 4638 3048 4642 3052
rect 4654 3038 4658 3042
rect 4582 3008 4586 3012
rect 4558 2998 4562 3002
rect 4582 2948 4586 2952
rect 4550 2928 4554 2932
rect 4534 2918 4538 2922
rect 4566 2938 4570 2942
rect 4558 2898 4562 2902
rect 4590 2898 4594 2902
rect 4534 2878 4538 2882
rect 4566 2878 4570 2882
rect 4478 2848 4482 2852
rect 4542 2868 4546 2872
rect 4574 2868 4578 2872
rect 4598 2888 4602 2892
rect 4526 2858 4530 2862
rect 4582 2858 4586 2862
rect 4510 2838 4514 2842
rect 4510 2818 4514 2822
rect 4486 2808 4490 2812
rect 4734 3108 4738 3112
rect 4710 3098 4714 3102
rect 4758 3098 4762 3102
rect 4694 3058 4698 3062
rect 4686 2988 4690 2992
rect 4678 2948 4682 2952
rect 4662 2938 4666 2942
rect 4742 3088 4746 3092
rect 4718 3058 4722 3062
rect 4758 3058 4762 3062
rect 4774 3058 4778 3062
rect 4718 3048 4722 3052
rect 4766 3048 4770 3052
rect 4694 2978 4698 2982
rect 4702 2958 4706 2962
rect 4622 2928 4626 2932
rect 4694 2918 4698 2922
rect 4638 2858 4642 2862
rect 4678 2858 4682 2862
rect 4646 2818 4650 2822
rect 4614 2788 4618 2792
rect 4558 2758 4562 2762
rect 4574 2758 4578 2762
rect 4622 2768 4626 2772
rect 4478 2748 4482 2752
rect 4590 2748 4594 2752
rect 4478 2738 4482 2742
rect 4462 2688 4466 2692
rect 4526 2688 4530 2692
rect 4462 2658 4466 2662
rect 4510 2658 4514 2662
rect 4454 2648 4458 2652
rect 4426 2603 4430 2607
rect 4433 2603 4437 2607
rect 4470 2598 4474 2602
rect 4454 2578 4458 2582
rect 4446 2548 4450 2552
rect 4430 2538 4434 2542
rect 4422 2468 4426 2472
rect 4406 2448 4410 2452
rect 4462 2538 4466 2542
rect 4462 2478 4466 2482
rect 4486 2528 4490 2532
rect 4534 2668 4538 2672
rect 4526 2648 4530 2652
rect 4518 2548 4522 2552
rect 4510 2498 4514 2502
rect 4494 2478 4498 2482
rect 4478 2468 4482 2472
rect 4510 2468 4514 2472
rect 4446 2458 4450 2462
rect 4470 2458 4474 2462
rect 4462 2448 4466 2452
rect 4454 2428 4458 2432
rect 4382 2418 4386 2422
rect 4398 2418 4402 2422
rect 4430 2418 4434 2422
rect 4366 2348 4370 2352
rect 4426 2403 4430 2407
rect 4433 2403 4437 2407
rect 4398 2398 4402 2402
rect 4406 2368 4410 2372
rect 4398 2318 4402 2322
rect 4358 2268 4362 2272
rect 4334 2258 4338 2262
rect 4318 2248 4322 2252
rect 4350 2248 4354 2252
rect 4478 2418 4482 2422
rect 4494 2408 4498 2412
rect 4502 2388 4506 2392
rect 4486 2358 4490 2362
rect 4486 2348 4490 2352
rect 4510 2368 4514 2372
rect 4550 2738 4554 2742
rect 4582 2738 4586 2742
rect 4566 2728 4570 2732
rect 4550 2678 4554 2682
rect 4550 2668 4554 2672
rect 4582 2688 4586 2692
rect 4598 2598 4602 2602
rect 4542 2548 4546 2552
rect 4566 2528 4570 2532
rect 4534 2388 4538 2392
rect 4606 2568 4610 2572
rect 4670 2778 4674 2782
rect 4654 2738 4658 2742
rect 4622 2688 4626 2692
rect 4638 2708 4642 2712
rect 4670 2708 4674 2712
rect 4662 2668 4666 2672
rect 4630 2658 4634 2662
rect 4638 2588 4642 2592
rect 4622 2578 4626 2582
rect 4614 2548 4618 2552
rect 4614 2538 4618 2542
rect 4638 2518 4642 2522
rect 4646 2518 4650 2522
rect 4590 2498 4594 2502
rect 4622 2468 4626 2472
rect 4654 2468 4658 2472
rect 4630 2458 4634 2462
rect 4630 2448 4634 2452
rect 4574 2378 4578 2382
rect 4558 2368 4562 2372
rect 4526 2348 4530 2352
rect 4406 2258 4410 2262
rect 4398 2238 4402 2242
rect 4414 2238 4418 2242
rect 4358 2218 4362 2222
rect 4426 2203 4430 2207
rect 4433 2203 4437 2207
rect 4414 2198 4418 2202
rect 4270 2188 4274 2192
rect 4294 2188 4298 2192
rect 4302 2188 4306 2192
rect 4238 2158 4242 2162
rect 4174 2148 4178 2152
rect 4206 2148 4210 2152
rect 4254 2148 4258 2152
rect 4286 2148 4290 2152
rect 4310 2148 4314 2152
rect 4438 2148 4442 2152
rect 4142 2118 4146 2122
rect 4150 2068 4154 2072
rect 4142 2058 4146 2062
rect 4126 2038 4130 2042
rect 4166 2068 4170 2072
rect 4182 2138 4186 2142
rect 4246 2138 4250 2142
rect 4198 2108 4202 2112
rect 4214 2088 4218 2092
rect 4190 2078 4194 2082
rect 4198 2068 4202 2072
rect 4142 2048 4146 2052
rect 4158 2048 4162 2052
rect 4134 1998 4138 2002
rect 4094 1988 4098 1992
rect 4086 1978 4090 1982
rect 4110 1958 4114 1962
rect 4150 2028 4154 2032
rect 4054 1948 4058 1952
rect 4054 1938 4058 1942
rect 4070 1938 4074 1942
rect 4086 1938 4090 1942
rect 4094 1938 4098 1942
rect 4110 1938 4114 1942
rect 4126 1938 4130 1942
rect 4102 1918 4106 1922
rect 4070 1908 4074 1912
rect 4062 1848 4066 1852
rect 4062 1768 4066 1772
rect 4046 1758 4050 1762
rect 3918 1738 3922 1742
rect 3982 1738 3986 1742
rect 4062 1738 4066 1742
rect 3894 1728 3898 1732
rect 3902 1708 3906 1712
rect 3922 1703 3926 1707
rect 3929 1703 3933 1707
rect 3902 1678 3906 1682
rect 4038 1698 4042 1702
rect 4102 1878 4106 1882
rect 4110 1878 4114 1882
rect 4094 1858 4098 1862
rect 4110 1768 4114 1772
rect 4118 1728 4122 1732
rect 3950 1668 3954 1672
rect 4030 1668 4034 1672
rect 4094 1668 4098 1672
rect 3942 1658 3946 1662
rect 4014 1658 4018 1662
rect 4030 1658 4034 1662
rect 3998 1648 4002 1652
rect 4030 1648 4034 1652
rect 4086 1638 4090 1642
rect 3886 1568 3890 1572
rect 3910 1568 3914 1572
rect 3862 1558 3866 1562
rect 3878 1548 3882 1552
rect 3982 1608 3986 1612
rect 4038 1598 4042 1602
rect 4030 1578 4034 1582
rect 3982 1538 3986 1542
rect 3966 1528 3970 1532
rect 3902 1518 3906 1522
rect 3790 1478 3794 1482
rect 3854 1478 3858 1482
rect 3894 1478 3898 1482
rect 3790 1448 3794 1452
rect 3806 1448 3810 1452
rect 3790 1438 3794 1442
rect 3766 1398 3770 1402
rect 3750 1368 3754 1372
rect 3774 1358 3778 1362
rect 3870 1468 3874 1472
rect 3846 1448 3850 1452
rect 3838 1428 3842 1432
rect 3798 1408 3802 1412
rect 3822 1408 3826 1412
rect 3734 1348 3738 1352
rect 3766 1348 3770 1352
rect 3502 1338 3506 1342
rect 3558 1338 3562 1342
rect 3582 1338 3586 1342
rect 3678 1338 3682 1342
rect 3462 1278 3466 1282
rect 3478 1278 3482 1282
rect 3502 1278 3506 1282
rect 3470 1268 3474 1272
rect 3510 1268 3514 1272
rect 3542 1268 3546 1272
rect 3390 1218 3394 1222
rect 3510 1218 3514 1222
rect 3402 1203 3406 1207
rect 3409 1203 3413 1207
rect 3374 1198 3378 1202
rect 3526 1198 3530 1202
rect 3430 1188 3434 1192
rect 3374 1158 3378 1162
rect 3414 1158 3418 1162
rect 3406 1148 3410 1152
rect 3310 1138 3314 1142
rect 3358 1138 3362 1142
rect 3310 1118 3314 1122
rect 3326 1118 3330 1122
rect 3334 1118 3338 1122
rect 3302 1108 3306 1112
rect 3302 1078 3306 1082
rect 3294 1058 3298 1062
rect 3238 1028 3242 1032
rect 3334 1098 3338 1102
rect 3334 1068 3338 1072
rect 3374 1138 3378 1142
rect 3366 1098 3370 1102
rect 3366 1088 3370 1092
rect 3350 1068 3354 1072
rect 3558 1258 3562 1262
rect 3550 1228 3554 1232
rect 3590 1298 3594 1302
rect 3606 1298 3610 1302
rect 3622 1278 3626 1282
rect 3598 1258 3602 1262
rect 3566 1198 3570 1202
rect 3822 1388 3826 1392
rect 3798 1338 3802 1342
rect 3718 1328 3722 1332
rect 3694 1308 3698 1312
rect 3542 1188 3546 1192
rect 3654 1188 3658 1192
rect 3686 1188 3690 1192
rect 3550 1178 3554 1182
rect 3478 1158 3482 1162
rect 3518 1158 3522 1162
rect 3542 1158 3546 1162
rect 3606 1168 3610 1172
rect 3566 1158 3570 1162
rect 3438 1098 3442 1102
rect 3430 1068 3434 1072
rect 3326 1058 3330 1062
rect 3342 1058 3346 1062
rect 3390 1058 3394 1062
rect 3198 1018 3202 1022
rect 3318 1018 3322 1022
rect 3142 998 3146 1002
rect 3142 978 3146 982
rect 3094 968 3098 972
rect 3102 968 3106 972
rect 3174 958 3178 962
rect 3006 948 3010 952
rect 3078 948 3082 952
rect 3086 938 3090 942
rect 3142 938 3146 942
rect 2966 928 2970 932
rect 2982 928 2986 932
rect 2982 918 2986 922
rect 2926 858 2930 862
rect 2982 858 2986 862
rect 2910 828 2914 832
rect 2958 848 2962 852
rect 2974 848 2978 852
rect 2934 818 2938 822
rect 2878 778 2882 782
rect 2902 778 2906 782
rect 2862 768 2866 772
rect 2886 758 2890 762
rect 2702 738 2706 742
rect 2734 738 2738 742
rect 2782 738 2786 742
rect 2662 708 2666 712
rect 2622 668 2626 672
rect 2654 668 2658 672
rect 2686 698 2690 702
rect 2630 658 2634 662
rect 2646 658 2650 662
rect 2646 598 2650 602
rect 2662 568 2666 572
rect 2630 548 2634 552
rect 2606 528 2610 532
rect 2622 528 2626 532
rect 2646 528 2650 532
rect 2670 528 2674 532
rect 2654 518 2658 522
rect 2670 508 2674 512
rect 2774 728 2778 732
rect 2710 668 2714 672
rect 2742 668 2746 672
rect 2702 658 2706 662
rect 2710 638 2714 642
rect 2790 568 2794 572
rect 2782 548 2786 552
rect 2726 538 2730 542
rect 2718 518 2722 522
rect 2686 508 2690 512
rect 2670 478 2674 482
rect 2678 478 2682 482
rect 2734 488 2738 492
rect 2686 468 2690 472
rect 2702 468 2706 472
rect 2718 468 2722 472
rect 2630 459 2634 463
rect 2694 458 2698 462
rect 2606 448 2610 452
rect 2742 448 2746 452
rect 2774 538 2778 542
rect 2910 768 2914 772
rect 2982 838 2986 842
rect 2918 748 2922 752
rect 2830 738 2834 742
rect 2814 678 2818 682
rect 2838 678 2842 682
rect 2846 668 2850 672
rect 2814 658 2818 662
rect 2822 648 2826 652
rect 2806 598 2810 602
rect 2822 558 2826 562
rect 2806 538 2810 542
rect 2798 498 2802 502
rect 2822 488 2826 492
rect 2766 448 2770 452
rect 2782 448 2786 452
rect 2758 398 2762 402
rect 2614 378 2618 382
rect 2702 378 2706 382
rect 2702 358 2706 362
rect 2638 348 2642 352
rect 2726 348 2730 352
rect 2542 338 2546 342
rect 2614 338 2618 342
rect 2630 338 2634 342
rect 2670 338 2674 342
rect 2686 338 2690 342
rect 2598 328 2602 332
rect 2630 328 2634 332
rect 2662 328 2666 332
rect 2694 328 2698 332
rect 2526 268 2530 272
rect 2478 228 2482 232
rect 2462 208 2466 212
rect 2430 138 2434 142
rect 2438 138 2442 142
rect 2318 128 2322 132
rect 2350 128 2354 132
rect 2366 128 2370 132
rect 2286 108 2290 112
rect 2302 108 2306 112
rect 2254 88 2258 92
rect 2414 78 2418 82
rect 2326 68 2330 72
rect 2678 308 2682 312
rect 2638 288 2642 292
rect 2646 288 2650 292
rect 2606 268 2610 272
rect 2630 268 2634 272
rect 2590 258 2594 262
rect 2614 258 2618 262
rect 2710 288 2714 292
rect 2670 268 2674 272
rect 2718 268 2722 272
rect 2694 258 2698 262
rect 2598 248 2602 252
rect 2678 248 2682 252
rect 2710 248 2714 252
rect 2614 238 2618 242
rect 2542 148 2546 152
rect 2518 138 2522 142
rect 2566 138 2570 142
rect 2494 98 2498 102
rect 2646 218 2650 222
rect 2814 438 2818 442
rect 2814 358 2818 362
rect 2758 338 2762 342
rect 2766 338 2770 342
rect 2774 248 2778 252
rect 2726 168 2730 172
rect 2654 158 2658 162
rect 2638 148 2642 152
rect 2670 148 2674 152
rect 2518 78 2522 82
rect 2846 638 2850 642
rect 2926 728 2930 732
rect 2910 718 2914 722
rect 2890 703 2894 707
rect 2897 703 2901 707
rect 2878 688 2882 692
rect 2894 688 2898 692
rect 2870 678 2874 682
rect 2862 668 2866 672
rect 2958 748 2962 752
rect 2974 728 2978 732
rect 2990 718 2994 722
rect 2934 708 2938 712
rect 2982 708 2986 712
rect 2958 678 2962 682
rect 2966 668 2970 672
rect 2894 658 2898 662
rect 2862 648 2866 652
rect 2846 568 2850 572
rect 2854 568 2858 572
rect 2894 568 2898 572
rect 2894 558 2898 562
rect 2878 548 2882 552
rect 2838 538 2842 542
rect 2854 528 2858 532
rect 2870 528 2874 532
rect 2838 478 2842 482
rect 2838 438 2842 442
rect 2854 438 2858 442
rect 2890 503 2894 507
rect 2897 503 2901 507
rect 2878 498 2882 502
rect 2870 468 2874 472
rect 2870 438 2874 442
rect 2942 658 2946 662
rect 2934 568 2938 572
rect 2918 508 2922 512
rect 2894 458 2898 462
rect 2958 648 2962 652
rect 2966 638 2970 642
rect 2982 638 2986 642
rect 2966 618 2970 622
rect 3102 928 3106 932
rect 3094 888 3098 892
rect 3046 878 3050 882
rect 3070 878 3074 882
rect 3086 868 3090 872
rect 3014 858 3018 862
rect 3022 848 3026 852
rect 3046 858 3050 862
rect 3038 838 3042 842
rect 3062 788 3066 792
rect 3022 768 3026 772
rect 3030 768 3034 772
rect 3046 748 3050 752
rect 3054 748 3058 752
rect 3038 738 3042 742
rect 3014 728 3018 732
rect 3030 658 3034 662
rect 3062 698 3066 702
rect 3134 918 3138 922
rect 3142 888 3146 892
rect 3118 858 3122 862
rect 3134 858 3138 862
rect 3182 858 3186 862
rect 3078 848 3082 852
rect 3182 848 3186 852
rect 3118 838 3122 842
rect 3078 808 3082 812
rect 3086 788 3090 792
rect 3078 738 3082 742
rect 3078 698 3082 702
rect 3070 688 3074 692
rect 3078 648 3082 652
rect 3046 618 3050 622
rect 2998 608 3002 612
rect 3062 578 3066 582
rect 3030 558 3034 562
rect 3006 548 3010 552
rect 3038 548 3042 552
rect 2982 538 2986 542
rect 3054 508 3058 512
rect 3014 488 3018 492
rect 3022 488 3026 492
rect 2950 468 2954 472
rect 2974 468 2978 472
rect 2990 468 2994 472
rect 2910 448 2914 452
rect 2878 428 2882 432
rect 2846 368 2850 372
rect 2846 308 2850 312
rect 2830 298 2834 302
rect 2838 298 2842 302
rect 2822 278 2826 282
rect 2870 388 2874 392
rect 3030 458 3034 462
rect 2958 398 2962 402
rect 2990 398 2994 402
rect 2942 358 2946 362
rect 3022 438 3026 442
rect 3030 438 3034 442
rect 3038 398 3042 402
rect 3054 378 3058 382
rect 3062 368 3066 372
rect 3038 358 3042 362
rect 2902 348 2906 352
rect 3046 348 3050 352
rect 2982 338 2986 342
rect 2998 338 3002 342
rect 2862 328 2866 332
rect 2862 298 2866 302
rect 2846 268 2850 272
rect 2830 228 2834 232
rect 3046 338 3050 342
rect 3006 328 3010 332
rect 2878 318 2882 322
rect 2870 208 2874 212
rect 2854 198 2858 202
rect 2830 178 2834 182
rect 2814 158 2818 162
rect 2846 168 2850 172
rect 2846 148 2850 152
rect 2862 158 2866 162
rect 2890 303 2894 307
rect 2897 303 2901 307
rect 3030 318 3034 322
rect 2958 298 2962 302
rect 3022 298 3026 302
rect 2926 288 2930 292
rect 2918 278 2922 282
rect 2990 278 2994 282
rect 2942 268 2946 272
rect 2902 258 2906 262
rect 2886 248 2890 252
rect 2942 228 2946 232
rect 2918 218 2922 222
rect 2894 198 2898 202
rect 2934 148 2938 152
rect 2662 138 2666 142
rect 2710 138 2714 142
rect 2742 138 2746 142
rect 2750 138 2754 142
rect 2878 138 2882 142
rect 2926 138 2930 142
rect 2718 128 2722 132
rect 2710 108 2714 112
rect 2702 98 2706 102
rect 2886 128 2890 132
rect 2782 118 2786 122
rect 2910 118 2914 122
rect 2890 103 2894 107
rect 2897 103 2901 107
rect 2926 98 2930 102
rect 2918 88 2922 92
rect 2742 78 2746 82
rect 2886 78 2890 82
rect 2894 78 2898 82
rect 2502 68 2506 72
rect 2558 68 2562 72
rect 2574 68 2578 72
rect 2646 68 2650 72
rect 2742 68 2746 72
rect 2838 68 2842 72
rect 3022 268 3026 272
rect 3006 218 3010 222
rect 3006 178 3010 182
rect 3078 508 3082 512
rect 3070 338 3074 342
rect 3094 758 3098 762
rect 3166 738 3170 742
rect 3150 718 3154 722
rect 3142 688 3146 692
rect 3110 678 3114 682
rect 3118 668 3122 672
rect 3126 658 3130 662
rect 3142 658 3146 662
rect 3102 638 3106 642
rect 3094 528 3098 532
rect 3166 648 3170 652
rect 3118 638 3122 642
rect 3310 958 3314 962
rect 3318 958 3322 962
rect 3278 948 3282 952
rect 3246 938 3250 942
rect 3286 938 3290 942
rect 3254 878 3258 882
rect 3310 888 3314 892
rect 3270 858 3274 862
rect 3206 848 3210 852
rect 3206 828 3210 832
rect 3238 798 3242 802
rect 3206 788 3210 792
rect 3230 758 3234 762
rect 3358 938 3362 942
rect 3366 888 3370 892
rect 3402 1003 3406 1007
rect 3409 1003 3413 1007
rect 3510 1138 3514 1142
rect 3502 1128 3506 1132
rect 3454 1108 3458 1112
rect 3494 1098 3498 1102
rect 3486 1088 3490 1092
rect 3462 1028 3466 1032
rect 3462 998 3466 1002
rect 3446 948 3450 952
rect 3470 948 3474 952
rect 3486 948 3490 952
rect 3438 928 3442 932
rect 3478 938 3482 942
rect 3510 988 3514 992
rect 3574 1148 3578 1152
rect 3534 1078 3538 1082
rect 3574 1138 3578 1142
rect 3558 1118 3562 1122
rect 3566 1088 3570 1092
rect 3534 1058 3538 1062
rect 3542 1058 3546 1062
rect 3526 1048 3530 1052
rect 3550 1048 3554 1052
rect 3598 1148 3602 1152
rect 3638 1158 3642 1162
rect 3606 1138 3610 1142
rect 3622 1118 3626 1122
rect 3654 1118 3658 1122
rect 3630 1088 3634 1092
rect 3662 1088 3666 1092
rect 3590 1078 3594 1082
rect 3630 1078 3634 1082
rect 3646 1078 3650 1082
rect 3622 1068 3626 1072
rect 3726 1258 3730 1262
rect 3710 1248 3714 1252
rect 3742 1328 3746 1332
rect 3742 1258 3746 1262
rect 3734 1238 3738 1242
rect 3726 1188 3730 1192
rect 3710 1148 3714 1152
rect 3718 1088 3722 1092
rect 3670 1068 3674 1072
rect 3686 1068 3690 1072
rect 3638 1058 3642 1062
rect 3638 1048 3642 1052
rect 3590 1018 3594 1022
rect 3582 998 3586 1002
rect 3542 978 3546 982
rect 3622 998 3626 1002
rect 3518 938 3522 942
rect 3550 938 3554 942
rect 3574 938 3578 942
rect 3590 938 3594 942
rect 3606 938 3610 942
rect 3622 938 3626 942
rect 3518 928 3522 932
rect 3502 908 3506 912
rect 3494 888 3498 892
rect 3382 878 3386 882
rect 3438 878 3442 882
rect 3462 878 3466 882
rect 3358 868 3362 872
rect 3390 868 3394 872
rect 3430 868 3434 872
rect 3454 868 3458 872
rect 3486 868 3490 872
rect 3406 858 3410 862
rect 3462 858 3466 862
rect 3494 858 3498 862
rect 3350 848 3354 852
rect 3486 848 3490 852
rect 3358 838 3362 842
rect 3402 803 3406 807
rect 3409 803 3413 807
rect 3318 798 3322 802
rect 3310 778 3314 782
rect 3462 778 3466 782
rect 3334 768 3338 772
rect 3222 748 3226 752
rect 3246 748 3250 752
rect 3270 748 3274 752
rect 3302 748 3306 752
rect 3206 718 3210 722
rect 3198 658 3202 662
rect 3190 648 3194 652
rect 3174 628 3178 632
rect 3182 628 3186 632
rect 3134 568 3138 572
rect 3182 608 3186 612
rect 3230 588 3234 592
rect 3198 568 3202 572
rect 3126 528 3130 532
rect 3174 498 3178 502
rect 3382 758 3386 762
rect 3446 758 3450 762
rect 3358 748 3362 752
rect 3446 748 3450 752
rect 3334 738 3338 742
rect 3478 738 3482 742
rect 3318 728 3322 732
rect 3302 698 3306 702
rect 3286 688 3290 692
rect 3254 638 3258 642
rect 3214 528 3218 532
rect 3158 488 3162 492
rect 3182 488 3186 492
rect 3110 478 3114 482
rect 3102 468 3106 472
rect 3166 468 3170 472
rect 3110 458 3114 462
rect 3086 308 3090 312
rect 3054 298 3058 302
rect 3062 298 3066 302
rect 3070 278 3074 282
rect 3086 248 3090 252
rect 3102 308 3106 312
rect 3118 428 3122 432
rect 3158 428 3162 432
rect 3134 398 3138 402
rect 3206 468 3210 472
rect 3214 458 3218 462
rect 3214 368 3218 372
rect 3206 358 3210 362
rect 3246 468 3250 472
rect 3238 388 3242 392
rect 3222 348 3226 352
rect 3158 328 3162 332
rect 3110 278 3114 282
rect 3118 278 3122 282
rect 3158 268 3162 272
rect 3198 338 3202 342
rect 3214 288 3218 292
rect 3222 278 3226 282
rect 3174 258 3178 262
rect 3094 218 3098 222
rect 3062 198 3066 202
rect 3070 158 3074 162
rect 3086 158 3090 162
rect 3118 248 3122 252
rect 3182 248 3186 252
rect 3206 248 3210 252
rect 3222 248 3226 252
rect 3118 238 3122 242
rect 3142 218 3146 222
rect 3110 158 3114 162
rect 2990 148 2994 152
rect 3054 148 3058 152
rect 3102 148 3106 152
rect 3062 138 3066 142
rect 3110 138 3114 142
rect 3014 108 3018 112
rect 3110 98 3114 102
rect 3126 88 3130 92
rect 3214 208 3218 212
rect 3158 188 3162 192
rect 3230 228 3234 232
rect 3222 168 3226 172
rect 3230 158 3234 162
rect 3214 148 3218 152
rect 3158 138 3162 142
rect 3174 138 3178 142
rect 3142 98 3146 102
rect 3030 78 3034 82
rect 3054 78 3058 82
rect 3134 78 3138 82
rect 3198 78 3202 82
rect 2958 68 2962 72
rect 3182 68 3186 72
rect 2126 58 2130 62
rect 2158 58 2162 62
rect 2374 58 2378 62
rect 2486 58 2490 62
rect 2550 58 2554 62
rect 2566 58 2570 62
rect 2646 58 2650 62
rect 2734 58 2738 62
rect 2830 58 2834 62
rect 2894 58 2898 62
rect 2966 58 2970 62
rect 3262 628 3266 632
rect 3278 558 3282 562
rect 3278 508 3282 512
rect 3302 598 3306 602
rect 3302 548 3306 552
rect 3294 538 3298 542
rect 3310 528 3314 532
rect 3302 488 3306 492
rect 3286 478 3290 482
rect 3310 478 3314 482
rect 3430 728 3434 732
rect 3406 718 3410 722
rect 3422 718 3426 722
rect 3390 678 3394 682
rect 3494 758 3498 762
rect 3526 888 3530 892
rect 3510 848 3514 852
rect 3542 878 3546 882
rect 3534 798 3538 802
rect 3710 1068 3714 1072
rect 3814 1318 3818 1322
rect 3806 1308 3810 1312
rect 3758 1288 3762 1292
rect 3782 1278 3786 1282
rect 3806 1288 3810 1292
rect 3758 1268 3762 1272
rect 3822 1308 3826 1312
rect 3854 1308 3858 1312
rect 3838 1298 3842 1302
rect 3830 1288 3834 1292
rect 3822 1268 3826 1272
rect 3846 1268 3850 1272
rect 3766 1238 3770 1242
rect 3766 1228 3770 1232
rect 3790 1228 3794 1232
rect 3886 1438 3890 1442
rect 3922 1503 3926 1507
rect 3929 1503 3933 1507
rect 3910 1478 3914 1482
rect 4070 1558 4074 1562
rect 4046 1538 4050 1542
rect 4062 1518 4066 1522
rect 4030 1498 4034 1502
rect 3974 1488 3978 1492
rect 4046 1488 4050 1492
rect 3958 1438 3962 1442
rect 3958 1428 3962 1432
rect 3910 1328 3914 1332
rect 3922 1303 3926 1307
rect 3929 1303 3933 1307
rect 3902 1288 3906 1292
rect 3982 1478 3986 1482
rect 3982 1468 3986 1472
rect 3974 1308 3978 1312
rect 3974 1268 3978 1272
rect 3846 1258 3850 1262
rect 3862 1258 3866 1262
rect 3878 1238 3882 1242
rect 3918 1248 3922 1252
rect 3846 1228 3850 1232
rect 3894 1228 3898 1232
rect 3814 1198 3818 1202
rect 3926 1218 3930 1222
rect 3782 1188 3786 1192
rect 3750 1168 3754 1172
rect 3838 1158 3842 1162
rect 3742 1108 3746 1112
rect 3958 1168 3962 1172
rect 3766 1148 3770 1152
rect 3782 1148 3786 1152
rect 3806 1118 3810 1122
rect 3822 1118 3826 1122
rect 3806 1088 3810 1092
rect 3758 1078 3762 1082
rect 3806 1078 3810 1082
rect 3678 1058 3682 1062
rect 3710 1058 3714 1062
rect 3758 1068 3762 1072
rect 3742 1018 3746 1022
rect 3686 988 3690 992
rect 3854 1108 3858 1112
rect 3966 1148 3970 1152
rect 3922 1103 3926 1107
rect 3929 1103 3933 1107
rect 3958 1098 3962 1102
rect 3902 1078 3906 1082
rect 3870 1068 3874 1072
rect 3774 1058 3778 1062
rect 3806 1058 3810 1062
rect 3822 1058 3826 1062
rect 3822 1038 3826 1042
rect 3766 998 3770 1002
rect 3782 998 3786 1002
rect 3734 958 3738 962
rect 3758 958 3762 962
rect 3670 948 3674 952
rect 3750 948 3754 952
rect 3734 938 3738 942
rect 3670 918 3674 922
rect 3726 918 3730 922
rect 3750 918 3754 922
rect 3654 898 3658 902
rect 3718 898 3722 902
rect 3774 988 3778 992
rect 3782 988 3786 992
rect 3782 968 3786 972
rect 3798 958 3802 962
rect 3830 1008 3834 1012
rect 4030 1458 4034 1462
rect 4054 1438 4058 1442
rect 4062 1418 4066 1422
rect 4014 1408 4018 1412
rect 4046 1408 4050 1412
rect 4006 1368 4010 1372
rect 4102 1558 4106 1562
rect 4102 1538 4106 1542
rect 4142 1908 4146 1912
rect 4158 1948 4162 1952
rect 4238 2088 4242 2092
rect 4238 2068 4242 2072
rect 4230 2048 4234 2052
rect 4222 2028 4226 2032
rect 4222 1998 4226 2002
rect 4198 1978 4202 1982
rect 4198 1968 4202 1972
rect 4190 1948 4194 1952
rect 4174 1898 4178 1902
rect 4182 1898 4186 1902
rect 4214 1888 4218 1892
rect 4206 1878 4210 1882
rect 4150 1868 4154 1872
rect 4190 1868 4194 1872
rect 4158 1858 4162 1862
rect 4174 1838 4178 1842
rect 4166 1808 4170 1812
rect 4214 1858 4218 1862
rect 4214 1818 4218 1822
rect 4198 1788 4202 1792
rect 4182 1758 4186 1762
rect 4246 1868 4250 1872
rect 4286 2138 4290 2142
rect 4382 2138 4386 2142
rect 4342 2118 4346 2122
rect 4286 2108 4290 2112
rect 4302 2088 4306 2092
rect 4262 1948 4266 1952
rect 4334 2078 4338 2082
rect 4302 1968 4306 1972
rect 4374 2108 4378 2112
rect 4390 2108 4394 2112
rect 4358 2088 4362 2092
rect 4350 2068 4354 2072
rect 4350 2038 4354 2042
rect 4454 2248 4458 2252
rect 4486 2298 4490 2302
rect 4470 2278 4474 2282
rect 4502 2278 4506 2282
rect 4478 2268 4482 2272
rect 4462 2168 4466 2172
rect 4462 2128 4466 2132
rect 4470 2128 4474 2132
rect 4446 2098 4450 2102
rect 4446 2088 4450 2092
rect 4462 2088 4466 2092
rect 4406 2068 4410 2072
rect 4366 2038 4370 2042
rect 4358 1998 4362 2002
rect 4310 1958 4314 1962
rect 4342 1958 4346 1962
rect 4318 1948 4322 1952
rect 4366 1948 4370 1952
rect 4398 2058 4402 2062
rect 4470 2078 4474 2082
rect 4526 2248 4530 2252
rect 4526 2238 4530 2242
rect 4518 2218 4522 2222
rect 4494 2158 4498 2162
rect 4502 2158 4506 2162
rect 4550 2318 4554 2322
rect 4542 2278 4546 2282
rect 4550 2268 4554 2272
rect 4582 2358 4586 2362
rect 4654 2368 4658 2372
rect 4686 2768 4690 2772
rect 4694 2768 4698 2772
rect 4710 2788 4714 2792
rect 4686 2688 4690 2692
rect 4678 2658 4682 2662
rect 4774 3028 4778 3032
rect 4798 3038 4802 3042
rect 4782 2998 4786 3002
rect 4894 3138 4898 3142
rect 4870 3128 4874 3132
rect 4838 3108 4842 3112
rect 4838 3098 4842 3102
rect 4854 3098 4858 3102
rect 4894 3108 4898 3112
rect 4910 3108 4914 3112
rect 4870 3088 4874 3092
rect 4886 3048 4890 3052
rect 4886 2998 4890 3002
rect 4822 2958 4826 2962
rect 4870 2958 4874 2962
rect 4734 2948 4738 2952
rect 4782 2948 4786 2952
rect 4830 2938 4834 2942
rect 4758 2928 4762 2932
rect 4902 3088 4906 3092
rect 4918 3098 4922 3102
rect 4902 3048 4906 3052
rect 4910 3048 4914 3052
rect 4918 3038 4922 3042
rect 4966 3228 4970 3232
rect 4990 3208 4994 3212
rect 4990 3188 4994 3192
rect 4934 3148 4938 3152
rect 4974 3128 4978 3132
rect 4938 3103 4942 3107
rect 4945 3103 4949 3107
rect 4966 3098 4970 3102
rect 5038 3448 5042 3452
rect 5030 3398 5034 3402
rect 5038 3278 5042 3282
rect 5038 3208 5042 3212
rect 5030 3198 5034 3202
rect 5094 3558 5098 3562
rect 5078 3478 5082 3482
rect 5086 3468 5090 3472
rect 5150 3788 5154 3792
rect 5158 3768 5162 3772
rect 5126 3748 5130 3752
rect 5126 3728 5130 3732
rect 5142 3718 5146 3722
rect 5134 3698 5138 3702
rect 5166 3718 5170 3722
rect 5182 3728 5186 3732
rect 5158 3698 5162 3702
rect 5174 3698 5178 3702
rect 5150 3688 5154 3692
rect 5142 3678 5146 3682
rect 5126 3658 5130 3662
rect 5110 3648 5114 3652
rect 5142 3648 5146 3652
rect 5118 3638 5122 3642
rect 5142 3638 5146 3642
rect 5150 3618 5154 3622
rect 5182 3668 5186 3672
rect 5166 3598 5170 3602
rect 5158 3558 5162 3562
rect 5150 3548 5154 3552
rect 5134 3518 5138 3522
rect 5102 3378 5106 3382
rect 5102 3368 5106 3372
rect 5062 3338 5066 3342
rect 5054 3328 5058 3332
rect 5102 3318 5106 3322
rect 5070 3288 5074 3292
rect 5062 3198 5066 3202
rect 5054 3158 5058 3162
rect 4998 3148 5002 3152
rect 4934 3068 4938 3072
rect 4998 3068 5002 3072
rect 4942 3058 4946 3062
rect 4926 3028 4930 3032
rect 4958 3028 4962 3032
rect 4902 2978 4906 2982
rect 4910 2978 4914 2982
rect 4846 2938 4850 2942
rect 4878 2938 4882 2942
rect 4838 2918 4842 2922
rect 4798 2878 4802 2882
rect 4750 2868 4754 2872
rect 4734 2768 4738 2772
rect 4750 2758 4754 2762
rect 4862 2928 4866 2932
rect 4854 2908 4858 2912
rect 4838 2868 4842 2872
rect 4878 2898 4882 2902
rect 4862 2878 4866 2882
rect 4782 2858 4786 2862
rect 4806 2858 4810 2862
rect 4798 2848 4802 2852
rect 4830 2848 4834 2852
rect 4774 2838 4778 2842
rect 4806 2798 4810 2802
rect 4790 2768 4794 2772
rect 4766 2748 4770 2752
rect 4790 2748 4794 2752
rect 4790 2728 4794 2732
rect 4774 2718 4778 2722
rect 4742 2708 4746 2712
rect 4702 2628 4706 2632
rect 4686 2598 4690 2602
rect 4670 2538 4674 2542
rect 4710 2618 4714 2622
rect 4758 2688 4762 2692
rect 4782 2688 4786 2692
rect 4830 2788 4834 2792
rect 4886 2868 4890 2872
rect 4942 2948 4946 2952
rect 4974 3048 4978 3052
rect 4998 3048 5002 3052
rect 4966 2998 4970 3002
rect 4990 2988 4994 2992
rect 4966 2968 4970 2972
rect 4934 2938 4938 2942
rect 4982 2928 4986 2932
rect 4942 2918 4946 2922
rect 4938 2903 4942 2907
rect 4945 2903 4949 2907
rect 4950 2858 4954 2862
rect 4990 2868 4994 2872
rect 4958 2838 4962 2842
rect 4942 2828 4946 2832
rect 4878 2778 4882 2782
rect 4854 2768 4858 2772
rect 4918 2768 4922 2772
rect 4974 2768 4978 2772
rect 4902 2758 4906 2762
rect 4926 2758 4930 2762
rect 4902 2748 4906 2752
rect 4926 2748 4930 2752
rect 4862 2728 4866 2732
rect 4918 2728 4922 2732
rect 4854 2718 4858 2722
rect 4838 2678 4842 2682
rect 4870 2708 4874 2712
rect 4966 2728 4970 2732
rect 4958 2718 4962 2722
rect 4918 2708 4922 2712
rect 4938 2703 4942 2707
rect 4945 2703 4949 2707
rect 4894 2698 4898 2702
rect 4910 2688 4914 2692
rect 4902 2678 4906 2682
rect 5030 3138 5034 3142
rect 5046 3138 5050 3142
rect 5102 3248 5106 3252
rect 5086 3218 5090 3222
rect 5142 3468 5146 3472
rect 5158 3528 5162 3532
rect 5230 4188 5234 4192
rect 5222 4158 5226 4162
rect 5238 4148 5242 4152
rect 5214 4138 5218 4142
rect 5222 4098 5226 4102
rect 5230 4038 5234 4042
rect 5222 3838 5226 3842
rect 5246 4138 5250 4142
rect 5262 4178 5266 4182
rect 5278 4158 5282 4162
rect 5270 4068 5274 4072
rect 5270 3938 5274 3942
rect 5254 3858 5258 3862
rect 5222 3738 5226 3742
rect 5206 3678 5210 3682
rect 5206 3648 5210 3652
rect 5198 3538 5202 3542
rect 5190 3518 5194 3522
rect 5182 3468 5186 3472
rect 5126 3448 5130 3452
rect 5126 3438 5130 3442
rect 5134 3428 5138 3432
rect 5118 3338 5122 3342
rect 5126 3338 5130 3342
rect 5126 3328 5130 3332
rect 5118 3268 5122 3272
rect 5118 3228 5122 3232
rect 5118 3218 5122 3222
rect 5078 3158 5082 3162
rect 5094 3158 5098 3162
rect 5110 3158 5114 3162
rect 5126 3158 5130 3162
rect 5038 3128 5042 3132
rect 5054 3128 5058 3132
rect 5078 3128 5082 3132
rect 5094 3108 5098 3112
rect 5046 3078 5050 3082
rect 5078 3078 5082 3082
rect 5014 3008 5018 3012
rect 5022 2998 5026 3002
rect 5110 3128 5114 3132
rect 5118 3108 5122 3112
rect 5126 3068 5130 3072
rect 5110 3058 5114 3062
rect 5094 3008 5098 3012
rect 5102 3008 5106 3012
rect 5102 2998 5106 3002
rect 5094 2958 5098 2962
rect 5030 2948 5034 2952
rect 5126 2988 5130 2992
rect 5118 2888 5122 2892
rect 5022 2878 5026 2882
rect 5078 2878 5082 2882
rect 5062 2858 5066 2862
rect 5038 2818 5042 2822
rect 5054 2808 5058 2812
rect 5054 2788 5058 2792
rect 5038 2768 5042 2772
rect 5014 2758 5018 2762
rect 5022 2748 5026 2752
rect 4998 2678 5002 2682
rect 4878 2668 4882 2672
rect 4910 2668 4914 2672
rect 4942 2668 4946 2672
rect 4766 2658 4770 2662
rect 4726 2648 4730 2652
rect 4838 2648 4842 2652
rect 4718 2608 4722 2612
rect 4766 2608 4770 2612
rect 4718 2578 4722 2582
rect 4710 2538 4714 2542
rect 4702 2508 4706 2512
rect 4710 2488 4714 2492
rect 4694 2478 4698 2482
rect 4678 2468 4682 2472
rect 4686 2468 4690 2472
rect 4862 2628 4866 2632
rect 4790 2578 4794 2582
rect 4806 2568 4810 2572
rect 4766 2558 4770 2562
rect 4790 2558 4794 2562
rect 4814 2558 4818 2562
rect 4782 2538 4786 2542
rect 4750 2518 4754 2522
rect 4782 2518 4786 2522
rect 4734 2498 4738 2502
rect 4774 2478 4778 2482
rect 4790 2478 4794 2482
rect 4798 2468 4802 2472
rect 4934 2648 4938 2652
rect 4942 2628 4946 2632
rect 4902 2598 4906 2602
rect 5030 2728 5034 2732
rect 4918 2568 4922 2572
rect 5014 2568 5018 2572
rect 4886 2558 4890 2562
rect 4910 2558 4914 2562
rect 4870 2538 4874 2542
rect 4990 2558 4994 2562
rect 4926 2548 4930 2552
rect 4958 2548 4962 2552
rect 4838 2498 4842 2502
rect 4902 2518 4906 2522
rect 4870 2488 4874 2492
rect 4886 2488 4890 2492
rect 4694 2458 4698 2462
rect 4766 2458 4770 2462
rect 4750 2448 4754 2452
rect 4686 2378 4690 2382
rect 4734 2358 4738 2362
rect 4638 2348 4642 2352
rect 4662 2348 4666 2352
rect 4702 2348 4706 2352
rect 4606 2338 4610 2342
rect 4662 2338 4666 2342
rect 4678 2338 4682 2342
rect 4710 2338 4714 2342
rect 4726 2338 4730 2342
rect 4542 2258 4546 2262
rect 4574 2258 4578 2262
rect 4590 2258 4594 2262
rect 4550 2248 4554 2252
rect 4566 2248 4570 2252
rect 4542 2158 4546 2162
rect 4534 2128 4538 2132
rect 4526 2118 4530 2122
rect 4510 2108 4514 2112
rect 4486 2078 4490 2082
rect 4494 2078 4498 2082
rect 4590 2218 4594 2222
rect 4574 2148 4578 2152
rect 4670 2328 4674 2332
rect 4678 2328 4682 2332
rect 4718 2328 4722 2332
rect 4686 2318 4690 2322
rect 4702 2318 4706 2322
rect 4606 2248 4610 2252
rect 4686 2288 4690 2292
rect 4718 2268 4722 2272
rect 4790 2448 4794 2452
rect 4806 2448 4810 2452
rect 4782 2378 4786 2382
rect 4814 2368 4818 2372
rect 4926 2528 4930 2532
rect 4934 2518 4938 2522
rect 4926 2508 4930 2512
rect 4938 2503 4942 2507
rect 4945 2503 4949 2507
rect 4934 2478 4938 2482
rect 4942 2458 4946 2462
rect 4966 2538 4970 2542
rect 4990 2538 4994 2542
rect 4966 2518 4970 2522
rect 4974 2498 4978 2502
rect 4926 2448 4930 2452
rect 4958 2448 4962 2452
rect 4918 2438 4922 2442
rect 4894 2428 4898 2432
rect 4910 2428 4914 2432
rect 4886 2378 4890 2382
rect 4798 2348 4802 2352
rect 4758 2318 4762 2322
rect 4766 2318 4770 2322
rect 4782 2318 4786 2322
rect 4774 2308 4778 2312
rect 4766 2298 4770 2302
rect 4758 2288 4762 2292
rect 4750 2278 4754 2282
rect 4814 2328 4818 2332
rect 4902 2328 4906 2332
rect 4838 2318 4842 2322
rect 4846 2308 4850 2312
rect 4838 2298 4842 2302
rect 4814 2288 4818 2292
rect 4822 2288 4826 2292
rect 4830 2288 4834 2292
rect 4854 2288 4858 2292
rect 4734 2258 4738 2262
rect 4678 2248 4682 2252
rect 4734 2228 4738 2232
rect 4694 2218 4698 2222
rect 4654 2188 4658 2192
rect 4614 2148 4618 2152
rect 4598 2128 4602 2132
rect 4590 2098 4594 2102
rect 4662 2168 4666 2172
rect 4670 2158 4674 2162
rect 4646 2138 4650 2142
rect 4678 2148 4682 2152
rect 4622 2118 4626 2122
rect 4678 2118 4682 2122
rect 4630 2108 4634 2112
rect 4646 2108 4650 2112
rect 4622 2078 4626 2082
rect 4542 2068 4546 2072
rect 4566 2068 4570 2072
rect 4614 2068 4618 2072
rect 4486 2058 4490 2062
rect 4518 2058 4522 2062
rect 4542 2058 4546 2062
rect 4406 2048 4410 2052
rect 4486 2048 4490 2052
rect 4494 2038 4498 2042
rect 4486 2018 4490 2022
rect 4426 2003 4430 2007
rect 4433 2003 4437 2007
rect 4478 1978 4482 1982
rect 4270 1938 4274 1942
rect 4286 1898 4290 1902
rect 4342 1898 4346 1902
rect 4294 1888 4298 1892
rect 4278 1868 4282 1872
rect 4414 1898 4418 1902
rect 4446 1898 4450 1902
rect 4470 1898 4474 1902
rect 4366 1868 4370 1872
rect 4390 1868 4394 1872
rect 4414 1868 4418 1872
rect 4414 1858 4418 1862
rect 4254 1848 4258 1852
rect 4406 1848 4410 1852
rect 4342 1838 4346 1842
rect 4230 1828 4234 1832
rect 4238 1828 4242 1832
rect 4262 1808 4266 1812
rect 4246 1758 4250 1762
rect 4134 1738 4138 1742
rect 4134 1708 4138 1712
rect 4166 1698 4170 1702
rect 4198 1738 4202 1742
rect 4198 1718 4202 1722
rect 4206 1708 4210 1712
rect 4238 1728 4242 1732
rect 4214 1688 4218 1692
rect 4230 1688 4234 1692
rect 4174 1678 4178 1682
rect 4222 1678 4226 1682
rect 4158 1668 4162 1672
rect 4198 1668 4202 1672
rect 4214 1668 4218 1672
rect 4158 1658 4162 1662
rect 4174 1658 4178 1662
rect 4206 1658 4210 1662
rect 4190 1648 4194 1652
rect 4134 1608 4138 1612
rect 4238 1648 4242 1652
rect 4230 1598 4234 1602
rect 4166 1588 4170 1592
rect 4222 1588 4226 1592
rect 4190 1578 4194 1582
rect 4174 1568 4178 1572
rect 4230 1568 4234 1572
rect 4254 1688 4258 1692
rect 4294 1788 4298 1792
rect 4366 1788 4370 1792
rect 4278 1768 4282 1772
rect 4270 1748 4274 1752
rect 4286 1748 4290 1752
rect 4382 1778 4386 1782
rect 4334 1758 4338 1762
rect 4278 1738 4282 1742
rect 4270 1718 4274 1722
rect 4286 1668 4290 1672
rect 4254 1658 4258 1662
rect 4270 1648 4274 1652
rect 4262 1578 4266 1582
rect 4254 1568 4258 1572
rect 4246 1558 4250 1562
rect 4158 1548 4162 1552
rect 4142 1538 4146 1542
rect 4166 1538 4170 1542
rect 4206 1538 4210 1542
rect 4238 1538 4242 1542
rect 4102 1518 4106 1522
rect 4086 1508 4090 1512
rect 4174 1498 4178 1502
rect 4142 1478 4146 1482
rect 4078 1468 4082 1472
rect 4094 1468 4098 1472
rect 4118 1458 4122 1462
rect 4190 1468 4194 1472
rect 4158 1458 4162 1462
rect 4190 1458 4194 1462
rect 4158 1438 4162 1442
rect 4182 1438 4186 1442
rect 4222 1528 4226 1532
rect 4206 1518 4210 1522
rect 4230 1518 4234 1522
rect 4238 1498 4242 1502
rect 4206 1468 4210 1472
rect 4198 1428 4202 1432
rect 4150 1398 4154 1402
rect 4078 1378 4082 1382
rect 4062 1338 4066 1342
rect 4070 1288 4074 1292
rect 4046 1268 4050 1272
rect 4118 1368 4122 1372
rect 4102 1348 4106 1352
rect 4094 1338 4098 1342
rect 4134 1338 4138 1342
rect 4094 1328 4098 1332
rect 4102 1258 4106 1262
rect 4126 1258 4130 1262
rect 4022 1238 4026 1242
rect 4214 1438 4218 1442
rect 4262 1508 4266 1512
rect 4254 1388 4258 1392
rect 4246 1378 4250 1382
rect 4214 1358 4218 1362
rect 4230 1348 4234 1352
rect 4270 1498 4274 1502
rect 4286 1608 4290 1612
rect 4302 1728 4306 1732
rect 4426 1803 4430 1807
rect 4433 1803 4437 1807
rect 4406 1758 4410 1762
rect 4318 1718 4322 1722
rect 4358 1718 4362 1722
rect 4374 1718 4378 1722
rect 4390 1718 4394 1722
rect 4334 1698 4338 1702
rect 4358 1698 4362 1702
rect 4326 1688 4330 1692
rect 4318 1668 4322 1672
rect 4334 1648 4338 1652
rect 4326 1638 4330 1642
rect 4294 1568 4298 1572
rect 4310 1568 4314 1572
rect 4286 1538 4290 1542
rect 4278 1478 4282 1482
rect 4270 1468 4274 1472
rect 4278 1458 4282 1462
rect 4278 1398 4282 1402
rect 4334 1548 4338 1552
rect 4318 1538 4322 1542
rect 4318 1498 4322 1502
rect 4350 1478 4354 1482
rect 4318 1468 4322 1472
rect 4302 1378 4306 1382
rect 4278 1358 4282 1362
rect 4310 1358 4314 1362
rect 4270 1348 4274 1352
rect 4206 1328 4210 1332
rect 4286 1328 4290 1332
rect 4254 1318 4258 1322
rect 4270 1318 4274 1322
rect 4246 1308 4250 1312
rect 4190 1288 4194 1292
rect 4174 1268 4178 1272
rect 4070 1168 4074 1172
rect 4166 1168 4170 1172
rect 4038 1158 4042 1162
rect 4182 1158 4186 1162
rect 4006 1148 4010 1152
rect 4022 1148 4026 1152
rect 4014 1118 4018 1122
rect 4022 1118 4026 1122
rect 4030 1118 4034 1122
rect 4086 1128 4090 1132
rect 4038 1108 4042 1112
rect 4078 1108 4082 1112
rect 4118 1118 4122 1122
rect 4110 1108 4114 1112
rect 4054 1078 4058 1082
rect 3982 1068 3986 1072
rect 3990 1068 3994 1072
rect 3998 1068 4002 1072
rect 3918 1058 3922 1062
rect 3926 1048 3930 1052
rect 3958 1048 3962 1052
rect 3902 1018 3906 1022
rect 3774 918 3778 922
rect 3822 928 3826 932
rect 3870 928 3874 932
rect 3814 898 3818 902
rect 3766 878 3770 882
rect 3806 878 3810 882
rect 3822 878 3826 882
rect 3678 868 3682 872
rect 3630 858 3634 862
rect 3646 858 3650 862
rect 3662 858 3666 862
rect 3558 808 3562 812
rect 3518 778 3522 782
rect 3542 778 3546 782
rect 3566 778 3570 782
rect 3510 758 3514 762
rect 3502 748 3506 752
rect 3510 738 3514 742
rect 3526 768 3530 772
rect 3494 698 3498 702
rect 3430 688 3434 692
rect 3454 688 3458 692
rect 3558 748 3562 752
rect 3534 738 3538 742
rect 3550 738 3554 742
rect 3526 688 3530 692
rect 3502 678 3506 682
rect 3558 728 3562 732
rect 3614 728 3618 732
rect 3606 718 3610 722
rect 3614 698 3618 702
rect 3550 678 3554 682
rect 3422 668 3426 672
rect 3438 668 3442 672
rect 3502 668 3506 672
rect 3366 638 3370 642
rect 3422 638 3426 642
rect 3402 603 3406 607
rect 3409 603 3413 607
rect 3326 468 3330 472
rect 3342 468 3346 472
rect 3358 468 3362 472
rect 3278 458 3282 462
rect 3262 448 3266 452
rect 3254 388 3258 392
rect 3246 298 3250 302
rect 3294 448 3298 452
rect 3302 348 3306 352
rect 3294 338 3298 342
rect 3302 328 3306 332
rect 3262 288 3266 292
rect 3278 288 3282 292
rect 3294 288 3298 292
rect 3254 268 3258 272
rect 3278 268 3282 272
rect 3254 248 3258 252
rect 3262 238 3266 242
rect 3278 198 3282 202
rect 3262 178 3266 182
rect 3238 138 3242 142
rect 3230 88 3234 92
rect 3230 68 3234 72
rect 3310 298 3314 302
rect 3350 448 3354 452
rect 3326 438 3330 442
rect 3358 438 3362 442
rect 3326 428 3330 432
rect 3326 388 3330 392
rect 3374 518 3378 522
rect 3454 658 3458 662
rect 3534 658 3538 662
rect 3462 648 3466 652
rect 3478 648 3482 652
rect 3446 628 3450 632
rect 3454 568 3458 572
rect 3566 648 3570 652
rect 3510 638 3514 642
rect 3582 628 3586 632
rect 3534 618 3538 622
rect 3518 608 3522 612
rect 3486 558 3490 562
rect 3462 548 3466 552
rect 3494 548 3498 552
rect 3430 538 3434 542
rect 3486 538 3490 542
rect 3526 538 3530 542
rect 3478 518 3482 522
rect 3486 518 3490 522
rect 3502 518 3506 522
rect 3542 488 3546 492
rect 3622 668 3626 672
rect 3670 828 3674 832
rect 3694 808 3698 812
rect 3702 798 3706 802
rect 3814 868 3818 872
rect 3726 858 3730 862
rect 3742 858 3746 862
rect 3798 858 3802 862
rect 3790 848 3794 852
rect 3798 838 3802 842
rect 3806 838 3810 842
rect 4094 1068 4098 1072
rect 4142 1148 4146 1152
rect 4158 1148 4162 1152
rect 4310 1288 4314 1292
rect 4270 1278 4274 1282
rect 4246 1268 4250 1272
rect 4262 1268 4266 1272
rect 4294 1268 4298 1272
rect 4294 1248 4298 1252
rect 4342 1458 4346 1462
rect 4542 2048 4546 2052
rect 4502 1968 4506 1972
rect 4510 1938 4514 1942
rect 4534 1888 4538 1892
rect 4598 2048 4602 2052
rect 4582 2038 4586 2042
rect 4566 1968 4570 1972
rect 4630 2048 4634 2052
rect 4630 1968 4634 1972
rect 4606 1958 4610 1962
rect 4598 1948 4602 1952
rect 4558 1928 4562 1932
rect 4566 1928 4570 1932
rect 4526 1878 4530 1882
rect 4526 1868 4530 1872
rect 4454 1818 4458 1822
rect 4438 1688 4442 1692
rect 4502 1778 4506 1782
rect 4574 1868 4578 1872
rect 4598 1918 4602 1922
rect 4590 1888 4594 1892
rect 4558 1848 4562 1852
rect 4582 1848 4586 1852
rect 4574 1818 4578 1822
rect 4542 1798 4546 1802
rect 4638 1948 4642 1952
rect 4662 2098 4666 2102
rect 4710 2158 4714 2162
rect 4710 2148 4714 2152
rect 4958 2358 4962 2362
rect 5038 2648 5042 2652
rect 5078 2828 5082 2832
rect 5062 2778 5066 2782
rect 5070 2778 5074 2782
rect 5062 2738 5066 2742
rect 5086 2818 5090 2822
rect 5110 2798 5114 2802
rect 5102 2788 5106 2792
rect 5150 3368 5154 3372
rect 5150 3318 5154 3322
rect 5182 3458 5186 3462
rect 5190 3388 5194 3392
rect 5270 3748 5274 3752
rect 5294 3748 5298 3752
rect 5246 3698 5250 3702
rect 5294 3728 5298 3732
rect 5294 3698 5298 3702
rect 5278 3688 5282 3692
rect 5238 3638 5242 3642
rect 5230 3508 5234 3512
rect 5214 3498 5218 3502
rect 5246 3558 5250 3562
rect 5238 3478 5242 3482
rect 5294 3658 5298 3662
rect 5286 3558 5290 3562
rect 5294 3548 5298 3552
rect 5278 3538 5282 3542
rect 5230 3468 5234 3472
rect 5246 3448 5250 3452
rect 5198 3358 5202 3362
rect 5206 3348 5210 3352
rect 5222 3348 5226 3352
rect 5246 3338 5250 3342
rect 5174 3318 5178 3322
rect 5158 3288 5162 3292
rect 5150 3268 5154 3272
rect 5150 3248 5154 3252
rect 5166 3248 5170 3252
rect 5142 3168 5146 3172
rect 5166 3238 5170 3242
rect 5182 3288 5186 3292
rect 5198 3288 5202 3292
rect 5182 3268 5186 3272
rect 5246 3268 5250 3272
rect 5158 3218 5162 3222
rect 5174 3218 5178 3222
rect 5150 3138 5154 3142
rect 5142 3058 5146 3062
rect 5134 2978 5138 2982
rect 5150 2938 5154 2942
rect 5134 2928 5138 2932
rect 5142 2868 5146 2872
rect 5166 3188 5170 3192
rect 5174 3138 5178 3142
rect 5174 3118 5178 3122
rect 5206 3258 5210 3262
rect 5190 3148 5194 3152
rect 5238 3158 5242 3162
rect 5222 3148 5226 3152
rect 5198 3138 5202 3142
rect 5206 3138 5210 3142
rect 5190 3088 5194 3092
rect 5198 3078 5202 3082
rect 5214 3078 5218 3082
rect 5174 3018 5178 3022
rect 5182 2958 5186 2962
rect 5166 2938 5170 2942
rect 5166 2898 5170 2902
rect 5294 3528 5298 3532
rect 5302 3518 5306 3522
rect 5286 3488 5290 3492
rect 5286 3478 5290 3482
rect 5262 3418 5266 3422
rect 5254 3258 5258 3262
rect 5246 3088 5250 3092
rect 5238 3018 5242 3022
rect 5254 3018 5258 3022
rect 5166 2878 5170 2882
rect 5158 2798 5162 2802
rect 5134 2778 5138 2782
rect 5126 2768 5130 2772
rect 5086 2758 5090 2762
rect 5230 2898 5234 2902
rect 5214 2848 5218 2852
rect 5230 2848 5234 2852
rect 5214 2838 5218 2842
rect 5222 2818 5226 2822
rect 5198 2748 5202 2752
rect 5214 2748 5218 2752
rect 5126 2738 5130 2742
rect 5198 2738 5202 2742
rect 5086 2728 5090 2732
rect 5078 2678 5082 2682
rect 5086 2658 5090 2662
rect 5142 2658 5146 2662
rect 5046 2548 5050 2552
rect 5030 2528 5034 2532
rect 5046 2528 5050 2532
rect 5070 2498 5074 2502
rect 5006 2488 5010 2492
rect 5102 2618 5106 2622
rect 5094 2568 5098 2572
rect 5094 2538 5098 2542
rect 5270 3338 5274 3342
rect 5286 3338 5290 3342
rect 5294 3338 5298 3342
rect 5270 3248 5274 3252
rect 5294 3118 5298 3122
rect 5286 3018 5290 3022
rect 5278 3008 5282 3012
rect 5270 2948 5274 2952
rect 5286 2938 5290 2942
rect 5294 2928 5298 2932
rect 5254 2918 5258 2922
rect 5246 2828 5250 2832
rect 5238 2788 5242 2792
rect 5238 2748 5242 2752
rect 5238 2718 5242 2722
rect 5286 2828 5290 2832
rect 5254 2788 5258 2792
rect 5254 2738 5258 2742
rect 5238 2648 5242 2652
rect 5198 2608 5202 2612
rect 5158 2588 5162 2592
rect 5158 2568 5162 2572
rect 5126 2558 5130 2562
rect 5142 2548 5146 2552
rect 5094 2498 5098 2502
rect 5118 2498 5122 2502
rect 5038 2478 5042 2482
rect 5078 2478 5082 2482
rect 5054 2438 5058 2442
rect 5062 2378 5066 2382
rect 5014 2358 5018 2362
rect 4982 2348 4986 2352
rect 4926 2318 4930 2322
rect 4918 2298 4922 2302
rect 4798 2268 4802 2272
rect 4806 2268 4810 2272
rect 4838 2268 4842 2272
rect 4910 2268 4914 2272
rect 4846 2258 4850 2262
rect 4774 2178 4778 2182
rect 4782 2178 4786 2182
rect 4822 2158 4826 2162
rect 4854 2218 4858 2222
rect 4854 2208 4858 2212
rect 4938 2303 4942 2307
rect 4945 2303 4949 2307
rect 4966 2338 4970 2342
rect 4998 2338 5002 2342
rect 4990 2328 4994 2332
rect 5046 2328 5050 2332
rect 5030 2318 5034 2322
rect 5022 2288 5026 2292
rect 4982 2278 4986 2282
rect 5006 2248 5010 2252
rect 4958 2198 4962 2202
rect 4942 2168 4946 2172
rect 4910 2158 4914 2162
rect 4774 2148 4778 2152
rect 4830 2148 4834 2152
rect 4846 2148 4850 2152
rect 4878 2148 4882 2152
rect 4910 2148 4914 2152
rect 4726 2138 4730 2142
rect 4918 2138 4922 2142
rect 4750 2128 4754 2132
rect 4726 2108 4730 2112
rect 4734 2078 4738 2082
rect 4654 2068 4658 2072
rect 4742 2068 4746 2072
rect 4662 2058 4666 2062
rect 4678 2058 4682 2062
rect 4798 2058 4802 2062
rect 4830 2058 4834 2062
rect 4750 2048 4754 2052
rect 4654 2038 4658 2042
rect 4710 2038 4714 2042
rect 4654 2028 4658 2032
rect 4614 1908 4618 1912
rect 4638 1908 4642 1912
rect 4630 1898 4634 1902
rect 4638 1868 4642 1872
rect 4782 1978 4786 1982
rect 4830 1978 4834 1982
rect 4862 2088 4866 2092
rect 4886 2068 4890 2072
rect 4870 2018 4874 2022
rect 4862 2008 4866 2012
rect 4854 1968 4858 1972
rect 4790 1958 4794 1962
rect 4822 1958 4826 1962
rect 4766 1938 4770 1942
rect 4838 1938 4842 1942
rect 4854 1938 4858 1942
rect 4750 1928 4754 1932
rect 4790 1908 4794 1912
rect 4758 1888 4762 1892
rect 4806 1888 4810 1892
rect 4846 1888 4850 1892
rect 4814 1878 4818 1882
rect 4686 1868 4690 1872
rect 4750 1868 4754 1872
rect 4614 1848 4618 1852
rect 4646 1858 4650 1862
rect 4758 1858 4762 1862
rect 4790 1858 4794 1862
rect 4846 1858 4850 1862
rect 4870 1968 4874 1972
rect 4878 1898 4882 1902
rect 4878 1858 4882 1862
rect 4654 1838 4658 1842
rect 4694 1838 4698 1842
rect 4630 1818 4634 1822
rect 4678 1818 4682 1822
rect 4622 1808 4626 1812
rect 4510 1768 4514 1772
rect 4574 1768 4578 1772
rect 4510 1758 4514 1762
rect 4542 1758 4546 1762
rect 4614 1758 4618 1762
rect 4550 1748 4554 1752
rect 4606 1748 4610 1752
rect 4462 1728 4466 1732
rect 4462 1698 4466 1702
rect 4518 1698 4522 1702
rect 4426 1603 4430 1607
rect 4433 1603 4437 1607
rect 4470 1668 4474 1672
rect 4486 1668 4490 1672
rect 4478 1658 4482 1662
rect 4502 1658 4506 1662
rect 4518 1658 4522 1662
rect 4582 1658 4586 1662
rect 4462 1588 4466 1592
rect 4454 1578 4458 1582
rect 4398 1568 4402 1572
rect 4438 1568 4442 1572
rect 4382 1538 4386 1542
rect 4366 1508 4370 1512
rect 4382 1498 4386 1502
rect 4390 1478 4394 1482
rect 4406 1538 4410 1542
rect 4438 1538 4442 1542
rect 4406 1478 4410 1482
rect 4398 1468 4402 1472
rect 4462 1518 4466 1522
rect 4470 1508 4474 1512
rect 4502 1618 4506 1622
rect 4494 1578 4498 1582
rect 4590 1648 4594 1652
rect 4582 1588 4586 1592
rect 4534 1558 4538 1562
rect 4542 1558 4546 1562
rect 4566 1558 4570 1562
rect 4494 1508 4498 1512
rect 4462 1468 4466 1472
rect 4478 1468 4482 1472
rect 4486 1468 4490 1472
rect 4454 1458 4458 1462
rect 4326 1408 4330 1412
rect 4398 1448 4402 1452
rect 4430 1418 4434 1422
rect 4382 1408 4386 1412
rect 4426 1403 4430 1407
rect 4433 1403 4437 1407
rect 4374 1398 4378 1402
rect 4438 1378 4442 1382
rect 4390 1358 4394 1362
rect 4422 1358 4426 1362
rect 4374 1348 4378 1352
rect 4326 1318 4330 1322
rect 4398 1298 4402 1302
rect 4326 1288 4330 1292
rect 4350 1278 4354 1282
rect 4374 1278 4378 1282
rect 4326 1268 4330 1272
rect 4342 1268 4346 1272
rect 4454 1338 4458 1342
rect 4486 1458 4490 1462
rect 4494 1388 4498 1392
rect 4478 1358 4482 1362
rect 4502 1378 4506 1382
rect 4502 1368 4506 1372
rect 4494 1338 4498 1342
rect 4478 1318 4482 1322
rect 4470 1288 4474 1292
rect 4566 1548 4570 1552
rect 4558 1508 4562 1512
rect 4574 1498 4578 1502
rect 4590 1558 4594 1562
rect 4598 1558 4602 1562
rect 4702 1758 4706 1762
rect 4670 1748 4674 1752
rect 4686 1748 4690 1752
rect 4702 1748 4706 1752
rect 4638 1738 4642 1742
rect 4742 1828 4746 1832
rect 4758 1828 4762 1832
rect 4766 1828 4770 1832
rect 4726 1768 4730 1772
rect 4718 1758 4722 1762
rect 4734 1758 4738 1762
rect 4654 1728 4658 1732
rect 4710 1728 4714 1732
rect 4734 1728 4738 1732
rect 4662 1688 4666 1692
rect 4718 1688 4722 1692
rect 4678 1668 4682 1672
rect 4718 1668 4722 1672
rect 4694 1658 4698 1662
rect 4710 1658 4714 1662
rect 4646 1628 4650 1632
rect 4702 1598 4706 1602
rect 4670 1578 4674 1582
rect 4702 1578 4706 1582
rect 4662 1568 4666 1572
rect 4630 1558 4634 1562
rect 4646 1558 4650 1562
rect 4606 1508 4610 1512
rect 4590 1488 4594 1492
rect 4550 1448 4554 1452
rect 4574 1418 4578 1422
rect 4518 1368 4522 1372
rect 4598 1368 4602 1372
rect 4518 1358 4522 1362
rect 4582 1358 4586 1362
rect 4542 1338 4546 1342
rect 4510 1278 4514 1282
rect 4390 1268 4394 1272
rect 4406 1268 4410 1272
rect 4510 1268 4514 1272
rect 4334 1258 4338 1262
rect 4366 1258 4370 1262
rect 4398 1258 4402 1262
rect 4334 1248 4338 1252
rect 4382 1248 4386 1252
rect 4446 1248 4450 1252
rect 4286 1208 4290 1212
rect 4214 1188 4218 1192
rect 4190 1118 4194 1122
rect 4174 1108 4178 1112
rect 4126 1088 4130 1092
rect 4014 1058 4018 1062
rect 4046 1058 4050 1062
rect 4110 1058 4114 1062
rect 4054 1018 4058 1022
rect 3974 988 3978 992
rect 3918 928 3922 932
rect 3950 918 3954 922
rect 3902 908 3906 912
rect 3854 858 3858 862
rect 3838 848 3842 852
rect 3814 788 3818 792
rect 3846 788 3850 792
rect 3678 758 3682 762
rect 3694 758 3698 762
rect 3646 698 3650 702
rect 3670 688 3674 692
rect 3686 688 3690 692
rect 3686 658 3690 662
rect 3670 648 3674 652
rect 3686 648 3690 652
rect 3662 638 3666 642
rect 3678 638 3682 642
rect 3558 578 3562 582
rect 3566 568 3570 572
rect 3606 568 3610 572
rect 3582 548 3586 552
rect 3590 538 3594 542
rect 3550 478 3554 482
rect 3598 528 3602 532
rect 3686 558 3690 562
rect 3870 838 3874 842
rect 3922 903 3926 907
rect 3929 903 3933 907
rect 3950 888 3954 892
rect 3958 888 3962 892
rect 3886 838 3890 842
rect 3878 808 3882 812
rect 3862 768 3866 772
rect 3710 748 3714 752
rect 3798 748 3802 752
rect 3766 738 3770 742
rect 3806 738 3810 742
rect 3814 738 3818 742
rect 3886 788 3890 792
rect 3878 738 3882 742
rect 3814 728 3818 732
rect 3862 728 3866 732
rect 3734 718 3738 722
rect 3782 698 3786 702
rect 3718 678 3722 682
rect 3766 668 3770 672
rect 3710 658 3714 662
rect 3758 648 3762 652
rect 3646 548 3650 552
rect 3654 538 3658 542
rect 3670 538 3674 542
rect 3606 508 3610 512
rect 3590 498 3594 502
rect 3534 468 3538 472
rect 3558 468 3562 472
rect 3382 458 3386 462
rect 3470 458 3474 462
rect 3526 458 3530 462
rect 3550 458 3554 462
rect 3382 448 3386 452
rect 3470 418 3474 422
rect 3402 403 3406 407
rect 3409 403 3413 407
rect 3390 388 3394 392
rect 3382 348 3386 352
rect 3566 448 3570 452
rect 3582 448 3586 452
rect 3606 448 3610 452
rect 3526 438 3530 442
rect 3598 438 3602 442
rect 3534 418 3538 422
rect 3534 408 3538 412
rect 3486 398 3490 402
rect 3598 388 3602 392
rect 3558 378 3562 382
rect 3654 458 3658 462
rect 3662 418 3666 422
rect 3662 398 3666 402
rect 3726 528 3730 532
rect 3718 498 3722 502
rect 3870 698 3874 702
rect 3870 678 3874 682
rect 3966 878 3970 882
rect 3990 928 3994 932
rect 4014 928 4018 932
rect 4006 888 4010 892
rect 4014 878 4018 882
rect 3974 868 3978 872
rect 3918 858 3922 862
rect 3974 858 3978 862
rect 3942 848 3946 852
rect 3950 768 3954 772
rect 3918 758 3922 762
rect 3966 758 3970 762
rect 3974 748 3978 752
rect 3934 738 3938 742
rect 3958 738 3962 742
rect 3974 738 3978 742
rect 4014 798 4018 802
rect 3998 758 4002 762
rect 4038 788 4042 792
rect 4174 1068 4178 1072
rect 4166 1058 4170 1062
rect 4198 1058 4202 1062
rect 4422 1238 4426 1242
rect 4414 1208 4418 1212
rect 4326 1178 4330 1182
rect 4246 1168 4250 1172
rect 4382 1168 4386 1172
rect 4406 1168 4410 1172
rect 4358 1158 4362 1162
rect 4366 1148 4370 1152
rect 4390 1148 4394 1152
rect 4294 1138 4298 1142
rect 4326 1138 4330 1142
rect 4254 1128 4258 1132
rect 4350 1128 4354 1132
rect 4278 1118 4282 1122
rect 4398 1138 4402 1142
rect 4350 1118 4354 1122
rect 4358 1118 4362 1122
rect 4426 1203 4430 1207
rect 4433 1203 4437 1207
rect 4462 1178 4466 1182
rect 4574 1318 4578 1322
rect 4542 1298 4546 1302
rect 4574 1278 4578 1282
rect 4590 1348 4594 1352
rect 4622 1508 4626 1512
rect 4630 1508 4634 1512
rect 4614 1498 4618 1502
rect 4686 1568 4690 1572
rect 4702 1558 4706 1562
rect 4870 1848 4874 1852
rect 4878 1778 4882 1782
rect 4862 1758 4866 1762
rect 4830 1748 4834 1752
rect 4846 1748 4850 1752
rect 4862 1748 4866 1752
rect 4938 2103 4942 2107
rect 4945 2103 4949 2107
rect 5046 2268 5050 2272
rect 5030 2198 5034 2202
rect 4998 2178 5002 2182
rect 5022 2158 5026 2162
rect 5030 2158 5034 2162
rect 4966 2148 4970 2152
rect 4926 1998 4930 2002
rect 4894 1918 4898 1922
rect 4798 1738 4802 1742
rect 4846 1738 4850 1742
rect 4814 1728 4818 1732
rect 4886 1728 4890 1732
rect 4926 1918 4930 1922
rect 4918 1908 4922 1912
rect 4938 1903 4942 1907
rect 4945 1903 4949 1907
rect 4926 1888 4930 1892
rect 4958 1878 4962 1882
rect 4902 1718 4906 1722
rect 4750 1698 4754 1702
rect 4742 1658 4746 1662
rect 4654 1468 4658 1472
rect 4622 1458 4626 1462
rect 4638 1398 4642 1402
rect 4614 1358 4618 1362
rect 4694 1458 4698 1462
rect 4894 1688 4898 1692
rect 4774 1678 4778 1682
rect 4790 1668 4794 1672
rect 5054 2138 5058 2142
rect 4998 2128 5002 2132
rect 5046 2088 5050 2092
rect 5014 2068 5018 2072
rect 4998 2058 5002 2062
rect 5046 2058 5050 2062
rect 4974 2028 4978 2032
rect 5030 2028 5034 2032
rect 4990 2018 4994 2022
rect 5014 1948 5018 1952
rect 4998 1928 5002 1932
rect 4982 1908 4986 1912
rect 4982 1878 4986 1882
rect 4942 1738 4946 1742
rect 4938 1703 4942 1707
rect 4945 1703 4949 1707
rect 4918 1668 4922 1672
rect 4774 1658 4778 1662
rect 4862 1658 4866 1662
rect 4886 1658 4890 1662
rect 4758 1648 4762 1652
rect 4822 1648 4826 1652
rect 4862 1638 4866 1642
rect 4830 1558 4834 1562
rect 4838 1558 4842 1562
rect 4982 1838 4986 1842
rect 5014 1888 5018 1892
rect 5006 1878 5010 1882
rect 5046 1948 5050 1952
rect 5038 1938 5042 1942
rect 5046 1918 5050 1922
rect 5022 1868 5026 1872
rect 5014 1858 5018 1862
rect 5030 1858 5034 1862
rect 5046 1858 5050 1862
rect 5014 1808 5018 1812
rect 5158 2518 5162 2522
rect 5190 2498 5194 2502
rect 5214 2548 5218 2552
rect 5198 2488 5202 2492
rect 5286 2808 5290 2812
rect 5278 2748 5282 2752
rect 5262 2558 5266 2562
rect 5246 2538 5250 2542
rect 5254 2518 5258 2522
rect 5150 2468 5154 2472
rect 5206 2458 5210 2462
rect 5078 2448 5082 2452
rect 5126 2448 5130 2452
rect 5150 2438 5154 2442
rect 5078 2388 5082 2392
rect 5126 2388 5130 2392
rect 5134 2388 5138 2392
rect 5070 2248 5074 2252
rect 5070 2218 5074 2222
rect 5110 2358 5114 2362
rect 5246 2358 5250 2362
rect 5278 2518 5282 2522
rect 5262 2388 5266 2392
rect 5294 2408 5298 2412
rect 5270 2368 5274 2372
rect 5278 2358 5282 2362
rect 5302 2378 5306 2382
rect 5174 2348 5178 2352
rect 5086 2298 5090 2302
rect 5078 2208 5082 2212
rect 5078 2188 5082 2192
rect 5078 2168 5082 2172
rect 5150 2288 5154 2292
rect 5158 2288 5162 2292
rect 5214 2328 5218 2332
rect 5238 2338 5242 2342
rect 5214 2308 5218 2312
rect 5222 2308 5226 2312
rect 5254 2308 5258 2312
rect 5102 2278 5106 2282
rect 5174 2278 5178 2282
rect 5142 2268 5146 2272
rect 5198 2268 5202 2272
rect 5102 2258 5106 2262
rect 5150 2258 5154 2262
rect 5150 2248 5154 2252
rect 5142 2218 5146 2222
rect 5086 2158 5090 2162
rect 5134 2158 5138 2162
rect 5158 2238 5162 2242
rect 5182 2218 5186 2222
rect 5198 2198 5202 2202
rect 5182 2178 5186 2182
rect 5174 2158 5178 2162
rect 5110 2148 5114 2152
rect 5142 2148 5146 2152
rect 5166 2148 5170 2152
rect 5126 2138 5130 2142
rect 5150 2138 5154 2142
rect 5070 2078 5074 2082
rect 5118 2128 5122 2132
rect 5110 2118 5114 2122
rect 5102 2108 5106 2112
rect 5126 2088 5130 2092
rect 5086 2068 5090 2072
rect 5110 2058 5114 2062
rect 5086 2038 5090 2042
rect 5102 2028 5106 2032
rect 5062 1958 5066 1962
rect 5158 2078 5162 2082
rect 5062 1908 5066 1912
rect 5094 1868 5098 1872
rect 5126 1938 5130 1942
rect 5150 1928 5154 1932
rect 5190 2138 5194 2142
rect 5262 2288 5266 2292
rect 5270 2258 5274 2262
rect 5302 2258 5306 2262
rect 5238 2228 5242 2232
rect 5222 2098 5226 2102
rect 5198 2078 5202 2082
rect 5230 2078 5234 2082
rect 5222 2068 5226 2072
rect 5270 2218 5274 2222
rect 5262 2198 5266 2202
rect 5254 2168 5258 2172
rect 5254 2088 5258 2092
rect 5286 2178 5290 2182
rect 5270 2068 5274 2072
rect 5286 2058 5290 2062
rect 5246 2018 5250 2022
rect 5262 1958 5266 1962
rect 5230 1948 5234 1952
rect 5214 1938 5218 1942
rect 5126 1918 5130 1922
rect 5134 1918 5138 1922
rect 5150 1918 5154 1922
rect 5182 1918 5186 1922
rect 5142 1878 5146 1882
rect 5110 1858 5114 1862
rect 5046 1778 5050 1782
rect 4982 1768 4986 1772
rect 4998 1768 5002 1772
rect 4966 1758 4970 1762
rect 4974 1708 4978 1712
rect 4966 1678 4970 1682
rect 4958 1618 4962 1622
rect 4902 1598 4906 1602
rect 4878 1568 4882 1572
rect 4886 1568 4890 1572
rect 4758 1547 4762 1551
rect 4822 1548 4826 1552
rect 4854 1548 4858 1552
rect 4878 1548 4882 1552
rect 4894 1548 4898 1552
rect 4806 1538 4810 1542
rect 4814 1538 4818 1542
rect 4846 1538 4850 1542
rect 4798 1528 4802 1532
rect 4886 1538 4890 1542
rect 4758 1488 4762 1492
rect 4790 1488 4794 1492
rect 4838 1488 4842 1492
rect 4766 1478 4770 1482
rect 4670 1418 4674 1422
rect 4742 1418 4746 1422
rect 4702 1408 4706 1412
rect 4686 1378 4690 1382
rect 4814 1478 4818 1482
rect 4862 1518 4866 1522
rect 4806 1468 4810 1472
rect 4822 1468 4826 1472
rect 4782 1458 4786 1462
rect 4814 1458 4818 1462
rect 4846 1448 4850 1452
rect 4798 1428 4802 1432
rect 4790 1418 4794 1422
rect 4774 1378 4778 1382
rect 4830 1378 4834 1382
rect 4718 1358 4722 1362
rect 4806 1358 4810 1362
rect 4630 1348 4634 1352
rect 4678 1348 4682 1352
rect 4766 1348 4770 1352
rect 4622 1338 4626 1342
rect 4654 1338 4658 1342
rect 4670 1338 4674 1342
rect 4622 1288 4626 1292
rect 4542 1248 4546 1252
rect 4550 1148 4554 1152
rect 4470 1138 4474 1142
rect 4414 1118 4418 1122
rect 4398 1098 4402 1102
rect 4238 1088 4242 1092
rect 4254 1088 4258 1092
rect 4286 1088 4290 1092
rect 4326 1088 4330 1092
rect 4350 1088 4354 1092
rect 4238 1068 4242 1072
rect 4238 1058 4242 1062
rect 4150 1048 4154 1052
rect 4166 1048 4170 1052
rect 4174 1048 4178 1052
rect 4142 1038 4146 1042
rect 4110 1018 4114 1022
rect 4102 1008 4106 1012
rect 4190 998 4194 1002
rect 4142 988 4146 992
rect 4198 988 4202 992
rect 4134 978 4138 982
rect 4070 948 4074 952
rect 4070 938 4074 942
rect 4094 918 4098 922
rect 4134 938 4138 942
rect 4086 898 4090 902
rect 4110 898 4114 902
rect 4094 888 4098 892
rect 4102 878 4106 882
rect 4062 868 4066 872
rect 4078 838 4082 842
rect 4054 778 4058 782
rect 4086 778 4090 782
rect 4062 768 4066 772
rect 4006 748 4010 752
rect 3990 738 3994 742
rect 3982 728 3986 732
rect 3922 703 3926 707
rect 3929 703 3933 707
rect 3982 688 3986 692
rect 3926 678 3930 682
rect 3990 678 3994 682
rect 3838 668 3842 672
rect 3862 668 3866 672
rect 3910 668 3914 672
rect 4046 758 4050 762
rect 4078 758 4082 762
rect 4118 868 4122 872
rect 4198 968 4202 972
rect 4206 968 4210 972
rect 4206 948 4210 952
rect 4222 948 4226 952
rect 4174 938 4178 942
rect 4190 938 4194 942
rect 4222 928 4226 932
rect 4222 908 4226 912
rect 4150 898 4154 902
rect 4182 898 4186 902
rect 4214 898 4218 902
rect 4150 868 4154 872
rect 4134 768 4138 772
rect 4110 758 4114 762
rect 4030 748 4034 752
rect 4062 728 4066 732
rect 4094 728 4098 732
rect 4086 718 4090 722
rect 4062 698 4066 702
rect 4038 678 4042 682
rect 4030 668 4034 672
rect 3870 658 3874 662
rect 3846 648 3850 652
rect 3806 628 3810 632
rect 3790 578 3794 582
rect 3790 518 3794 522
rect 3782 508 3786 512
rect 3862 578 3866 582
rect 3958 648 3962 652
rect 3886 588 3890 592
rect 3878 578 3882 582
rect 3918 568 3922 572
rect 3830 548 3834 552
rect 3894 548 3898 552
rect 3822 528 3826 532
rect 3990 658 3994 662
rect 4006 658 4010 662
rect 4022 658 4026 662
rect 3998 588 4002 592
rect 4030 578 4034 582
rect 4006 568 4010 572
rect 3950 558 3954 562
rect 3974 558 3978 562
rect 3958 548 3962 552
rect 3982 548 3986 552
rect 3990 548 3994 552
rect 4022 548 4026 552
rect 3886 538 3890 542
rect 3958 538 3962 542
rect 3942 528 3946 532
rect 3950 528 3954 532
rect 3878 518 3882 522
rect 3854 508 3858 512
rect 3922 503 3926 507
rect 3929 503 3933 507
rect 3998 538 4002 542
rect 4030 538 4034 542
rect 4022 528 4026 532
rect 3982 518 3986 522
rect 3878 498 3882 502
rect 3974 498 3978 502
rect 4006 498 4010 502
rect 3718 468 3722 472
rect 3862 468 3866 472
rect 3702 448 3706 452
rect 3710 438 3714 442
rect 3694 428 3698 432
rect 3686 398 3690 402
rect 3622 358 3626 362
rect 3542 348 3546 352
rect 3574 348 3578 352
rect 3582 348 3586 352
rect 3366 338 3370 342
rect 3646 338 3650 342
rect 3390 328 3394 332
rect 3318 278 3322 282
rect 3342 278 3346 282
rect 3382 268 3386 272
rect 3342 258 3346 262
rect 3374 248 3378 252
rect 3334 238 3338 242
rect 3470 318 3474 322
rect 3438 298 3442 302
rect 3478 278 3482 282
rect 3518 278 3522 282
rect 3534 268 3538 272
rect 3478 258 3482 262
rect 3502 258 3506 262
rect 3454 228 3458 232
rect 3402 203 3406 207
rect 3409 203 3413 207
rect 3390 198 3394 202
rect 3318 168 3322 172
rect 3422 168 3426 172
rect 3334 158 3338 162
rect 3430 148 3434 152
rect 3414 138 3418 142
rect 3358 98 3362 102
rect 3310 78 3314 82
rect 3318 68 3322 72
rect 3462 188 3466 192
rect 3550 218 3554 222
rect 3478 168 3482 172
rect 3470 158 3474 162
rect 3574 328 3578 332
rect 3646 328 3650 332
rect 3614 318 3618 322
rect 3598 298 3602 302
rect 3622 298 3626 302
rect 3710 408 3714 412
rect 3742 458 3746 462
rect 3742 448 3746 452
rect 3758 428 3762 432
rect 3734 388 3738 392
rect 3718 378 3722 382
rect 3774 448 3778 452
rect 3830 458 3834 462
rect 3822 448 3826 452
rect 3798 398 3802 402
rect 3790 378 3794 382
rect 3734 368 3738 372
rect 3758 368 3762 372
rect 3766 368 3770 372
rect 3726 358 3730 362
rect 3662 348 3666 352
rect 3702 348 3706 352
rect 3686 328 3690 332
rect 3678 318 3682 322
rect 3678 298 3682 302
rect 3670 278 3674 282
rect 3670 238 3674 242
rect 3654 228 3658 232
rect 3646 218 3650 222
rect 3622 208 3626 212
rect 3654 198 3658 202
rect 3710 338 3714 342
rect 3710 288 3714 292
rect 3694 248 3698 252
rect 3702 238 3706 242
rect 3694 188 3698 192
rect 3582 168 3586 172
rect 3678 168 3682 172
rect 3606 158 3610 162
rect 3654 158 3658 162
rect 3726 218 3730 222
rect 3742 358 3746 362
rect 3750 348 3754 352
rect 3766 348 3770 352
rect 3766 338 3770 342
rect 3742 328 3746 332
rect 3782 328 3786 332
rect 3750 318 3754 322
rect 3758 298 3762 302
rect 3790 278 3794 282
rect 3990 478 3994 482
rect 4030 478 4034 482
rect 3894 468 3898 472
rect 3934 468 3938 472
rect 3974 468 3978 472
rect 4014 458 4018 462
rect 3926 448 3930 452
rect 3870 408 3874 412
rect 3814 358 3818 362
rect 3838 358 3842 362
rect 3830 338 3834 342
rect 3846 338 3850 342
rect 3822 328 3826 332
rect 3830 328 3834 332
rect 3822 308 3826 312
rect 3830 278 3834 282
rect 3798 268 3802 272
rect 3838 268 3842 272
rect 3806 258 3810 262
rect 3790 248 3794 252
rect 3750 238 3754 242
rect 3782 238 3786 242
rect 3814 238 3818 242
rect 3862 298 3866 302
rect 3854 288 3858 292
rect 3750 188 3754 192
rect 3766 188 3770 192
rect 3862 218 3866 222
rect 3734 178 3738 182
rect 3462 148 3466 152
rect 3486 148 3490 152
rect 3518 148 3522 152
rect 3526 148 3530 152
rect 3646 148 3650 152
rect 3838 168 3842 172
rect 3822 158 3826 162
rect 3526 128 3530 132
rect 3454 108 3458 112
rect 3438 88 3442 92
rect 3462 88 3466 92
rect 3486 88 3490 92
rect 3606 138 3610 142
rect 3622 138 3626 142
rect 3654 138 3658 142
rect 3686 138 3690 142
rect 3702 138 3706 142
rect 3630 128 3634 132
rect 3686 128 3690 132
rect 3566 118 3570 122
rect 3710 108 3714 112
rect 3534 98 3538 102
rect 3590 98 3594 102
rect 3606 98 3610 102
rect 3542 88 3546 92
rect 3494 78 3498 82
rect 3430 68 3434 72
rect 3942 448 3946 452
rect 3982 428 3986 432
rect 4022 428 4026 432
rect 3934 398 3938 402
rect 3886 368 3890 372
rect 3926 348 3930 352
rect 4022 418 4026 422
rect 3982 358 3986 362
rect 3886 338 3890 342
rect 3878 318 3882 322
rect 4062 668 4066 672
rect 4118 728 4122 732
rect 4102 718 4106 722
rect 4102 708 4106 712
rect 4086 678 4090 682
rect 4110 668 4114 672
rect 4142 758 4146 762
rect 4142 748 4146 752
rect 4206 868 4210 872
rect 4246 1028 4250 1032
rect 4254 978 4258 982
rect 4526 1118 4530 1122
rect 4462 1088 4466 1092
rect 4486 1088 4490 1092
rect 4302 1068 4306 1072
rect 4366 1058 4370 1062
rect 4382 1058 4386 1062
rect 4558 1138 4562 1142
rect 4566 1138 4570 1142
rect 4542 1068 4546 1072
rect 4414 1058 4418 1062
rect 4334 1048 4338 1052
rect 4390 1048 4394 1052
rect 4406 1048 4410 1052
rect 4390 1028 4394 1032
rect 4286 968 4290 972
rect 4270 958 4274 962
rect 4262 938 4266 942
rect 4526 1048 4530 1052
rect 4494 1008 4498 1012
rect 4526 1008 4530 1012
rect 4426 1003 4430 1007
rect 4433 1003 4437 1007
rect 4430 988 4434 992
rect 4486 988 4490 992
rect 4302 928 4306 932
rect 4278 908 4282 912
rect 4374 928 4378 932
rect 4374 918 4378 922
rect 4286 878 4290 882
rect 4358 868 4362 872
rect 4366 868 4370 872
rect 4406 928 4410 932
rect 4214 858 4218 862
rect 4198 848 4202 852
rect 4174 828 4178 832
rect 4182 828 4186 832
rect 4198 828 4202 832
rect 4158 808 4162 812
rect 4166 808 4170 812
rect 4166 778 4170 782
rect 4158 758 4162 762
rect 4182 728 4186 732
rect 4190 728 4194 732
rect 4150 708 4154 712
rect 4142 698 4146 702
rect 4238 848 4242 852
rect 4230 838 4234 842
rect 4222 708 4226 712
rect 4190 688 4194 692
rect 4198 678 4202 682
rect 4262 848 4266 852
rect 4286 838 4290 842
rect 4254 828 4258 832
rect 4310 858 4314 862
rect 4342 858 4346 862
rect 4294 758 4298 762
rect 4302 758 4306 762
rect 4342 748 4346 752
rect 4278 728 4282 732
rect 4334 728 4338 732
rect 4302 668 4306 672
rect 4078 658 4082 662
rect 4126 658 4130 662
rect 4198 658 4202 662
rect 4294 658 4298 662
rect 4070 648 4074 652
rect 4086 618 4090 622
rect 4046 498 4050 502
rect 4038 408 4042 412
rect 4038 388 4042 392
rect 4046 378 4050 382
rect 4054 378 4058 382
rect 4030 368 4034 372
rect 4046 368 4050 372
rect 3894 328 3898 332
rect 3886 308 3890 312
rect 3878 258 3882 262
rect 3870 148 3874 152
rect 3870 138 3874 142
rect 3870 98 3874 102
rect 3622 88 3626 92
rect 3710 88 3714 92
rect 3774 88 3778 92
rect 3854 88 3858 92
rect 3862 88 3866 92
rect 3582 78 3586 82
rect 3606 78 3610 82
rect 3686 78 3690 82
rect 3838 78 3842 82
rect 3214 58 3218 62
rect 3254 58 3258 62
rect 3310 58 3314 62
rect 3622 68 3626 72
rect 3558 58 3562 62
rect 3582 58 3586 62
rect 3598 58 3602 62
rect 3742 68 3746 72
rect 3758 68 3762 72
rect 3734 58 3738 62
rect 3922 303 3926 307
rect 3929 303 3933 307
rect 4022 328 4026 332
rect 4022 288 4026 292
rect 3910 278 3914 282
rect 4078 358 4082 362
rect 4054 288 4058 292
rect 3958 258 3962 262
rect 4014 258 4018 262
rect 4046 258 4050 262
rect 4038 248 4042 252
rect 4054 238 4058 242
rect 3902 218 3906 222
rect 3902 208 3906 212
rect 4046 228 4050 232
rect 4078 198 4082 202
rect 4054 178 4058 182
rect 3998 168 4002 172
rect 3926 158 3930 162
rect 4062 158 4066 162
rect 3918 148 3922 152
rect 3918 138 3922 142
rect 3974 138 3978 142
rect 4030 138 4034 142
rect 4054 138 4058 142
rect 4078 138 4082 142
rect 3886 128 3890 132
rect 3950 128 3954 132
rect 3922 103 3926 107
rect 3929 103 3933 107
rect 3942 98 3946 102
rect 3902 88 3906 92
rect 4038 118 4042 122
rect 4014 88 4018 92
rect 3966 78 3970 82
rect 3894 68 3898 72
rect 3910 68 3914 72
rect 4030 78 4034 82
rect 3886 58 3890 62
rect 4054 88 4058 92
rect 4174 648 4178 652
rect 4302 648 4306 652
rect 4318 648 4322 652
rect 4198 618 4202 622
rect 4134 598 4138 602
rect 4110 588 4114 592
rect 4318 638 4322 642
rect 4342 618 4346 622
rect 4150 568 4154 572
rect 4198 568 4202 572
rect 4214 568 4218 572
rect 4134 558 4138 562
rect 4222 558 4226 562
rect 4454 968 4458 972
rect 4446 958 4450 962
rect 4478 948 4482 952
rect 4470 938 4474 942
rect 4494 938 4498 942
rect 4510 938 4514 942
rect 4502 928 4506 932
rect 4510 918 4514 922
rect 4542 918 4546 922
rect 4446 908 4450 912
rect 4406 858 4410 862
rect 4430 848 4434 852
rect 4390 838 4394 842
rect 4390 808 4394 812
rect 4426 803 4430 807
rect 4433 803 4437 807
rect 4382 778 4386 782
rect 4414 778 4418 782
rect 4430 778 4434 782
rect 4422 758 4426 762
rect 4454 878 4458 882
rect 4606 1258 4610 1262
rect 4590 1248 4594 1252
rect 4654 1238 4658 1242
rect 4646 1198 4650 1202
rect 4662 1208 4666 1212
rect 4630 1188 4634 1192
rect 4638 1188 4642 1192
rect 4670 1188 4674 1192
rect 4662 1178 4666 1182
rect 4670 1168 4674 1172
rect 4702 1338 4706 1342
rect 4734 1338 4738 1342
rect 4758 1338 4762 1342
rect 4742 1328 4746 1332
rect 4774 1308 4778 1312
rect 4766 1288 4770 1292
rect 4694 1268 4698 1272
rect 4718 1258 4722 1262
rect 4686 1218 4690 1222
rect 4678 1158 4682 1162
rect 4590 1148 4594 1152
rect 4622 1148 4626 1152
rect 4678 1148 4682 1152
rect 4582 1138 4586 1142
rect 4598 1138 4602 1142
rect 4582 1128 4586 1132
rect 4590 1088 4594 1092
rect 4574 1078 4578 1082
rect 4566 1058 4570 1062
rect 4582 1048 4586 1052
rect 4558 998 4562 1002
rect 4558 918 4562 922
rect 4502 888 4506 892
rect 4526 888 4530 892
rect 4550 888 4554 892
rect 4454 858 4458 862
rect 4470 858 4474 862
rect 4454 838 4458 842
rect 4462 818 4466 822
rect 4446 768 4450 772
rect 4454 768 4458 772
rect 4438 758 4442 762
rect 4390 738 4394 742
rect 4414 728 4418 732
rect 4398 688 4402 692
rect 4390 678 4394 682
rect 4406 658 4410 662
rect 4478 738 4482 742
rect 4454 708 4458 712
rect 4398 618 4402 622
rect 4426 603 4430 607
rect 4433 603 4437 607
rect 4358 578 4362 582
rect 4190 548 4194 552
rect 4286 548 4290 552
rect 4150 538 4154 542
rect 4166 538 4170 542
rect 4182 538 4186 542
rect 4142 518 4146 522
rect 4334 538 4338 542
rect 4446 538 4450 542
rect 4190 528 4194 532
rect 4246 528 4250 532
rect 4230 508 4234 512
rect 4438 508 4442 512
rect 4166 478 4170 482
rect 4350 478 4354 482
rect 4358 478 4362 482
rect 4374 478 4378 482
rect 4102 468 4106 472
rect 4150 468 4154 472
rect 4174 468 4178 472
rect 4198 468 4202 472
rect 4246 468 4250 472
rect 4334 468 4338 472
rect 4126 428 4130 432
rect 4182 448 4186 452
rect 4166 418 4170 422
rect 4214 458 4218 462
rect 4294 459 4298 463
rect 4198 448 4202 452
rect 4270 428 4274 432
rect 4190 408 4194 412
rect 4182 398 4186 402
rect 4142 388 4146 392
rect 4102 358 4106 362
rect 4166 378 4170 382
rect 4238 388 4242 392
rect 4206 358 4210 362
rect 4246 368 4250 372
rect 4254 368 4258 372
rect 4158 348 4162 352
rect 4182 348 4186 352
rect 4230 348 4234 352
rect 4182 338 4186 342
rect 4134 328 4138 332
rect 4182 328 4186 332
rect 4110 308 4114 312
rect 4102 248 4106 252
rect 4142 288 4146 292
rect 4342 368 4346 372
rect 4286 358 4290 362
rect 4366 468 4370 472
rect 4382 468 4386 472
rect 4398 458 4402 462
rect 4478 668 4482 672
rect 4542 878 4546 882
rect 4526 858 4530 862
rect 4502 848 4506 852
rect 4494 808 4498 812
rect 4502 788 4506 792
rect 4494 778 4498 782
rect 4510 708 4514 712
rect 4510 698 4514 702
rect 4590 918 4594 922
rect 4614 1118 4618 1122
rect 4606 1098 4610 1102
rect 4654 1138 4658 1142
rect 4654 1118 4658 1122
rect 4694 1118 4698 1122
rect 4638 1098 4642 1102
rect 4662 1098 4666 1102
rect 4622 1088 4626 1092
rect 4630 1068 4634 1072
rect 4638 1058 4642 1062
rect 4670 1088 4674 1092
rect 4614 1038 4618 1042
rect 4630 1038 4634 1042
rect 4646 1038 4650 1042
rect 4678 1028 4682 1032
rect 4638 1008 4642 1012
rect 4654 978 4658 982
rect 4646 968 4650 972
rect 4638 958 4642 962
rect 4614 948 4618 952
rect 4614 938 4618 942
rect 4598 898 4602 902
rect 4670 948 4674 952
rect 4710 1088 4714 1092
rect 4710 1068 4714 1072
rect 4694 948 4698 952
rect 4686 908 4690 912
rect 4614 888 4618 892
rect 4582 878 4586 882
rect 4590 878 4594 882
rect 4694 878 4698 882
rect 4750 1228 4754 1232
rect 4734 1198 4738 1202
rect 4742 1158 4746 1162
rect 4782 1168 4786 1172
rect 4742 1128 4746 1132
rect 4750 1108 4754 1112
rect 4758 1098 4762 1102
rect 4758 1088 4762 1092
rect 4726 1068 4730 1072
rect 4734 1068 4738 1072
rect 4902 1488 4906 1492
rect 4894 1478 4898 1482
rect 4886 1448 4890 1452
rect 4878 1438 4882 1442
rect 4902 1428 4906 1432
rect 4886 1368 4890 1372
rect 4854 1358 4858 1362
rect 4938 1503 4942 1507
rect 4945 1503 4949 1507
rect 4950 1488 4954 1492
rect 4926 1468 4930 1472
rect 4918 1458 4922 1462
rect 4934 1458 4938 1462
rect 4910 1408 4914 1412
rect 4918 1388 4922 1392
rect 4934 1368 4938 1372
rect 5070 1768 5074 1772
rect 5078 1758 5082 1762
rect 5022 1748 5026 1752
rect 5038 1748 5042 1752
rect 5030 1708 5034 1712
rect 5030 1648 5034 1652
rect 5054 1728 5058 1732
rect 5086 1728 5090 1732
rect 5078 1678 5082 1682
rect 5046 1668 5050 1672
rect 5070 1668 5074 1672
rect 5046 1658 5050 1662
rect 5086 1658 5090 1662
rect 5062 1648 5066 1652
rect 5038 1638 5042 1642
rect 5062 1628 5066 1632
rect 5030 1618 5034 1622
rect 4990 1578 4994 1582
rect 5022 1578 5026 1582
rect 4974 1518 4978 1522
rect 5054 1568 5058 1572
rect 5014 1548 5018 1552
rect 5038 1548 5042 1552
rect 5006 1458 5010 1462
rect 4990 1448 4994 1452
rect 4966 1428 4970 1432
rect 4950 1378 4954 1382
rect 5054 1488 5058 1492
rect 5054 1478 5058 1482
rect 5118 1778 5122 1782
rect 5110 1738 5114 1742
rect 5126 1688 5130 1692
rect 5126 1648 5130 1652
rect 5094 1618 5098 1622
rect 5110 1618 5114 1622
rect 5094 1608 5098 1612
rect 5070 1548 5074 1552
rect 5086 1548 5090 1552
rect 5078 1528 5082 1532
rect 5062 1458 5066 1462
rect 5078 1428 5082 1432
rect 4998 1408 5002 1412
rect 5038 1408 5042 1412
rect 5070 1408 5074 1412
rect 5062 1388 5066 1392
rect 5054 1368 5058 1372
rect 5046 1358 5050 1362
rect 5022 1348 5026 1352
rect 5038 1348 5042 1352
rect 5062 1358 5066 1362
rect 4926 1338 4930 1342
rect 4942 1338 4946 1342
rect 5006 1338 5010 1342
rect 5030 1338 5034 1342
rect 5046 1338 5050 1342
rect 4854 1288 4858 1292
rect 4982 1328 4986 1332
rect 4926 1318 4930 1322
rect 4938 1303 4942 1307
rect 4945 1303 4949 1307
rect 4958 1288 4962 1292
rect 5046 1318 5050 1322
rect 5014 1308 5018 1312
rect 5006 1288 5010 1292
rect 4990 1278 4994 1282
rect 4822 1268 4826 1272
rect 4870 1268 4874 1272
rect 4902 1268 4906 1272
rect 4982 1268 4986 1272
rect 4830 1158 4834 1162
rect 4862 1258 4866 1262
rect 4894 1258 4898 1262
rect 4902 1198 4906 1202
rect 4886 1178 4890 1182
rect 4902 1168 4906 1172
rect 4870 1158 4874 1162
rect 4894 1158 4898 1162
rect 5102 1468 5106 1472
rect 5102 1368 5106 1372
rect 5094 1358 5098 1362
rect 5190 1908 5194 1912
rect 5166 1898 5170 1902
rect 5158 1878 5162 1882
rect 5166 1878 5170 1882
rect 5182 1868 5186 1872
rect 5206 1828 5210 1832
rect 5166 1768 5170 1772
rect 5142 1568 5146 1572
rect 5262 1938 5266 1942
rect 5222 1908 5226 1912
rect 5238 1908 5242 1912
rect 5230 1868 5234 1872
rect 5222 1848 5226 1852
rect 5214 1748 5218 1752
rect 5230 1748 5234 1752
rect 5174 1738 5178 1742
rect 5286 1978 5290 1982
rect 5278 1948 5282 1952
rect 5278 1898 5282 1902
rect 5278 1868 5282 1872
rect 5198 1688 5202 1692
rect 5254 1688 5258 1692
rect 5190 1668 5194 1672
rect 5238 1668 5242 1672
rect 5262 1668 5266 1672
rect 5166 1658 5170 1662
rect 5222 1658 5226 1662
rect 5238 1658 5242 1662
rect 5182 1648 5186 1652
rect 5134 1548 5138 1552
rect 5150 1548 5154 1552
rect 5150 1538 5154 1542
rect 5150 1508 5154 1512
rect 5118 1458 5122 1462
rect 5206 1508 5210 1512
rect 5190 1478 5194 1482
rect 5198 1478 5202 1482
rect 5150 1458 5154 1462
rect 5174 1458 5178 1462
rect 5198 1458 5202 1462
rect 5134 1448 5138 1452
rect 5126 1438 5130 1442
rect 5086 1348 5090 1352
rect 5094 1338 5098 1342
rect 5086 1318 5090 1322
rect 5094 1308 5098 1312
rect 5110 1308 5114 1312
rect 5078 1298 5082 1302
rect 5070 1288 5074 1292
rect 5054 1268 5058 1272
rect 4998 1258 5002 1262
rect 4918 1248 4922 1252
rect 4918 1158 4922 1162
rect 5054 1248 5058 1252
rect 4998 1188 5002 1192
rect 4982 1158 4986 1162
rect 5046 1158 5050 1162
rect 4966 1148 4970 1152
rect 5054 1148 5058 1152
rect 4894 1128 4898 1132
rect 4886 1118 4890 1122
rect 4846 1088 4850 1092
rect 4894 1078 4898 1082
rect 4798 1058 4802 1062
rect 4870 1058 4874 1062
rect 4886 1058 4890 1062
rect 4830 1048 4834 1052
rect 4878 1048 4882 1052
rect 4790 1008 4794 1012
rect 4806 968 4810 972
rect 4750 958 4754 962
rect 4862 1038 4866 1042
rect 4838 1028 4842 1032
rect 4854 968 4858 972
rect 4782 948 4786 952
rect 4742 928 4746 932
rect 4734 918 4738 922
rect 4742 918 4746 922
rect 4766 878 4770 882
rect 4606 868 4610 872
rect 4678 868 4682 872
rect 4702 868 4706 872
rect 4718 868 4722 872
rect 4614 848 4618 852
rect 4638 838 4642 842
rect 4638 818 4642 822
rect 4662 838 4666 842
rect 4614 798 4618 802
rect 4654 798 4658 802
rect 4574 758 4578 762
rect 4606 758 4610 762
rect 4550 748 4554 752
rect 4574 748 4578 752
rect 4542 708 4546 712
rect 4558 708 4562 712
rect 4590 678 4594 682
rect 4566 668 4570 672
rect 4502 658 4506 662
rect 4526 658 4530 662
rect 4550 658 4554 662
rect 4486 608 4490 612
rect 4510 578 4514 582
rect 4622 748 4626 752
rect 4582 658 4586 662
rect 4606 658 4610 662
rect 4646 738 4650 742
rect 4654 718 4658 722
rect 4654 678 4658 682
rect 4670 678 4674 682
rect 4638 648 4642 652
rect 4630 638 4634 642
rect 4742 828 4746 832
rect 4718 818 4722 822
rect 4694 728 4698 732
rect 4686 668 4690 672
rect 4654 608 4658 612
rect 4646 598 4650 602
rect 4598 588 4602 592
rect 4598 568 4602 572
rect 4638 568 4642 572
rect 4518 548 4522 552
rect 4566 548 4570 552
rect 4582 548 4586 552
rect 4630 548 4634 552
rect 4470 538 4474 542
rect 4534 538 4538 542
rect 4534 528 4538 532
rect 4510 518 4514 522
rect 4478 508 4482 512
rect 4470 498 4474 502
rect 4510 488 4514 492
rect 4518 478 4522 482
rect 4590 508 4594 512
rect 4606 488 4610 492
rect 4622 488 4626 492
rect 4646 508 4650 512
rect 4574 468 4578 472
rect 4494 458 4498 462
rect 4566 458 4570 462
rect 4406 448 4410 452
rect 4406 388 4410 392
rect 4390 358 4394 362
rect 4358 348 4362 352
rect 4398 348 4402 352
rect 4350 338 4354 342
rect 4198 308 4202 312
rect 4230 288 4234 292
rect 4174 268 4178 272
rect 4158 258 4162 262
rect 4190 258 4194 262
rect 4206 258 4210 262
rect 4214 258 4218 262
rect 4246 248 4250 252
rect 4278 248 4282 252
rect 4374 318 4378 322
rect 4334 288 4338 292
rect 4366 288 4370 292
rect 4350 278 4354 282
rect 4398 288 4402 292
rect 4382 278 4386 282
rect 4494 448 4498 452
rect 4518 448 4522 452
rect 4534 448 4538 452
rect 4438 428 4442 432
rect 4426 403 4430 407
rect 4433 403 4437 407
rect 4454 358 4458 362
rect 4310 258 4314 262
rect 4422 258 4426 262
rect 4366 248 4370 252
rect 4398 248 4402 252
rect 4174 238 4178 242
rect 4222 238 4226 242
rect 4294 238 4298 242
rect 4206 208 4210 212
rect 4142 188 4146 192
rect 4126 168 4130 172
rect 4102 158 4106 162
rect 4110 158 4114 162
rect 4118 88 4122 92
rect 4382 218 4386 222
rect 4430 218 4434 222
rect 4406 208 4410 212
rect 4426 203 4430 207
rect 4433 203 4437 207
rect 4374 168 4378 172
rect 4414 168 4418 172
rect 4446 168 4450 172
rect 4270 148 4274 152
rect 4302 148 4306 152
rect 4150 108 4154 112
rect 4174 98 4178 102
rect 4182 98 4186 102
rect 4254 98 4258 102
rect 4094 78 4098 82
rect 4126 78 4130 82
rect 4246 88 4250 92
rect 4262 78 4266 82
rect 4206 68 4210 72
rect 4286 138 4290 142
rect 4294 108 4298 112
rect 4286 88 4290 92
rect 4502 328 4506 332
rect 4494 268 4498 272
rect 4510 318 4514 322
rect 4518 288 4522 292
rect 4542 428 4546 432
rect 4622 428 4626 432
rect 4590 348 4594 352
rect 4542 318 4546 322
rect 4542 288 4546 292
rect 4582 308 4586 312
rect 4542 278 4546 282
rect 4566 258 4570 262
rect 4534 248 4538 252
rect 4566 248 4570 252
rect 4542 238 4546 242
rect 4510 228 4514 232
rect 4478 168 4482 172
rect 4518 158 4522 162
rect 4318 138 4322 142
rect 4366 128 4370 132
rect 4326 118 4330 122
rect 4302 78 4306 82
rect 4334 98 4338 102
rect 4406 108 4410 112
rect 4486 98 4490 102
rect 4414 88 4418 92
rect 4398 78 4402 82
rect 4550 158 4554 162
rect 4606 258 4610 262
rect 4590 248 4594 252
rect 4582 188 4586 192
rect 4590 178 4594 182
rect 4598 168 4602 172
rect 4654 448 4658 452
rect 4774 758 4778 762
rect 4774 728 4778 732
rect 4758 708 4762 712
rect 4670 658 4674 662
rect 4718 658 4722 662
rect 4670 548 4674 552
rect 4702 628 4706 632
rect 4734 618 4738 622
rect 4766 608 4770 612
rect 4718 578 4722 582
rect 4702 528 4706 532
rect 4750 528 4754 532
rect 4686 468 4690 472
rect 4718 468 4722 472
rect 4646 388 4650 392
rect 4638 368 4642 372
rect 4638 348 4642 352
rect 4654 318 4658 322
rect 4662 308 4666 312
rect 4646 298 4650 302
rect 4678 448 4682 452
rect 4686 438 4690 442
rect 4750 468 4754 472
rect 4734 448 4738 452
rect 4718 398 4722 402
rect 4758 448 4762 452
rect 4750 428 4754 432
rect 4838 938 4842 942
rect 4878 948 4882 952
rect 4862 938 4866 942
rect 4918 1138 4922 1142
rect 4934 1138 4938 1142
rect 4950 1118 4954 1122
rect 4938 1103 4942 1107
rect 4945 1103 4949 1107
rect 4910 1088 4914 1092
rect 4982 1138 4986 1142
rect 4918 958 4922 962
rect 4934 958 4938 962
rect 4926 948 4930 952
rect 4974 1048 4978 1052
rect 5038 1138 5042 1142
rect 5006 1108 5010 1112
rect 5014 1098 5018 1102
rect 5110 1278 5114 1282
rect 5094 1248 5098 1252
rect 5102 1218 5106 1222
rect 5238 1538 5242 1542
rect 5238 1518 5242 1522
rect 5246 1468 5250 1472
rect 5222 1458 5226 1462
rect 5206 1438 5210 1442
rect 5158 1418 5162 1422
rect 5206 1398 5210 1402
rect 5182 1358 5186 1362
rect 5142 1348 5146 1352
rect 5182 1348 5186 1352
rect 5246 1348 5250 1352
rect 5142 1338 5146 1342
rect 5198 1338 5202 1342
rect 5222 1328 5226 1332
rect 5206 1318 5210 1322
rect 5150 1298 5154 1302
rect 5126 1268 5130 1272
rect 5118 1208 5122 1212
rect 5118 1168 5122 1172
rect 5086 1108 5090 1112
rect 5110 1148 5114 1152
rect 5214 1308 5218 1312
rect 5190 1258 5194 1262
rect 5174 1228 5178 1232
rect 5158 1218 5162 1222
rect 5150 1198 5154 1202
rect 5134 1168 5138 1172
rect 5166 1158 5170 1162
rect 5246 1268 5250 1272
rect 5214 1178 5218 1182
rect 5190 1148 5194 1152
rect 5110 1138 5114 1142
rect 5118 1138 5122 1142
rect 5102 1098 5106 1102
rect 5126 1128 5130 1132
rect 5150 1128 5154 1132
rect 5094 1078 5098 1082
rect 5078 1068 5082 1072
rect 5014 978 5018 982
rect 5054 968 5058 972
rect 4998 958 5002 962
rect 4998 948 5002 952
rect 5038 948 5042 952
rect 4918 938 4922 942
rect 4966 938 4970 942
rect 4910 928 4914 932
rect 4798 888 4802 892
rect 4878 918 4882 922
rect 4822 888 4826 892
rect 4838 878 4842 882
rect 4942 928 4946 932
rect 5038 928 5042 932
rect 4958 918 4962 922
rect 5014 918 5018 922
rect 4938 903 4942 907
rect 4945 903 4949 907
rect 4934 888 4938 892
rect 4958 888 4962 892
rect 4998 878 5002 882
rect 4902 868 4906 872
rect 4966 868 4970 872
rect 5062 948 5066 952
rect 5054 908 5058 912
rect 5078 908 5082 912
rect 5158 1088 5162 1092
rect 5134 1068 5138 1072
rect 5158 1068 5162 1072
rect 5166 1068 5170 1072
rect 5134 1048 5138 1052
rect 5150 988 5154 992
rect 5102 948 5106 952
rect 5134 948 5138 952
rect 5150 888 5154 892
rect 5006 868 5010 872
rect 5206 1138 5210 1142
rect 5198 1068 5202 1072
rect 5198 1038 5202 1042
rect 5190 1018 5194 1022
rect 5190 968 5194 972
rect 5206 948 5210 952
rect 5206 938 5210 942
rect 5166 878 5170 882
rect 5158 868 5162 872
rect 5206 868 5210 872
rect 5054 858 5058 862
rect 5086 858 5090 862
rect 5126 858 5130 862
rect 5182 858 5186 862
rect 5198 858 5202 862
rect 4998 848 5002 852
rect 5030 848 5034 852
rect 4918 838 4922 842
rect 5022 838 5026 842
rect 4830 778 4834 782
rect 4814 768 4818 772
rect 4894 768 4898 772
rect 4790 748 4794 752
rect 4798 748 4802 752
rect 4878 748 4882 752
rect 4790 718 4794 722
rect 4790 698 4794 702
rect 4806 668 4810 672
rect 4854 688 4858 692
rect 4878 698 4882 702
rect 4910 678 4914 682
rect 4902 668 4906 672
rect 5102 848 5106 852
rect 5014 828 5018 832
rect 5046 828 5050 832
rect 4966 808 4970 812
rect 4958 778 4962 782
rect 4926 728 4930 732
rect 4950 718 4954 722
rect 4938 703 4942 707
rect 4945 703 4949 707
rect 4934 688 4938 692
rect 5094 758 5098 762
rect 4974 748 4978 752
rect 5030 748 5034 752
rect 4966 738 4970 742
rect 4998 738 5002 742
rect 5006 728 5010 732
rect 4982 718 4986 722
rect 4998 698 5002 702
rect 4990 688 4994 692
rect 5006 678 5010 682
rect 5046 748 5050 752
rect 5078 748 5082 752
rect 5038 728 5042 732
rect 5022 718 5026 722
rect 5062 718 5066 722
rect 5094 718 5098 722
rect 5014 668 5018 672
rect 4870 658 4874 662
rect 4918 658 4922 662
rect 4958 658 4962 662
rect 5062 678 5066 682
rect 5038 658 5042 662
rect 5062 658 5066 662
rect 4830 648 4834 652
rect 4806 618 4810 622
rect 4822 618 4826 622
rect 4798 608 4802 612
rect 4798 538 4802 542
rect 4790 458 4794 462
rect 4782 368 4786 372
rect 4678 348 4682 352
rect 4702 348 4706 352
rect 4718 348 4722 352
rect 4742 348 4746 352
rect 4750 338 4754 342
rect 4678 308 4682 312
rect 4670 278 4674 282
rect 4630 268 4634 272
rect 4702 308 4706 312
rect 4734 318 4738 322
rect 4718 278 4722 282
rect 4814 338 4818 342
rect 4790 328 4794 332
rect 4766 318 4770 322
rect 4758 288 4762 292
rect 4782 278 4786 282
rect 4742 268 4746 272
rect 4694 258 4698 262
rect 4654 208 4658 212
rect 4638 168 4642 172
rect 4638 138 4642 142
rect 4614 128 4618 132
rect 4598 118 4602 122
rect 4566 88 4570 92
rect 4622 88 4626 92
rect 4454 78 4458 82
rect 4590 78 4594 82
rect 4422 68 4426 72
rect 4446 68 4450 72
rect 4486 68 4490 72
rect 4550 68 4554 72
rect 4718 258 4722 262
rect 4806 298 4810 302
rect 4782 248 4786 252
rect 4774 238 4778 242
rect 4806 228 4810 232
rect 4806 218 4810 222
rect 4718 168 4722 172
rect 4766 168 4770 172
rect 4782 168 4786 172
rect 4710 158 4714 162
rect 4694 148 4698 152
rect 4750 158 4754 162
rect 4758 148 4762 152
rect 4734 138 4738 142
rect 4766 138 4770 142
rect 4766 128 4770 132
rect 4782 88 4786 92
rect 4750 78 4754 82
rect 4638 68 4642 72
rect 4798 98 4802 102
rect 4814 158 4818 162
rect 4934 648 4938 652
rect 4950 648 4954 652
rect 5006 648 5010 652
rect 5038 648 5042 652
rect 5046 648 5050 652
rect 5086 648 5090 652
rect 4982 628 4986 632
rect 5030 638 5034 642
rect 4982 558 4986 562
rect 5030 558 5034 562
rect 4926 548 4930 552
rect 4982 548 4986 552
rect 4998 538 5002 542
rect 4934 528 4938 532
rect 4894 508 4898 512
rect 4958 508 4962 512
rect 4938 503 4942 507
rect 4945 503 4949 507
rect 4918 498 4922 502
rect 4918 488 4922 492
rect 4870 478 4874 482
rect 4886 478 4890 482
rect 4830 468 4834 472
rect 4830 458 4834 462
rect 4926 478 4930 482
rect 4958 478 4962 482
rect 4870 458 4874 462
rect 4894 448 4898 452
rect 4958 448 4962 452
rect 4974 448 4978 452
rect 4878 418 4882 422
rect 4886 378 4890 382
rect 4910 378 4914 382
rect 4878 358 4882 362
rect 4870 328 4874 332
rect 4846 268 4850 272
rect 4830 258 4834 262
rect 5006 528 5010 532
rect 5030 528 5034 532
rect 5022 518 5026 522
rect 5030 508 5034 512
rect 5038 508 5042 512
rect 5006 448 5010 452
rect 4982 418 4986 422
rect 4902 348 4906 352
rect 4942 328 4946 332
rect 4966 328 4970 332
rect 4950 318 4954 322
rect 4938 303 4942 307
rect 4945 303 4949 307
rect 4926 268 4930 272
rect 4902 258 4906 262
rect 4990 368 4994 372
rect 5014 368 5018 372
rect 5070 628 5074 632
rect 5126 798 5130 802
rect 5126 778 5130 782
rect 5118 748 5122 752
rect 5126 698 5130 702
rect 5110 658 5114 662
rect 5110 568 5114 572
rect 5086 548 5090 552
rect 5078 538 5082 542
rect 5054 518 5058 522
rect 5102 518 5106 522
rect 5062 508 5066 512
rect 5094 508 5098 512
rect 5094 488 5098 492
rect 5046 478 5050 482
rect 5070 468 5074 472
rect 5046 458 5050 462
rect 5070 458 5074 462
rect 5078 448 5082 452
rect 4998 348 5002 352
rect 5070 348 5074 352
rect 4982 338 4986 342
rect 5014 338 5018 342
rect 5006 288 5010 292
rect 5038 288 5042 292
rect 4990 278 4994 282
rect 4974 268 4978 272
rect 5006 258 5010 262
rect 5014 258 5018 262
rect 4974 248 4978 252
rect 4990 218 4994 222
rect 4926 178 4930 182
rect 5006 248 5010 252
rect 5070 248 5074 252
rect 5086 218 5090 222
rect 5022 198 5026 202
rect 4998 188 5002 192
rect 4990 168 4994 172
rect 5014 168 5018 172
rect 5062 188 5066 192
rect 5086 188 5090 192
rect 5030 168 5034 172
rect 5030 158 5034 162
rect 5038 158 5042 162
rect 4878 148 4882 152
rect 5070 148 5074 152
rect 5022 138 5026 142
rect 4894 128 4898 132
rect 4950 118 4954 122
rect 4938 103 4942 107
rect 4945 103 4949 107
rect 5102 468 5106 472
rect 5118 528 5122 532
rect 5158 818 5162 822
rect 5158 808 5162 812
rect 5150 768 5154 772
rect 5166 788 5170 792
rect 5158 748 5162 752
rect 5174 748 5178 752
rect 5158 728 5162 732
rect 5166 688 5170 692
rect 5150 678 5154 682
rect 5166 648 5170 652
rect 5150 568 5154 572
rect 5166 548 5170 552
rect 5198 738 5202 742
rect 5182 578 5186 582
rect 5206 558 5210 562
rect 5190 548 5194 552
rect 5166 538 5170 542
rect 5174 538 5178 542
rect 5182 538 5186 542
rect 5262 1178 5266 1182
rect 5294 1758 5298 1762
rect 5302 1368 5306 1372
rect 5286 1188 5290 1192
rect 5270 1148 5274 1152
rect 5254 1138 5258 1142
rect 5246 1068 5250 1072
rect 5278 1018 5282 1022
rect 5222 988 5226 992
rect 5262 988 5266 992
rect 5270 988 5274 992
rect 5238 918 5242 922
rect 5286 958 5290 962
rect 5286 948 5290 952
rect 5246 908 5250 912
rect 5238 868 5242 872
rect 5246 868 5250 872
rect 5222 758 5226 762
rect 5262 898 5266 902
rect 5278 818 5282 822
rect 5254 768 5258 772
rect 5262 728 5266 732
rect 5278 728 5282 732
rect 5246 668 5250 672
rect 5254 608 5258 612
rect 5294 598 5298 602
rect 5182 528 5186 532
rect 5214 528 5218 532
rect 5142 518 5146 522
rect 5174 518 5178 522
rect 5158 508 5162 512
rect 5126 458 5130 462
rect 5102 438 5106 442
rect 5166 458 5170 462
rect 5142 418 5146 422
rect 5142 408 5146 412
rect 5158 408 5162 412
rect 5134 398 5138 402
rect 5166 378 5170 382
rect 5134 328 5138 332
rect 5142 298 5146 302
rect 5126 288 5130 292
rect 5166 338 5170 342
rect 5214 488 5218 492
rect 5198 448 5202 452
rect 5198 418 5202 422
rect 5190 388 5194 392
rect 5182 358 5186 362
rect 5182 328 5186 332
rect 5142 278 5146 282
rect 5150 278 5154 282
rect 5270 538 5274 542
rect 5270 528 5274 532
rect 5262 488 5266 492
rect 5222 468 5226 472
rect 5270 468 5274 472
rect 5278 458 5282 462
rect 5238 398 5242 402
rect 5286 388 5290 392
rect 5262 368 5266 372
rect 5246 348 5250 352
rect 5222 338 5226 342
rect 5214 328 5218 332
rect 5278 338 5282 342
rect 5238 318 5242 322
rect 5206 308 5210 312
rect 5230 308 5234 312
rect 5246 298 5250 302
rect 5214 288 5218 292
rect 5222 278 5226 282
rect 5246 278 5250 282
rect 5166 268 5170 272
rect 5238 268 5242 272
rect 5182 258 5186 262
rect 5142 208 5146 212
rect 5222 218 5226 222
rect 5198 198 5202 202
rect 5270 318 5274 322
rect 5278 308 5282 312
rect 5294 328 5298 332
rect 5286 298 5290 302
rect 5278 278 5282 282
rect 5254 268 5258 272
rect 5278 268 5282 272
rect 5286 258 5290 262
rect 5230 188 5234 192
rect 5158 178 5162 182
rect 5126 148 5130 152
rect 5230 158 5234 162
rect 5246 158 5250 162
rect 5110 138 5114 142
rect 4838 88 4842 92
rect 4934 88 4938 92
rect 4790 78 4794 82
rect 4830 78 4834 82
rect 4910 78 4914 82
rect 5038 78 5042 82
rect 5174 128 5178 132
rect 5214 78 5218 82
rect 5102 68 5106 72
rect 4070 58 4074 62
rect 4246 58 4250 62
rect 4286 58 4290 62
rect 4382 58 4386 62
rect 4414 58 4418 62
rect 4422 58 4426 62
rect 4622 58 4626 62
rect 4646 58 4650 62
rect 4710 58 4714 62
rect 4790 58 4794 62
rect 4886 59 4890 63
rect 4998 59 5002 63
rect 1494 48 1498 52
rect 2230 48 2234 52
rect 3654 48 3658 52
rect 3806 48 3810 52
rect 4094 48 4098 52
rect 4454 48 4458 52
rect 5278 148 5282 152
rect 5262 138 5266 142
rect 5286 68 5290 72
rect 5174 58 5178 62
rect 4774 48 4778 52
rect 5022 48 5026 52
rect 5174 48 5178 52
rect 5198 48 5202 52
rect 710 38 714 42
rect 822 38 826 42
rect 1350 38 1354 42
rect 3750 38 3754 42
rect 4086 38 4090 42
rect 4606 38 4610 42
rect 2230 8 2234 12
rect 4526 8 4530 12
rect 330 3 334 7
rect 337 3 341 7
rect 1354 3 1358 7
rect 1361 3 1365 7
rect 2386 3 2390 7
rect 2393 3 2397 7
rect 3402 3 3406 7
rect 3409 3 3413 7
rect 4426 3 4430 7
rect 4433 3 4437 7
<< metal3 >>
rect 848 5103 850 5107
rect 854 5103 857 5107
rect 862 5103 864 5107
rect 1872 5103 1874 5107
rect 1878 5103 1881 5107
rect 1886 5103 1888 5107
rect 2888 5103 2890 5107
rect 2894 5103 2897 5107
rect 2902 5103 2904 5107
rect 3920 5103 3922 5107
rect 3926 5103 3929 5107
rect 3934 5103 3936 5107
rect 4936 5103 4938 5107
rect 4942 5103 4945 5107
rect 4950 5103 4952 5107
rect 314 5098 318 5101
rect 1658 5098 1662 5101
rect 514 5088 654 5091
rect 754 5088 814 5091
rect 2314 5088 2454 5091
rect 2530 5088 2614 5091
rect 2618 5088 2750 5091
rect 4154 5088 4238 5091
rect 114 5078 150 5081
rect 178 5078 294 5081
rect 306 5078 318 5081
rect 322 5078 382 5081
rect 702 5081 705 5088
rect 562 5078 705 5081
rect 802 5078 822 5081
rect 826 5078 910 5081
rect 1126 5081 1129 5088
rect 1126 5078 1134 5081
rect 1230 5081 1233 5088
rect 4486 5082 4489 5088
rect 1138 5078 1233 5081
rect 1726 5078 1734 5081
rect 1738 5078 1822 5081
rect 1826 5078 1934 5081
rect 2434 5078 2462 5081
rect 4498 5078 4502 5081
rect 5026 5078 5206 5081
rect 42 5068 193 5071
rect 314 5068 318 5071
rect 658 5068 694 5071
rect 722 5068 742 5071
rect 746 5068 846 5071
rect 1122 5068 1134 5071
rect 1242 5068 1270 5071
rect 1538 5068 1542 5071
rect 1546 5068 1590 5071
rect 1594 5068 1662 5071
rect 1666 5068 1734 5071
rect 2126 5071 2129 5078
rect 1986 5068 2129 5071
rect 2250 5068 2406 5071
rect 2450 5068 2486 5071
rect 2514 5068 2558 5071
rect 2666 5068 2742 5071
rect 3026 5068 3078 5071
rect 3122 5068 3150 5071
rect 3186 5068 3262 5071
rect 3474 5068 3566 5071
rect 3930 5068 3958 5071
rect 3962 5068 4030 5071
rect 4034 5068 4390 5071
rect 4394 5068 4854 5071
rect 5014 5071 5017 5078
rect 5014 5068 5046 5071
rect 5050 5068 5166 5071
rect 5170 5068 5238 5071
rect 190 5062 193 5068
rect 58 5058 118 5061
rect 154 5058 158 5061
rect 170 5058 174 5061
rect 210 5059 214 5061
rect 210 5058 217 5059
rect 450 5058 462 5061
rect 466 5058 470 5061
rect 562 5058 566 5061
rect 570 5058 582 5061
rect 666 5058 774 5061
rect 842 5058 870 5061
rect 1058 5058 1182 5061
rect 1190 5061 1193 5068
rect 1190 5058 1270 5061
rect 1406 5061 1409 5068
rect 1406 5058 1478 5061
rect 1578 5058 1782 5061
rect 1802 5058 2062 5061
rect 2066 5058 2222 5061
rect 2226 5058 2318 5061
rect 2322 5058 2502 5061
rect 2506 5058 2542 5061
rect 2546 5058 2638 5061
rect 2642 5058 2790 5061
rect 2826 5058 2894 5061
rect 3074 5058 3198 5061
rect 3366 5061 3369 5068
rect 3366 5058 3446 5061
rect 3546 5058 3574 5061
rect 3578 5058 3670 5061
rect 3766 5061 3769 5068
rect 3710 5058 3769 5061
rect 4082 5058 4086 5061
rect 4226 5058 4406 5061
rect 4594 5058 4782 5061
rect 4786 5058 4902 5061
rect 5002 5058 5022 5061
rect 5058 5058 5238 5061
rect 5242 5058 5246 5061
rect 130 5048 294 5051
rect 386 5048 462 5051
rect 506 5048 542 5051
rect 546 5048 761 5051
rect 830 5051 833 5058
rect 3710 5052 3713 5058
rect 3950 5052 3953 5058
rect 4310 5052 4313 5058
rect 4574 5052 4577 5058
rect 4926 5052 4929 5058
rect 794 5048 833 5051
rect 938 5048 1070 5051
rect 1078 5048 1230 5051
rect 1234 5048 1246 5051
rect 2154 5048 2350 5051
rect 2458 5048 2614 5051
rect 2778 5048 3054 5051
rect 3126 5048 3158 5051
rect 3178 5048 3214 5051
rect 3218 5048 3278 5051
rect 3346 5048 3558 5051
rect 3730 5048 3838 5051
rect 4906 5048 4910 5051
rect 4986 5048 5014 5051
rect 5334 5051 5338 5052
rect 5306 5048 5338 5051
rect 758 5042 761 5048
rect 1078 5042 1081 5048
rect 3126 5042 3129 5048
rect 442 5038 454 5041
rect 602 5038 622 5041
rect 626 5038 737 5041
rect 810 5038 822 5041
rect 1098 5038 1334 5041
rect 2346 5038 2454 5041
rect 2490 5038 2510 5041
rect 2514 5038 2742 5041
rect 2746 5038 2766 5041
rect 2770 5038 3097 5041
rect 3170 5038 3182 5041
rect 3202 5038 3262 5041
rect 3434 5038 3694 5041
rect 3706 5038 3718 5041
rect 4290 5038 4566 5041
rect 4690 5038 5014 5041
rect 734 5032 737 5038
rect 370 5028 494 5031
rect 610 5028 662 5031
rect 746 5028 942 5031
rect 954 5028 1038 5031
rect 1042 5028 1382 5031
rect 2090 5028 2518 5031
rect 2970 5028 2998 5031
rect 3002 5028 3086 5031
rect 3094 5031 3097 5038
rect 3094 5028 4014 5031
rect 4210 5028 4342 5031
rect 4402 5028 4782 5031
rect 226 5018 414 5021
rect 418 5018 470 5021
rect 474 5018 486 5021
rect 1914 5018 1958 5021
rect 2034 5018 2262 5021
rect 2410 5018 2430 5021
rect 2442 5018 2446 5021
rect 2450 5018 2638 5021
rect 2730 5018 2958 5021
rect 3042 5018 3166 5021
rect 3690 5018 3734 5021
rect 3738 5018 3998 5021
rect 4138 5018 4142 5021
rect 4522 5018 4526 5021
rect 4970 5018 5054 5021
rect 5146 5018 5150 5021
rect 926 5012 929 5018
rect 410 5008 502 5011
rect 538 5008 926 5011
rect 946 5008 1046 5011
rect 1658 5008 2302 5011
rect 2946 5008 3214 5011
rect 3474 5008 3494 5011
rect 3498 5008 3654 5011
rect 3658 5008 3766 5011
rect 328 5003 330 5007
rect 334 5003 337 5007
rect 342 5003 344 5007
rect 1352 5003 1354 5007
rect 1358 5003 1361 5007
rect 1366 5003 1368 5007
rect 2384 5003 2386 5007
rect 2390 5003 2393 5007
rect 2398 5003 2400 5007
rect 3400 5003 3402 5007
rect 3406 5003 3409 5007
rect 3414 5003 3416 5007
rect 4424 5003 4426 5007
rect 4430 5003 4433 5007
rect 4438 5003 4440 5007
rect 378 4998 494 5001
rect 498 4998 614 5001
rect 898 4998 942 5001
rect 946 4998 1254 5001
rect 1258 4998 1278 5001
rect 1658 4998 1662 5001
rect 1850 4998 1942 5001
rect 1970 4998 2134 5001
rect 2482 4998 3206 5001
rect 3562 4998 3702 5001
rect 3842 4998 4302 5001
rect 4482 4998 4758 5001
rect 3550 4992 3553 4998
rect 18 4988 534 4991
rect 2210 4988 2390 4991
rect 3154 4988 3310 4991
rect 3802 4988 3846 4991
rect 458 4978 502 4981
rect 778 4978 862 4981
rect 866 4978 894 4981
rect 958 4981 961 4988
rect 898 4978 961 4981
rect 2410 4978 2558 4981
rect 2794 4978 3046 4981
rect 3058 4978 3150 4981
rect 3234 4978 3350 4981
rect 3354 4978 3462 4981
rect 3562 4978 3630 4981
rect 3634 4978 4190 4981
rect 4362 4978 4526 4981
rect 4530 4978 4558 4981
rect 226 4968 278 4971
rect 442 4968 486 4971
rect 534 4971 537 4978
rect 490 4968 537 4971
rect 730 4968 734 4971
rect 746 4968 838 4971
rect 850 4968 886 4971
rect 978 4968 1006 4971
rect 1266 4968 1294 4971
rect 1458 4968 1542 4971
rect 2150 4968 2582 4971
rect 2866 4968 2894 4971
rect 2930 4968 3110 4971
rect 3258 4968 3294 4971
rect 3442 4968 3534 4971
rect 3542 4971 3545 4978
rect 3542 4968 3558 4971
rect 4250 4968 4358 4971
rect 4362 4968 4422 4971
rect 4610 4968 4614 4971
rect 4762 4968 4806 4971
rect 5010 4968 5118 4971
rect 286 4962 289 4968
rect 266 4958 278 4961
rect 298 4958 374 4961
rect 394 4958 422 4961
rect 426 4958 454 4961
rect 474 4958 478 4961
rect 622 4961 625 4968
rect 490 4958 625 4961
rect 630 4958 814 4961
rect 818 4958 830 4961
rect 902 4961 905 4968
rect 834 4958 905 4961
rect 950 4961 953 4968
rect 2150 4962 2153 4968
rect 938 4958 953 4961
rect 970 4958 1222 4961
rect 1226 4958 1270 4961
rect 1274 4958 1350 4961
rect 1354 4958 1390 4961
rect 1930 4958 1934 4961
rect 2082 4958 2150 4961
rect 2202 4958 2214 4961
rect 2218 4958 2222 4961
rect 2418 4958 2566 4961
rect 2626 4958 2630 4961
rect 2662 4961 2665 4968
rect 2662 4958 2694 4961
rect 3130 4958 3302 4961
rect 3306 4958 3334 4961
rect 3338 4958 3510 4961
rect 3514 4958 3542 4961
rect 3662 4961 3665 4968
rect 3658 4958 3665 4961
rect 3794 4958 3862 4961
rect 4074 4958 4230 4961
rect 4522 4958 4542 4961
rect 4610 4958 4806 4961
rect 5042 4958 5086 4961
rect 158 4951 161 4958
rect 146 4948 161 4951
rect 186 4948 190 4951
rect 210 4948 214 4951
rect 242 4948 246 4951
rect 250 4948 326 4951
rect 354 4948 366 4951
rect 370 4948 518 4951
rect 630 4951 633 4958
rect 610 4948 633 4951
rect 762 4948 918 4951
rect 922 4948 990 4951
rect 1066 4948 1166 4951
rect 1226 4948 1302 4951
rect 1346 4948 1406 4951
rect 1430 4948 1438 4951
rect 1442 4948 1454 4951
rect 1474 4948 1497 4951
rect 1590 4951 1593 4958
rect 1710 4951 1713 4958
rect 1522 4948 1713 4951
rect 1730 4948 1734 4951
rect 2018 4948 2070 4951
rect 2138 4948 2182 4951
rect 2194 4948 2238 4951
rect 2246 4948 2318 4951
rect 2338 4948 2350 4951
rect 2354 4948 2438 4951
rect 2442 4948 2470 4951
rect 2498 4948 2526 4951
rect 2530 4948 2550 4951
rect 2622 4951 2625 4958
rect 2570 4948 2625 4951
rect 2650 4948 2870 4951
rect 2874 4948 2942 4951
rect 3118 4951 3121 4958
rect 3010 4948 3121 4951
rect 3202 4948 3278 4951
rect 3290 4948 3366 4951
rect 1494 4942 1497 4948
rect 74 4938 118 4941
rect 122 4938 185 4941
rect 250 4938 270 4941
rect 274 4938 310 4941
rect 362 4938 366 4941
rect 394 4938 446 4941
rect 466 4938 558 4941
rect 578 4938 638 4941
rect 642 4938 766 4941
rect 778 4938 785 4941
rect 794 4938 806 4941
rect 834 4938 1014 4941
rect 1138 4938 1174 4941
rect 1402 4938 1489 4941
rect 1658 4938 1894 4941
rect 2194 4938 2217 4941
rect 2246 4941 2249 4948
rect 3490 4948 3550 4951
rect 3618 4948 3654 4951
rect 3698 4948 3702 4951
rect 3786 4948 3878 4951
rect 4070 4951 4073 4958
rect 3986 4948 4073 4951
rect 4098 4948 4134 4951
rect 4170 4948 4246 4951
rect 4322 4948 4494 4951
rect 4530 4948 4593 4951
rect 4642 4948 4710 4951
rect 4786 4948 4798 4951
rect 4870 4951 4873 4958
rect 4870 4948 4918 4951
rect 4978 4948 5302 4951
rect 3574 4942 3577 4948
rect 3590 4942 3593 4948
rect 3726 4942 3729 4948
rect 4590 4942 4593 4948
rect 2226 4938 2249 4941
rect 2330 4938 2510 4941
rect 2546 4938 2638 4941
rect 2882 4938 2926 4941
rect 3082 4938 3126 4941
rect 3210 4938 3246 4941
rect 3266 4938 3382 4941
rect 3682 4938 3686 4941
rect 3690 4938 3694 4941
rect 4130 4938 4137 4941
rect 182 4932 185 4938
rect 782 4932 785 4938
rect 106 4928 137 4931
rect 186 4928 206 4931
rect 210 4928 214 4931
rect 234 4928 342 4931
rect 418 4928 486 4931
rect 522 4928 534 4931
rect 538 4928 542 4931
rect 738 4928 758 4931
rect 842 4928 929 4931
rect 134 4922 137 4928
rect 170 4918 190 4921
rect 194 4918 350 4921
rect 358 4921 361 4928
rect 606 4922 609 4928
rect 926 4922 929 4928
rect 986 4928 1054 4931
rect 1226 4928 1254 4931
rect 1258 4928 1270 4931
rect 1378 4928 1430 4931
rect 1486 4931 1489 4938
rect 1486 4928 1614 4931
rect 1866 4928 1902 4931
rect 2162 4928 2206 4931
rect 2214 4931 2217 4938
rect 2214 4928 2254 4931
rect 2266 4928 2486 4931
rect 2802 4928 2881 4931
rect 2966 4931 2969 4938
rect 4134 4932 4137 4938
rect 4210 4938 4430 4941
rect 4742 4941 4745 4948
rect 4822 4941 4825 4948
rect 4742 4938 4825 4941
rect 4866 4938 4910 4941
rect 4914 4938 4966 4941
rect 5018 4938 5078 4941
rect 5130 4938 5153 4941
rect 4190 4932 4193 4938
rect 5150 4932 5153 4938
rect 2946 4928 2969 4931
rect 3114 4928 3278 4931
rect 3706 4928 3822 4931
rect 3826 4928 3846 4931
rect 4458 4928 4486 4931
rect 4490 4928 4694 4931
rect 5018 4928 5094 4931
rect 934 4922 937 4928
rect 2878 4922 2881 4928
rect 354 4918 361 4921
rect 378 4918 470 4921
rect 650 4918 670 4921
rect 722 4918 782 4921
rect 1082 4918 1198 4921
rect 1858 4918 1870 4921
rect 2034 4918 2054 4921
rect 2058 4918 2086 4921
rect 2098 4918 2158 4921
rect 2162 4918 2406 4921
rect 2426 4918 2598 4921
rect 2674 4918 2750 4921
rect 3570 4918 3582 4921
rect 3586 4918 3622 4921
rect 3658 4918 3758 4921
rect 3778 4918 3822 4921
rect 4050 4918 4054 4921
rect 4138 4918 4142 4921
rect 4162 4918 4182 4921
rect 4186 4918 4190 4921
rect 4374 4921 4377 4928
rect 5006 4922 5009 4928
rect 4250 4918 4377 4921
rect 4682 4918 4862 4921
rect 4866 4918 4894 4921
rect 5026 4918 5030 4921
rect 5090 4918 5174 4921
rect 5230 4912 5233 4918
rect 130 4908 430 4911
rect 466 4908 566 4911
rect 706 4908 750 4911
rect 754 4908 766 4911
rect 1810 4908 1862 4911
rect 3146 4908 3590 4911
rect 3978 4908 4006 4911
rect 4290 4908 4310 4911
rect 4650 4908 4838 4911
rect 848 4903 850 4907
rect 854 4903 857 4907
rect 862 4903 864 4907
rect 1872 4903 1874 4907
rect 1878 4903 1881 4907
rect 1886 4903 1888 4907
rect 2102 4902 2105 4908
rect 2888 4903 2890 4907
rect 2894 4903 2897 4907
rect 2902 4903 2904 4907
rect 3920 4903 3922 4907
rect 3926 4903 3929 4907
rect 3934 4903 3936 4907
rect 4936 4903 4938 4907
rect 4942 4903 4945 4907
rect 4950 4903 4952 4907
rect 74 4898 190 4901
rect 250 4898 390 4901
rect 466 4898 582 4901
rect 874 4898 950 4901
rect 954 4898 1318 4901
rect 1322 4898 1342 4901
rect 1410 4898 1422 4901
rect 2634 4898 2878 4901
rect 3074 4898 3414 4901
rect 4242 4898 4294 4901
rect 4298 4898 4446 4901
rect 4450 4898 4478 4901
rect 4482 4898 4526 4901
rect 4546 4898 4678 4901
rect 5046 4892 5049 4898
rect 170 4888 182 4891
rect 314 4888 798 4891
rect 802 4888 1006 4891
rect 1154 4888 1182 4891
rect 1186 4888 1350 4891
rect 1354 4888 1486 4891
rect 1730 4888 1742 4891
rect 1746 4888 1910 4891
rect 2578 4888 2582 4891
rect 2854 4888 2966 4891
rect 2986 4888 3022 4891
rect 3138 4888 3233 4891
rect 3442 4888 3598 4891
rect 3618 4888 3758 4891
rect 3762 4888 3934 4891
rect 3938 4888 4094 4891
rect 4278 4888 4286 4891
rect 4290 4888 4294 4891
rect 4966 4888 4974 4891
rect 4978 4888 5022 4891
rect 5170 4888 5190 4891
rect 114 4878 302 4881
rect 346 4878 374 4881
rect 394 4878 406 4881
rect 434 4878 454 4881
rect 546 4878 550 4881
rect 586 4878 646 4881
rect 650 4878 694 4881
rect 714 4878 822 4881
rect 930 4878 982 4881
rect 986 4878 1046 4881
rect 1050 4878 1054 4881
rect 1218 4878 1230 4881
rect 1418 4878 1470 4881
rect 1986 4878 2326 4881
rect 2414 4881 2417 4888
rect 2854 4882 2857 4888
rect 3230 4882 3233 4888
rect 2414 4878 2454 4881
rect 2562 4878 2574 4881
rect 2578 4878 2646 4881
rect 2922 4878 3022 4881
rect 3234 4878 3430 4881
rect 3506 4878 3550 4881
rect 3554 4878 3622 4881
rect 3674 4878 3734 4881
rect 4102 4881 4105 4888
rect 5030 4882 5033 4888
rect 4102 4878 4118 4881
rect 4210 4878 4230 4881
rect 4274 4878 4286 4881
rect 4290 4878 4326 4881
rect 4882 4878 4974 4881
rect 5170 4878 5246 4881
rect 5258 4878 5262 4881
rect 122 4868 126 4871
rect 130 4868 254 4871
rect 314 4868 422 4871
rect 426 4868 478 4871
rect 482 4868 950 4871
rect 1026 4868 1086 4871
rect 1090 4868 1174 4871
rect 1178 4868 1182 4871
rect 1242 4868 1254 4871
rect 1386 4870 1494 4871
rect 1386 4868 1438 4870
rect 1442 4868 1494 4870
rect 1666 4868 1745 4871
rect 2074 4868 2166 4871
rect 2410 4868 2430 4871
rect 2594 4868 2726 4871
rect 2962 4868 2982 4871
rect 2986 4868 3030 4871
rect 3034 4868 3054 4871
rect 3218 4868 3254 4871
rect 3290 4868 3302 4871
rect 3530 4868 3550 4871
rect 3554 4868 3806 4871
rect 4002 4868 4022 4871
rect 4058 4868 4110 4871
rect 4274 4868 4302 4871
rect 4306 4868 4366 4871
rect 4370 4868 4406 4871
rect 4498 4868 4566 4871
rect 4570 4868 4577 4871
rect 4730 4868 4790 4871
rect 4810 4868 5006 4871
rect 5066 4868 5070 4871
rect 5082 4868 5110 4871
rect 5250 4868 5254 4871
rect 1742 4862 1745 4868
rect 154 4858 310 4861
rect 362 4858 510 4861
rect 530 4858 606 4861
rect 626 4858 638 4861
rect 706 4858 774 4861
rect 794 4858 798 4861
rect 810 4858 862 4861
rect 874 4858 878 4861
rect 898 4858 950 4861
rect 1010 4858 1078 4861
rect 1082 4858 1086 4861
rect 1178 4858 1230 4861
rect 1458 4858 1462 4861
rect 1506 4858 1574 4861
rect 1778 4858 1862 4861
rect 1890 4858 1982 4861
rect 1994 4858 2022 4861
rect 2026 4858 2142 4861
rect 2146 4858 2182 4861
rect 2194 4858 2225 4861
rect 2442 4858 2478 4861
rect 2502 4861 2505 4868
rect 2502 4858 2582 4861
rect 2594 4858 2606 4861
rect 2794 4858 2862 4861
rect 2902 4858 3078 4861
rect 3166 4861 3169 4868
rect 3122 4858 3169 4861
rect 3250 4858 3278 4861
rect 3402 4858 3630 4861
rect 3682 4858 3686 4861
rect 3858 4858 3958 4861
rect 4018 4858 4086 4861
rect 4090 4858 4118 4861
rect 4138 4858 4142 4861
rect 4214 4861 4217 4868
rect 4230 4861 4233 4868
rect 4214 4858 4233 4861
rect 4302 4858 4310 4861
rect 4314 4858 4374 4861
rect 4570 4858 4582 4861
rect 5014 4861 5017 4868
rect 4690 4858 5017 4861
rect 5090 4858 5134 4861
rect 5242 4858 5278 4861
rect 38 4852 41 4858
rect 2222 4852 2225 4858
rect 2902 4852 2905 4858
rect 4606 4852 4609 4858
rect 138 4848 158 4851
rect 170 4848 174 4851
rect 322 4848 374 4851
rect 410 4848 486 4851
rect 506 4848 638 4851
rect 642 4848 694 4851
rect 746 4848 806 4851
rect 850 4848 1078 4851
rect 1106 4848 1134 4851
rect 1138 4848 1158 4851
rect 1162 4848 1185 4851
rect 2146 4848 2158 4851
rect 2330 4848 2441 4851
rect 2522 4848 2542 4851
rect 2562 4848 2622 4851
rect 3258 4848 3262 4851
rect 3578 4848 3582 4851
rect 3602 4848 3617 4851
rect 154 4838 214 4841
rect 254 4841 257 4848
rect 254 4838 278 4841
rect 338 4838 342 4841
rect 398 4841 401 4848
rect 1182 4842 1185 4848
rect 2438 4842 2441 4848
rect 398 4838 446 4841
rect 522 4838 566 4841
rect 578 4838 702 4841
rect 738 4838 886 4841
rect 978 4838 1030 4841
rect 2634 4838 2926 4841
rect 2930 4838 2934 4841
rect 2954 4838 3262 4841
rect 3350 4841 3353 4848
rect 3614 4842 3617 4848
rect 3654 4848 3673 4851
rect 3722 4848 3742 4851
rect 3746 4848 3838 4851
rect 4026 4848 4046 4851
rect 4082 4848 4094 4851
rect 4106 4848 4190 4851
rect 4218 4848 4222 4851
rect 4226 4848 4270 4851
rect 4634 4848 4694 4851
rect 4698 4848 4894 4851
rect 4978 4848 5046 4851
rect 5074 4848 5094 4851
rect 5258 4848 5262 4851
rect 5334 4851 5338 4852
rect 5306 4848 5338 4851
rect 3654 4842 3657 4848
rect 3670 4842 3673 4848
rect 3350 4838 3478 4841
rect 3506 4838 3606 4841
rect 3914 4838 3950 4841
rect 3994 4838 4318 4841
rect 4322 4838 4406 4841
rect 4538 4838 4686 4841
rect 5058 4838 5078 4841
rect 5226 4838 5270 4841
rect 106 4828 118 4831
rect 574 4831 577 4838
rect 122 4828 577 4831
rect 658 4828 766 4831
rect 778 4828 838 4831
rect 866 4828 1038 4831
rect 1098 4828 1126 4831
rect 1130 4828 1166 4831
rect 1170 4828 1246 4831
rect 2682 4828 3270 4831
rect 3314 4828 3326 4831
rect 3330 4828 3750 4831
rect 3754 4828 3926 4831
rect 3930 4828 4126 4831
rect 114 4818 214 4821
rect 218 4818 246 4821
rect 370 4818 438 4821
rect 554 4818 558 4821
rect 618 4818 670 4821
rect 674 4818 878 4821
rect 1282 4818 1430 4821
rect 1434 4818 1654 4821
rect 2354 4818 2918 4821
rect 2922 4818 2926 4821
rect 3426 4818 3798 4821
rect 3802 4818 3974 4821
rect 3978 4818 4182 4821
rect 4186 4818 4214 4821
rect 4426 4818 4726 4821
rect 4994 4818 5278 4821
rect 5286 4812 5289 4818
rect 418 4808 526 4811
rect 818 4808 1118 4811
rect 2210 4808 2262 4811
rect 2266 4808 2334 4811
rect 2418 4808 2438 4811
rect 2514 4808 2566 4811
rect 3626 4808 3662 4811
rect 3666 4808 3678 4811
rect 4042 4808 4174 4811
rect 5002 4808 5006 4811
rect 5018 4808 5150 4811
rect 328 4803 330 4807
rect 334 4803 337 4807
rect 342 4803 344 4807
rect 1352 4803 1354 4807
rect 1358 4803 1361 4807
rect 1366 4803 1368 4807
rect 2384 4803 2386 4807
rect 2390 4803 2393 4807
rect 2398 4803 2400 4807
rect 3400 4803 3402 4807
rect 3406 4803 3409 4807
rect 3414 4803 3416 4807
rect 4424 4803 4426 4807
rect 4430 4803 4433 4807
rect 4438 4803 4440 4807
rect 402 4798 590 4801
rect 594 4798 606 4801
rect 610 4798 958 4801
rect 1658 4798 2174 4801
rect 2186 4798 2190 4801
rect 2218 4798 2222 4801
rect 3530 4798 3582 4801
rect 3794 4798 3806 4801
rect 3986 4798 4150 4801
rect 4154 4798 4334 4801
rect 4338 4798 4398 4801
rect 4554 4798 4558 4801
rect 4586 4798 5054 4801
rect 338 4788 582 4791
rect 646 4788 662 4791
rect 666 4788 710 4791
rect 746 4788 926 4791
rect 954 4788 1126 4791
rect 1362 4788 1406 4791
rect 1842 4788 1870 4791
rect 1874 4788 2126 4791
rect 2426 4788 2462 4791
rect 2834 4788 2958 4791
rect 3306 4788 3686 4791
rect 3738 4788 4038 4791
rect 4082 4788 4126 4791
rect 4138 4788 4166 4791
rect 4170 4788 4454 4791
rect 4458 4788 4502 4791
rect 4506 4788 4630 4791
rect 4658 4788 4686 4791
rect 4978 4788 5238 4791
rect 5266 4788 5302 4791
rect 606 4782 609 4788
rect 210 4778 278 4781
rect 434 4778 438 4781
rect 490 4778 494 4781
rect 554 4778 566 4781
rect 622 4781 625 4788
rect 646 4782 649 4788
rect 2158 4782 2161 4788
rect 622 4778 638 4781
rect 798 4778 806 4781
rect 810 4778 953 4781
rect 962 4778 982 4781
rect 986 4778 1158 4781
rect 1186 4778 1366 4781
rect 1522 4778 1846 4781
rect 2122 4778 2158 4781
rect 2218 4778 2358 4781
rect 2362 4778 2430 4781
rect 2882 4778 2894 4781
rect 2898 4778 3150 4781
rect 3154 4778 3430 4781
rect 3754 4778 3990 4781
rect 4002 4778 4046 4781
rect 4090 4778 4710 4781
rect 4714 4778 4750 4781
rect 4754 4778 4798 4781
rect 5010 4778 5134 4781
rect 462 4772 465 4778
rect 66 4768 126 4771
rect 194 4768 222 4771
rect 234 4768 318 4771
rect 394 4768 422 4771
rect 426 4768 438 4771
rect 586 4768 662 4771
rect 666 4768 817 4771
rect 834 4768 918 4771
rect 950 4771 953 4778
rect 1854 4772 1857 4778
rect 950 4768 1014 4771
rect 1162 4768 1238 4771
rect 1338 4768 1342 4771
rect 1394 4768 1606 4771
rect 1970 4768 2190 4771
rect 2198 4768 2254 4771
rect 2986 4768 3182 4771
rect 3386 4768 3422 4771
rect 3706 4768 3814 4771
rect 3842 4768 3950 4771
rect 4002 4768 4182 4771
rect 4674 4768 4686 4771
rect 4738 4768 4998 4771
rect 5010 4768 5046 4771
rect 5082 4768 5102 4771
rect 814 4762 817 4768
rect 1038 4762 1041 4768
rect 90 4758 142 4761
rect 146 4758 286 4761
rect 290 4758 470 4761
rect 474 4758 550 4761
rect 554 4758 662 4761
rect 738 4758 750 4761
rect 858 4758 998 4761
rect 1106 4758 1134 4761
rect 1202 4758 1278 4761
rect 1314 4758 1574 4761
rect 1858 4758 1878 4761
rect 1970 4758 2046 4761
rect 2098 4758 2102 4761
rect 2114 4758 2134 4761
rect 2198 4761 2201 4768
rect 2138 4758 2201 4761
rect 2254 4761 2257 4768
rect 2254 4758 2294 4761
rect 2298 4758 2422 4761
rect 2642 4758 2654 4761
rect 3058 4758 3094 4761
rect 3778 4758 3846 4761
rect 3874 4758 3910 4761
rect 3914 4758 3982 4761
rect 3986 4758 4070 4761
rect 4414 4761 4417 4768
rect 4414 4758 4446 4761
rect 4450 4758 4494 4761
rect 4522 4758 4534 4761
rect 4550 4758 4638 4761
rect 4746 4758 4806 4761
rect 5190 4761 5193 4768
rect 5034 4758 5193 4761
rect 1310 4752 1313 4758
rect 50 4748 102 4751
rect 106 4748 126 4751
rect 130 4748 158 4751
rect 190 4748 198 4751
rect 202 4748 414 4751
rect 426 4748 430 4751
rect 546 4748 846 4751
rect 858 4748 990 4751
rect 1042 4748 1094 4751
rect 1114 4748 1142 4751
rect 1174 4748 1209 4751
rect 1250 4748 1254 4751
rect 1274 4748 1302 4751
rect 1490 4748 1526 4751
rect 1586 4748 1614 4751
rect 1618 4748 1646 4751
rect 1690 4748 1710 4751
rect 1730 4748 1798 4751
rect 1890 4748 2158 4751
rect 2162 4748 2206 4751
rect 2274 4748 2350 4751
rect 2490 4748 2534 4751
rect 2610 4748 2614 4751
rect 2634 4748 2710 4751
rect 2802 4748 2854 4751
rect 2926 4751 2929 4758
rect 2882 4748 2929 4751
rect 3058 4748 3062 4751
rect 3290 4748 3310 4751
rect 90 4738 142 4741
rect 146 4738 150 4741
rect 234 4738 262 4741
rect 422 4741 425 4748
rect 1174 4742 1177 4748
rect 1206 4742 1209 4748
rect 1446 4742 1449 4748
rect 1566 4742 1569 4748
rect 394 4738 425 4741
rect 490 4738 502 4741
rect 522 4738 561 4741
rect 578 4738 598 4741
rect 674 4738 742 4741
rect 802 4738 814 4741
rect 834 4738 854 4741
rect 906 4738 918 4741
rect 922 4738 1110 4741
rect 1138 4738 1142 4741
rect 1270 4738 1382 4741
rect 1582 4741 1585 4748
rect 1570 4738 1585 4741
rect 1602 4738 1670 4741
rect 1830 4741 1833 4748
rect 1830 4738 1894 4741
rect 1946 4738 2022 4741
rect 2074 4738 2150 4741
rect 2186 4738 2278 4741
rect 2454 4741 2457 4748
rect 3414 4751 3417 4758
rect 3378 4748 3417 4751
rect 3638 4751 3641 4758
rect 4550 4752 4553 4758
rect 3546 4748 3641 4751
rect 3706 4748 3878 4751
rect 4154 4748 4161 4751
rect 4194 4748 4286 4751
rect 4578 4748 4614 4751
rect 4650 4748 4681 4751
rect 4706 4748 4782 4751
rect 5042 4748 5046 4751
rect 5162 4748 5238 4751
rect 2362 4738 2457 4741
rect 2482 4738 2558 4741
rect 2586 4738 2606 4741
rect 2610 4738 2638 4741
rect 2874 4738 2902 4741
rect 2994 4738 3070 4741
rect 3270 4738 3358 4741
rect 3494 4741 3497 4748
rect 3450 4738 3497 4741
rect 3662 4741 3665 4748
rect 3662 4738 3766 4741
rect 3770 4738 3854 4741
rect 4006 4741 4009 4748
rect 3962 4738 4009 4741
rect 4030 4742 4033 4748
rect 4158 4742 4161 4748
rect 4050 4738 4078 4741
rect 4082 4738 4094 4741
rect 4318 4741 4321 4748
rect 4334 4741 4337 4748
rect 4574 4742 4577 4748
rect 4678 4742 4681 4748
rect 4318 4738 4358 4741
rect 4362 4738 4454 4741
rect 4770 4738 4774 4741
rect 4914 4738 5070 4741
rect 5138 4738 5166 4741
rect 214 4732 217 4738
rect 558 4732 561 4738
rect 10 4728 158 4731
rect 594 4728 622 4731
rect 626 4728 630 4731
rect 738 4728 742 4731
rect 754 4728 854 4731
rect 890 4728 902 4731
rect 922 4728 974 4731
rect 978 4728 1054 4731
rect 1074 4728 1102 4731
rect 1106 4728 1110 4731
rect 1158 4731 1161 4738
rect 1270 4732 1273 4738
rect 2870 4732 2873 4738
rect 3270 4732 3273 4738
rect 1138 4728 1161 4731
rect 1178 4728 1182 4731
rect 1194 4728 1230 4731
rect 1306 4728 1342 4731
rect 1466 4728 1566 4731
rect 1618 4728 1641 4731
rect 1802 4728 1886 4731
rect 2186 4728 2422 4731
rect 2438 4728 2454 4731
rect 2538 4728 2598 4731
rect 2602 4728 2606 4731
rect 2858 4728 2862 4731
rect 2890 4728 2894 4731
rect 2978 4728 3150 4731
rect 3570 4728 3734 4731
rect 3738 4728 3742 4731
rect 4002 4728 4134 4731
rect 4138 4728 4150 4731
rect 4450 4728 4470 4731
rect 4490 4728 4518 4731
rect 4522 4728 4582 4731
rect 4682 4728 4694 4731
rect 4698 4728 4966 4731
rect 4994 4728 5118 4731
rect 5122 4728 5222 4731
rect 1606 4722 1609 4728
rect 1638 4722 1641 4728
rect 34 4718 62 4721
rect 66 4718 86 4721
rect 122 4718 142 4721
rect 146 4718 238 4721
rect 442 4718 646 4721
rect 650 4718 726 4721
rect 794 4718 822 4721
rect 866 4718 942 4721
rect 1018 4718 1022 4721
rect 1154 4718 1222 4721
rect 1650 4718 1758 4721
rect 2430 4721 2433 4728
rect 2338 4718 2433 4721
rect 2438 4722 2441 4728
rect 2850 4718 2886 4721
rect 3154 4718 3238 4721
rect 3354 4718 3358 4721
rect 3990 4721 3993 4728
rect 3610 4718 3993 4721
rect 4138 4718 4206 4721
rect 4218 4718 4230 4721
rect 4482 4718 4526 4721
rect 4578 4718 4630 4721
rect 4730 4718 4742 4721
rect 4746 4718 4774 4721
rect 4922 4718 4990 4721
rect 5050 4718 5054 4721
rect 5178 4718 5182 4721
rect 2006 4712 2009 4718
rect 2662 4712 2665 4718
rect 2846 4712 2849 4718
rect 58 4708 222 4711
rect 466 4708 638 4711
rect 698 4708 774 4711
rect 906 4708 934 4711
rect 1050 4708 1054 4711
rect 1058 4708 1246 4711
rect 1634 4708 1726 4711
rect 2010 4708 2118 4711
rect 2394 4708 2438 4711
rect 2442 4708 2478 4711
rect 3026 4708 3190 4711
rect 3194 4708 3206 4711
rect 3210 4708 3489 4711
rect 3506 4708 3526 4711
rect 3554 4708 3574 4711
rect 3674 4708 3678 4711
rect 3714 4708 3774 4711
rect 3834 4708 3838 4711
rect 4066 4708 4238 4711
rect 4242 4708 4342 4711
rect 4410 4708 4758 4711
rect 4762 4708 4926 4711
rect 5146 4708 5174 4711
rect 38 4702 41 4708
rect 848 4703 850 4707
rect 854 4703 857 4707
rect 862 4703 864 4707
rect 1872 4703 1874 4707
rect 1878 4703 1881 4707
rect 1886 4703 1888 4707
rect 2888 4703 2890 4707
rect 2894 4703 2897 4707
rect 2902 4703 2904 4707
rect 3486 4702 3489 4708
rect 3920 4703 3922 4707
rect 3926 4703 3929 4707
rect 3934 4703 3936 4707
rect 4936 4703 4938 4707
rect 4942 4703 4945 4707
rect 4950 4703 4952 4707
rect 42 4698 246 4701
rect 250 4698 318 4701
rect 498 4698 606 4701
rect 666 4698 726 4701
rect 730 4698 790 4701
rect 922 4698 926 4701
rect 938 4698 950 4701
rect 994 4698 1006 4701
rect 1010 4698 1086 4701
rect 1090 4698 1102 4701
rect 1106 4698 1126 4701
rect 1138 4698 1169 4701
rect 1242 4698 1286 4701
rect 1290 4698 1310 4701
rect 1314 4698 1438 4701
rect 1562 4698 1646 4701
rect 1650 4698 1654 4701
rect 1682 4698 1742 4701
rect 1954 4698 2078 4701
rect 2290 4698 2374 4701
rect 3106 4698 3438 4701
rect 3490 4698 3902 4701
rect 4034 4698 4414 4701
rect 4418 4698 4430 4701
rect 4514 4698 4638 4701
rect 4682 4698 4710 4701
rect 5002 4698 5022 4701
rect 5026 4698 5038 4701
rect 5090 4698 5102 4701
rect 130 4688 134 4691
rect 370 4688 526 4691
rect 538 4688 598 4691
rect 934 4688 942 4691
rect 946 4688 966 4691
rect 1082 4688 1158 4691
rect 1166 4691 1169 4698
rect 1166 4688 1270 4691
rect 1370 4688 1462 4691
rect 1474 4688 1686 4691
rect 1802 4688 1886 4691
rect 2270 4688 2310 4691
rect 2434 4688 2462 4691
rect 2562 4688 2654 4691
rect 2938 4688 3094 4691
rect 3114 4688 3150 4691
rect 3162 4688 3302 4691
rect 3306 4688 3342 4691
rect 3402 4688 3641 4691
rect 3746 4688 3798 4691
rect 3890 4688 4070 4691
rect 4250 4688 4254 4691
rect 4290 4688 4366 4691
rect 4370 4688 4414 4691
rect 4538 4688 4622 4691
rect 4690 4688 4718 4691
rect 4858 4688 4902 4691
rect 4930 4688 5158 4691
rect 5162 4688 5166 4691
rect 210 4678 326 4681
rect 610 4678 734 4681
rect 822 4681 825 4688
rect 822 4678 870 4681
rect 886 4681 889 4688
rect 1342 4682 1345 4688
rect 2270 4682 2273 4688
rect 3638 4682 3641 4688
rect 886 4678 950 4681
rect 1002 4678 1134 4681
rect 1186 4678 1190 4681
rect 1194 4678 1198 4681
rect 1786 4678 2086 4681
rect 2538 4678 2638 4681
rect 2866 4678 2902 4681
rect 2914 4678 2926 4681
rect 3234 4678 3366 4681
rect 3370 4678 3422 4681
rect 3426 4678 3462 4681
rect 3466 4678 3566 4681
rect 3570 4678 3590 4681
rect 3866 4678 3910 4681
rect 4126 4681 4129 4688
rect 4126 4678 4206 4681
rect 4226 4678 4230 4681
rect 4570 4678 4654 4681
rect 4986 4678 5022 4681
rect 50 4668 102 4671
rect 122 4668 126 4671
rect 202 4668 206 4671
rect 298 4668 342 4671
rect 502 4671 505 4678
rect 370 4668 505 4671
rect 618 4668 638 4671
rect 674 4668 734 4671
rect 738 4668 758 4671
rect 762 4668 822 4671
rect 922 4668 1006 4671
rect 1142 4671 1145 4678
rect 1010 4668 1145 4671
rect 1246 4671 1249 4678
rect 1534 4672 1537 4678
rect 1226 4668 1249 4671
rect 1266 4668 1318 4671
rect 1410 4668 1422 4671
rect 1602 4668 1662 4671
rect 1762 4668 1782 4671
rect 2002 4668 2014 4671
rect 2058 4668 2110 4671
rect 2294 4671 2297 4678
rect 2218 4668 2297 4671
rect 2426 4668 2462 4671
rect 2490 4668 2590 4671
rect 2650 4668 2705 4671
rect 2754 4668 2870 4671
rect 2930 4668 3118 4671
rect 3230 4671 3233 4678
rect 3154 4668 3254 4671
rect 3322 4668 3350 4671
rect 3378 4668 3382 4671
rect 3682 4668 3758 4671
rect 3866 4668 3966 4671
rect 3994 4668 4094 4671
rect 4382 4671 4385 4678
rect 4382 4668 4478 4671
rect 4550 4671 4553 4678
rect 4522 4668 4553 4671
rect 4650 4668 4758 4671
rect 5046 4671 5049 4678
rect 4970 4668 5086 4671
rect 5202 4668 5246 4671
rect 98 4658 198 4661
rect 282 4658 422 4661
rect 426 4658 486 4661
rect 546 4658 606 4661
rect 634 4658 654 4661
rect 658 4658 694 4661
rect 746 4658 750 4661
rect 834 4658 838 4661
rect 874 4658 934 4661
rect 1050 4658 1078 4661
rect 1082 4658 1094 4661
rect 1106 4658 1198 4661
rect 1314 4658 1318 4661
rect 1402 4658 1406 4661
rect 1554 4659 1574 4661
rect 1554 4658 1577 4659
rect 1594 4659 1686 4661
rect 2702 4662 2705 4668
rect 3270 4662 3273 4668
rect 1594 4658 1689 4659
rect 1778 4658 1833 4661
rect 1850 4658 2126 4661
rect 2210 4658 2526 4661
rect 2530 4658 2582 4661
rect 2738 4658 2814 4661
rect 2858 4658 2934 4661
rect 3002 4658 3070 4661
rect 3170 4658 3190 4661
rect 3250 4658 3270 4661
rect 3438 4661 3441 4668
rect 3282 4658 3441 4661
rect 3634 4658 3654 4661
rect 3658 4658 3753 4661
rect 3778 4658 3814 4661
rect 3818 4658 3870 4661
rect 4018 4658 4030 4661
rect 4146 4658 4350 4661
rect 4354 4658 4390 4661
rect 4394 4658 4462 4661
rect 4466 4658 4526 4661
rect 4554 4658 4646 4661
rect 4666 4658 4670 4661
rect 4674 4658 4710 4661
rect 4714 4658 4774 4661
rect 4778 4658 4862 4661
rect 4866 4658 4894 4661
rect 5066 4658 5102 4661
rect 5106 4658 5134 4661
rect 278 4652 281 4658
rect 218 4648 222 4651
rect 226 4648 254 4651
rect 330 4648 334 4651
rect 346 4648 406 4651
rect 410 4648 478 4651
rect 482 4648 590 4651
rect 718 4651 721 4658
rect 1830 4652 1833 4658
rect 2006 4652 2009 4658
rect 3750 4652 3753 4658
rect 5142 4652 5145 4658
rect 602 4648 774 4651
rect 782 4648 982 4651
rect 1042 4648 1102 4651
rect 1130 4648 1158 4651
rect 1250 4648 1326 4651
rect 1714 4648 1814 4651
rect 2050 4648 2054 4651
rect 2290 4648 2326 4651
rect 2330 4648 2494 4651
rect 2498 4648 2518 4651
rect 2578 4648 2622 4651
rect 2850 4648 3054 4651
rect 3058 4648 3070 4651
rect 3090 4648 3198 4651
rect 3330 4648 3382 4651
rect 3466 4648 3486 4651
rect 3498 4648 3550 4651
rect 3554 4648 3742 4651
rect 3794 4648 3990 4651
rect 4082 4648 4278 4651
rect 4474 4648 4566 4651
rect 4674 4648 4694 4651
rect 4706 4648 4782 4651
rect 4890 4648 4982 4651
rect 5042 4648 5078 4651
rect 186 4638 198 4641
rect 218 4638 222 4641
rect 234 4638 398 4641
rect 402 4638 409 4641
rect 418 4638 486 4641
rect 490 4638 622 4641
rect 782 4641 785 4648
rect 690 4638 785 4641
rect 826 4638 846 4641
rect 982 4641 985 4648
rect 982 4638 1062 4641
rect 1234 4638 1302 4641
rect 1306 4638 1334 4641
rect 1370 4638 1406 4641
rect 1410 4638 1438 4641
rect 1778 4638 2094 4641
rect 2170 4638 2278 4641
rect 2370 4638 2518 4641
rect 3082 4638 3110 4641
rect 3114 4638 3230 4641
rect 3362 4638 3406 4641
rect 3634 4638 3638 4641
rect 3690 4638 3814 4641
rect 4030 4641 4033 4648
rect 4030 4638 4110 4641
rect 4906 4638 5022 4641
rect 5026 4638 5054 4641
rect 5122 4638 5150 4641
rect 2846 4632 2849 4638
rect 154 4628 350 4631
rect 618 4628 662 4631
rect 666 4628 694 4631
rect 762 4628 854 4631
rect 858 4628 1017 4631
rect 1058 4628 1078 4631
rect 1274 4628 1414 4631
rect 1754 4628 2038 4631
rect 2074 4628 2742 4631
rect 3018 4628 3046 4631
rect 3234 4628 3726 4631
rect 3730 4628 3998 4631
rect 4402 4628 4478 4631
rect 162 4618 214 4621
rect 322 4618 342 4621
rect 362 4618 390 4621
rect 702 4621 705 4628
rect 1014 4622 1017 4628
rect 602 4618 766 4621
rect 826 4618 934 4621
rect 1026 4618 1310 4621
rect 1322 4618 1366 4621
rect 2178 4618 2590 4621
rect 2802 4618 3342 4621
rect 3390 4618 3502 4621
rect 3730 4618 3782 4621
rect 4066 4618 4086 4621
rect 4418 4618 4846 4621
rect 4850 4618 5054 4621
rect 582 4612 585 4618
rect 1606 4612 1609 4618
rect 594 4608 622 4611
rect 698 4608 1030 4611
rect 1258 4608 1294 4611
rect 1898 4608 1974 4611
rect 2698 4608 2950 4611
rect 3390 4611 3393 4618
rect 3258 4608 3393 4611
rect 3826 4608 4142 4611
rect 4530 4608 4814 4611
rect 328 4603 330 4607
rect 334 4603 337 4607
rect 342 4603 344 4607
rect 1352 4603 1354 4607
rect 1358 4603 1361 4607
rect 1366 4603 1368 4607
rect 2384 4603 2386 4607
rect 2390 4603 2393 4607
rect 2398 4603 2400 4607
rect 3400 4603 3402 4607
rect 3406 4603 3409 4607
rect 3414 4603 3416 4607
rect 4424 4603 4426 4607
rect 4430 4603 4433 4607
rect 4438 4603 4440 4607
rect 98 4598 110 4601
rect 450 4598 526 4601
rect 538 4598 670 4601
rect 1746 4598 1758 4601
rect 2482 4598 2534 4601
rect 2674 4598 2702 4601
rect 3818 4598 4118 4601
rect 4506 4598 4574 4601
rect 4650 4598 4654 4601
rect 4978 4598 5094 4601
rect 114 4588 726 4591
rect 730 4588 894 4591
rect 978 4588 1118 4591
rect 1138 4588 1230 4591
rect 1250 4588 1305 4591
rect 1386 4588 1694 4591
rect 1698 4588 1745 4591
rect 2098 4588 2734 4591
rect 2746 4588 3478 4591
rect 3482 4588 3622 4591
rect 3842 4588 4038 4591
rect 4058 4588 4102 4591
rect 4106 4588 4526 4591
rect 4634 4588 4638 4591
rect 4650 4588 4654 4591
rect 4658 4588 4718 4591
rect 4922 4588 5145 4591
rect 5194 4588 5230 4591
rect 1302 4582 1305 4588
rect 1742 4582 1745 4588
rect 5142 4582 5145 4588
rect 138 4578 182 4581
rect 266 4578 358 4581
rect 362 4578 585 4581
rect 602 4578 654 4581
rect 658 4578 982 4581
rect 1050 4578 1110 4581
rect 1122 4578 1158 4581
rect 2234 4578 2366 4581
rect 2514 4578 2574 4581
rect 3266 4578 3494 4581
rect 3730 4578 3886 4581
rect 3946 4578 4134 4581
rect 4138 4578 4158 4581
rect 4234 4578 4606 4581
rect 4610 4578 4806 4581
rect 4810 4578 5046 4581
rect 582 4572 585 4578
rect 98 4568 134 4571
rect 150 4568 158 4571
rect 162 4568 174 4571
rect 234 4568 254 4571
rect 298 4568 414 4571
rect 474 4568 574 4571
rect 682 4568 694 4571
rect 1082 4568 1102 4571
rect 1106 4568 1182 4571
rect 1242 4568 1302 4571
rect 1474 4568 1478 4571
rect 2330 4568 2334 4571
rect 2362 4568 2510 4571
rect 2762 4568 2801 4571
rect 3034 4568 3118 4571
rect 3294 4568 3414 4571
rect 3418 4568 3518 4571
rect 3614 4568 3966 4571
rect 4122 4568 4166 4571
rect 4210 4568 4390 4571
rect 4402 4568 4854 4571
rect 5122 4568 5190 4571
rect 14 4561 17 4568
rect 14 4558 46 4561
rect 74 4558 94 4561
rect 98 4558 198 4561
rect 202 4558 318 4561
rect 450 4558 454 4561
rect 474 4558 566 4561
rect 570 4558 582 4561
rect 618 4558 702 4561
rect 742 4561 745 4568
rect 2358 4562 2361 4568
rect 2798 4562 2801 4568
rect 3294 4562 3297 4568
rect 3614 4562 3617 4568
rect 742 4558 798 4561
rect 802 4558 806 4561
rect 930 4558 950 4561
rect 954 4558 1038 4561
rect 1146 4558 1150 4561
rect 1170 4558 1190 4561
rect 1198 4558 1206 4561
rect 1210 4558 1214 4561
rect 1314 4558 1462 4561
rect 1578 4558 1662 4561
rect 1698 4558 1766 4561
rect 1950 4558 2038 4561
rect 2106 4558 2110 4561
rect 2138 4558 2190 4561
rect 2402 4558 2454 4561
rect 2594 4558 2766 4561
rect 2786 4558 2790 4561
rect 2802 4558 2870 4561
rect 3050 4558 3062 4561
rect 3218 4558 3222 4561
rect 3318 4558 3326 4561
rect 3330 4558 3358 4561
rect 3806 4558 3830 4561
rect 3874 4558 3878 4561
rect 4062 4561 4065 4568
rect 3890 4558 4065 4561
rect 4074 4558 4078 4561
rect 4146 4558 4150 4561
rect 4170 4558 4174 4561
rect 4218 4558 4222 4561
rect 4274 4558 4278 4561
rect 4418 4558 4430 4561
rect 4490 4558 4550 4561
rect 4626 4558 4662 4561
rect 4666 4558 4678 4561
rect 4682 4558 4686 4561
rect 4714 4558 4734 4561
rect 4842 4558 4974 4561
rect 4994 4558 4998 4561
rect 5162 4558 5190 4561
rect 5210 4558 5214 4561
rect 58 4548 86 4551
rect 170 4548 270 4551
rect 274 4548 494 4551
rect 498 4548 542 4551
rect 546 4548 638 4551
rect 642 4548 670 4551
rect 674 4548 710 4551
rect 786 4548 790 4551
rect 1118 4551 1121 4558
rect 1198 4551 1201 4558
rect 794 4548 1073 4551
rect 1118 4548 1201 4551
rect 1218 4548 1254 4551
rect 1274 4548 1350 4551
rect 1362 4548 1366 4551
rect 1470 4551 1473 4558
rect 1458 4548 1473 4551
rect 1502 4551 1505 4558
rect 1950 4552 1953 4558
rect 1502 4548 1614 4551
rect 1618 4548 1646 4551
rect 2122 4548 2190 4551
rect 2194 4548 2214 4551
rect 2218 4548 2414 4551
rect 2418 4548 2486 4551
rect 2490 4548 2782 4551
rect 2786 4548 2814 4551
rect 2818 4548 2838 4551
rect 2954 4548 2958 4551
rect 3034 4548 3153 4551
rect 3202 4548 3286 4551
rect 3290 4548 3321 4551
rect 1070 4542 1073 4548
rect 1958 4542 1961 4548
rect 50 4538 54 4541
rect 162 4538 174 4541
rect 234 4538 270 4541
rect 370 4538 374 4541
rect 386 4538 406 4541
rect 450 4538 462 4541
rect 514 4538 550 4541
rect 586 4538 598 4541
rect 818 4538 854 4541
rect 978 4538 1006 4541
rect 1010 4538 1014 4541
rect 1034 4538 1038 4541
rect 1074 4538 1134 4541
rect 1138 4538 1190 4541
rect 1210 4538 1238 4541
rect 1242 4538 1262 4541
rect 1266 4538 1382 4541
rect 1466 4538 1470 4541
rect 1498 4538 1542 4541
rect 1642 4538 1654 4541
rect 1778 4538 1918 4541
rect 1946 4538 1958 4541
rect 2194 4538 2222 4541
rect 2290 4538 2470 4541
rect 2474 4538 2678 4541
rect 2738 4538 2798 4541
rect 2818 4538 2822 4541
rect 3030 4541 3033 4548
rect 2986 4538 3033 4541
rect 3150 4542 3153 4548
rect 3318 4542 3321 4548
rect 3362 4548 3422 4551
rect 3478 4551 3481 4558
rect 3806 4552 3809 4558
rect 5150 4552 5153 4558
rect 3458 4548 3481 4551
rect 3530 4548 3534 4551
rect 3658 4548 3678 4551
rect 3682 4548 3710 4551
rect 3842 4548 3846 4551
rect 3882 4548 3942 4551
rect 3970 4548 4262 4551
rect 4410 4548 4446 4551
rect 4450 4548 4494 4551
rect 4506 4548 4510 4551
rect 4698 4548 4726 4551
rect 4762 4548 4830 4551
rect 4850 4548 4913 4551
rect 5082 4548 5134 4551
rect 3342 4542 3345 4548
rect 3734 4542 3737 4548
rect 4910 4542 4913 4548
rect 5182 4542 5185 4548
rect 3186 4538 3233 4541
rect 3434 4538 3446 4541
rect 3466 4538 3510 4541
rect 3522 4538 3526 4541
rect 3578 4538 3670 4541
rect 3906 4538 3918 4541
rect 3954 4538 3958 4541
rect 4106 4538 4110 4541
rect 4142 4538 4198 4541
rect 4202 4538 4238 4541
rect 4466 4538 4609 4541
rect 4658 4538 4702 4541
rect 4730 4538 4758 4541
rect 4778 4538 4790 4541
rect 4866 4538 4870 4541
rect 5002 4538 5025 4541
rect 5042 4538 5118 4541
rect 5146 4538 5166 4541
rect 26 4528 126 4531
rect 130 4528 206 4531
rect 210 4528 246 4531
rect 250 4528 278 4531
rect 430 4531 433 4538
rect 662 4532 665 4538
rect 2558 4532 2561 4538
rect 3230 4532 3233 4538
rect 410 4528 433 4531
rect 450 4528 518 4531
rect 546 4528 662 4531
rect 842 4528 918 4531
rect 922 4528 1038 4531
rect 1042 4528 1078 4531
rect 1130 4528 1174 4531
rect 1242 4528 1334 4531
rect 1338 4528 1358 4531
rect 1666 4528 1806 4531
rect 1810 4528 1950 4531
rect 2114 4528 2209 4531
rect 2266 4528 2334 4531
rect 2738 4528 2745 4531
rect 2866 4528 2870 4531
rect 2914 4528 3006 4531
rect 3010 4528 3134 4531
rect 3330 4528 3406 4531
rect 3466 4528 3470 4531
rect 3806 4531 3809 4538
rect 4142 4532 4145 4538
rect 4606 4532 4609 4538
rect 5022 4532 5025 4538
rect 3806 4528 3982 4531
rect 4002 4528 4110 4531
rect 4170 4528 4190 4531
rect 4210 4528 4246 4531
rect 4666 4528 4673 4531
rect 4706 4528 5014 4531
rect 5098 4528 5166 4531
rect 5194 4528 5214 4531
rect 82 4518 142 4521
rect 146 4518 230 4521
rect 466 4518 470 4521
rect 546 4518 590 4521
rect 694 4521 697 4528
rect 2206 4522 2209 4528
rect 2350 4522 2353 4528
rect 2742 4522 2745 4528
rect 3662 4522 3665 4528
rect 642 4518 697 4521
rect 786 4518 822 4521
rect 826 4518 902 4521
rect 906 4518 990 4521
rect 1050 4518 1166 4521
rect 1186 4518 1214 4521
rect 1218 4518 1270 4521
rect 1274 4518 1278 4521
rect 1282 4518 1342 4521
rect 1386 4518 1398 4521
rect 1402 4518 1406 4521
rect 1594 4518 1782 4521
rect 2378 4518 2398 4521
rect 3266 4518 3374 4521
rect 3458 4518 3494 4521
rect 3706 4518 3774 4521
rect 3778 4518 4054 4521
rect 4134 4521 4137 4528
rect 4670 4522 4673 4528
rect 4134 4518 4206 4521
rect 4242 4518 4350 4521
rect 4474 4518 4502 4521
rect 4730 4518 4750 4521
rect 4866 4518 4878 4521
rect 4882 4518 4974 4521
rect 4978 4518 5030 4521
rect 5138 4518 5254 4521
rect 2638 4512 2641 4518
rect 34 4508 110 4511
rect 218 4508 246 4511
rect 530 4508 598 4511
rect 642 4508 806 4511
rect 810 4508 830 4511
rect 1002 4508 1014 4511
rect 1018 4508 1158 4511
rect 1178 4508 1454 4511
rect 1514 4508 1542 4511
rect 1690 4508 1750 4511
rect 1842 4508 1862 4511
rect 2666 4508 2790 4511
rect 3034 4508 3102 4511
rect 3106 4508 3214 4511
rect 3218 4508 3398 4511
rect 3570 4508 3761 4511
rect 3770 4508 3878 4511
rect 3946 4508 4094 4511
rect 4298 4508 4318 4511
rect 4322 4508 4358 4511
rect 4690 4508 4734 4511
rect 4746 4508 4790 4511
rect 4986 4508 5006 4511
rect 5130 4508 5166 4511
rect 848 4503 850 4507
rect 854 4503 857 4507
rect 862 4503 864 4507
rect 1872 4503 1874 4507
rect 1878 4503 1881 4507
rect 1886 4503 1888 4507
rect 2888 4503 2890 4507
rect 2894 4503 2897 4507
rect 2902 4503 2904 4507
rect 370 4498 390 4501
rect 570 4498 590 4501
rect 634 4498 678 4501
rect 914 4498 934 4501
rect 938 4498 1174 4501
rect 1178 4498 1326 4501
rect 1330 4498 1438 4501
rect 1442 4498 1686 4501
rect 1898 4498 2022 4501
rect 2106 4498 2454 4501
rect 2618 4498 2686 4501
rect 2762 4498 2830 4501
rect 3098 4498 3166 4501
rect 3170 4498 3222 4501
rect 3226 4498 3270 4501
rect 3274 4498 3542 4501
rect 3690 4498 3694 4501
rect 3758 4501 3761 4508
rect 3920 4503 3922 4507
rect 3926 4503 3929 4507
rect 3934 4503 3936 4507
rect 4936 4503 4938 4507
rect 4942 4503 4945 4507
rect 4950 4503 4952 4507
rect 3758 4498 3846 4501
rect 3858 4498 3878 4501
rect 4098 4498 4350 4501
rect 4690 4498 4718 4501
rect 4722 4498 4790 4501
rect 4994 4498 4998 4501
rect 498 4488 574 4491
rect 578 4488 630 4491
rect 674 4488 678 4491
rect 802 4488 854 4491
rect 1130 4488 1225 4491
rect 1266 4488 1326 4491
rect 1362 4488 1390 4491
rect 1490 4488 1574 4491
rect 1578 4488 1782 4491
rect 2018 4488 2070 4491
rect 2162 4488 2726 4491
rect 2754 4488 2814 4491
rect 2826 4488 2846 4491
rect 2850 4488 2894 4491
rect 2946 4488 3006 4491
rect 3338 4488 3550 4491
rect 3586 4488 3670 4491
rect 3826 4488 3854 4491
rect 3866 4488 3934 4491
rect 3946 4488 4006 4491
rect 4290 4488 4398 4491
rect 4402 4488 4414 4491
rect 4418 4488 4462 4491
rect 4498 4488 4694 4491
rect 4858 4488 4902 4491
rect 4998 4488 5078 4491
rect 5114 4488 5126 4491
rect 5130 4488 5206 4491
rect 142 4482 145 4488
rect 1222 4482 1225 4488
rect 3718 4482 3721 4488
rect 4998 4482 5001 4488
rect 58 4478 142 4481
rect 170 4478 214 4481
rect 362 4478 390 4481
rect 442 4478 582 4481
rect 602 4478 806 4481
rect 978 4478 982 4481
rect 1278 4478 1286 4481
rect 1290 4478 1294 4481
rect 1314 4478 1342 4481
rect 1354 4478 1374 4481
rect 1618 4478 1662 4481
rect 1674 4478 1710 4481
rect 1714 4478 1718 4481
rect 1746 4478 1854 4481
rect 1922 4478 2238 4481
rect 2370 4478 2382 4481
rect 2690 4478 2742 4481
rect 2746 4478 2910 4481
rect 3102 4478 3110 4481
rect 3122 4478 3158 4481
rect 3162 4478 3246 4481
rect 3506 4478 3590 4481
rect 3594 4478 3686 4481
rect 3842 4478 3870 4481
rect 3946 4478 4166 4481
rect 4394 4478 4438 4481
rect 4482 4478 4534 4481
rect 4586 4478 4630 4481
rect 4818 4478 4942 4481
rect 4970 4478 4982 4481
rect 5066 4478 5102 4481
rect 5154 4478 5198 4481
rect 1070 4472 1073 4478
rect 66 4468 182 4471
rect 186 4468 262 4471
rect 298 4468 446 4471
rect 498 4468 502 4471
rect 554 4468 558 4471
rect 706 4468 710 4471
rect 714 4468 718 4471
rect 770 4468 798 4471
rect 834 4468 886 4471
rect 890 4468 894 4471
rect 946 4468 950 4471
rect 970 4468 982 4471
rect 1142 4471 1145 4478
rect 2406 4472 2409 4478
rect 3102 4472 3105 4478
rect 1078 4468 1145 4471
rect 1162 4468 1174 4471
rect 1250 4468 1286 4471
rect 1474 4468 1622 4471
rect 1626 4468 1654 4471
rect 1850 4468 2078 4471
rect 2106 4468 2190 4471
rect 2482 4468 2534 4471
rect 2602 4468 2702 4471
rect 2714 4468 2838 4471
rect 2842 4468 2854 4471
rect 2882 4468 2974 4471
rect 3026 4468 3078 4471
rect 3114 4468 3118 4471
rect 3154 4468 3174 4471
rect 3218 4468 3222 4471
rect 3382 4471 3385 4478
rect 3314 4468 3385 4471
rect 3418 4468 3438 4471
rect 3570 4468 3614 4471
rect 3730 4468 3734 4471
rect 3822 4468 3910 4471
rect 4098 4468 4102 4471
rect 4190 4468 4254 4471
rect 4514 4468 4574 4471
rect 4594 4468 4758 4471
rect 4762 4468 4894 4471
rect 4914 4468 4926 4471
rect 5018 4468 5118 4471
rect 5154 4468 5158 4471
rect 5186 4468 5254 4471
rect 106 4458 110 4461
rect 114 4458 166 4461
rect 234 4458 326 4461
rect 362 4458 401 4461
rect 410 4458 438 4461
rect 490 4458 518 4461
rect 522 4458 614 4461
rect 618 4458 654 4461
rect 706 4458 774 4461
rect 826 4458 862 4461
rect 938 4458 1030 4461
rect 1078 4461 1081 4468
rect 1158 4462 1161 4468
rect 1050 4458 1081 4461
rect 1106 4458 1118 4461
rect 1122 4458 1153 4461
rect 1226 4458 1254 4461
rect 1294 4461 1297 4468
rect 1846 4462 1849 4468
rect 3822 4462 3825 4468
rect 4190 4462 4193 4468
rect 1294 4458 1310 4461
rect 1314 4458 1414 4461
rect 1450 4458 1462 4461
rect 1634 4458 1742 4461
rect 1794 4458 1806 4461
rect 1834 4458 1846 4461
rect 2074 4458 2078 4461
rect 2098 4458 2126 4461
rect 2130 4458 2134 4461
rect 2226 4458 2342 4461
rect 2346 4458 2382 4461
rect 2570 4458 2630 4461
rect 2690 4458 2830 4461
rect 2874 4458 3062 4461
rect 3074 4458 3086 4461
rect 3122 4458 3126 4461
rect 3202 4458 3230 4461
rect 3546 4458 3566 4461
rect 3714 4458 3790 4461
rect 4026 4458 4030 4461
rect 4042 4458 4062 4461
rect 4094 4458 4161 4461
rect 4250 4458 4318 4461
rect 4498 4458 4518 4461
rect 4810 4458 4822 4461
rect 4858 4458 4862 4461
rect 4906 4458 5017 4461
rect 5122 4458 5166 4461
rect 5186 4458 5190 4461
rect 398 4452 401 4458
rect -26 4451 -22 4452
rect -26 4448 6 4451
rect 90 4448 118 4451
rect 122 4448 270 4451
rect 274 4448 310 4451
rect 474 4448 526 4451
rect 538 4448 566 4451
rect 578 4448 582 4451
rect 586 4448 638 4451
rect 714 4448 718 4451
rect 770 4448 814 4451
rect 874 4448 897 4451
rect 962 4448 998 4451
rect 1074 4448 1094 4451
rect 1150 4451 1153 4458
rect 1998 4452 2001 4458
rect 2598 4452 2601 4458
rect 1150 4448 1182 4451
rect 1202 4448 1214 4451
rect 1218 4448 1257 4451
rect 1290 4448 1342 4451
rect 1346 4448 1350 4451
rect 1386 4448 1462 4451
rect 1474 4448 1518 4451
rect 1570 4448 1582 4451
rect 1794 4448 1982 4451
rect 2018 4448 2022 4451
rect 2034 4448 2094 4451
rect 2306 4448 2526 4451
rect 2666 4448 2758 4451
rect 3058 4448 3062 4451
rect 3082 4448 3206 4451
rect 3258 4448 3350 4451
rect 3382 4451 3385 4458
rect 3838 4452 3841 4458
rect 4094 4452 4097 4458
rect 3362 4448 3385 4451
rect 3394 4448 3462 4451
rect 3570 4448 3726 4451
rect 3734 4448 3798 4451
rect 3894 4448 3974 4451
rect 4106 4448 4150 4451
rect 4158 4451 4161 4458
rect 4630 4452 4633 4458
rect 5014 4452 5017 4458
rect 4158 4448 4334 4451
rect 4634 4448 4654 4451
rect 4674 4448 4726 4451
rect 4730 4448 4830 4451
rect 5106 4448 5230 4451
rect 894 4442 897 4448
rect 1254 4442 1257 4448
rect 3222 4442 3225 4448
rect 3734 4442 3737 4448
rect 3894 4442 3897 4448
rect 10 4438 86 4441
rect 146 4438 681 4441
rect 690 4438 718 4441
rect 778 4438 830 4441
rect 834 4438 886 4441
rect 1090 4438 1102 4441
rect 1434 4438 1702 4441
rect 1706 4438 2086 4441
rect 2394 4438 2686 4441
rect 2698 4438 2814 4441
rect 3290 4438 3366 4441
rect 3370 4438 3390 4441
rect 3394 4438 3534 4441
rect 4010 4438 4014 4441
rect 4098 4438 4150 4441
rect 4186 4438 4198 4441
rect 4610 4438 4958 4441
rect 4986 4438 4998 4441
rect 5022 4441 5025 4448
rect 5002 4438 5025 4441
rect 114 4428 278 4431
rect 282 4428 342 4431
rect 402 4428 406 4431
rect 538 4428 582 4431
rect 586 4428 646 4431
rect 678 4431 681 4438
rect 678 4428 750 4431
rect 754 4428 822 4431
rect 1034 4428 1102 4431
rect 1706 4428 1798 4431
rect 1802 4428 2422 4431
rect 2426 4428 2438 4431
rect 2466 4428 2470 4431
rect 2666 4428 2686 4431
rect 2734 4428 2806 4431
rect 3194 4428 3238 4431
rect 3402 4428 3502 4431
rect 4162 4428 4278 4431
rect 194 4418 278 4421
rect 378 4418 550 4421
rect 554 4418 662 4421
rect 794 4418 862 4421
rect 950 4421 953 4428
rect 2734 4422 2737 4428
rect 882 4418 953 4421
rect 1346 4418 2198 4421
rect 2282 4418 2326 4421
rect 2330 4418 2358 4421
rect 2362 4418 2542 4421
rect 2546 4418 2718 4421
rect 2770 4418 3494 4421
rect 3642 4418 3982 4421
rect 4170 4418 4230 4421
rect 4266 4418 4886 4421
rect 5018 4418 5134 4421
rect 5138 4418 5142 4421
rect 5210 4418 5222 4421
rect 130 4408 190 4411
rect 826 4408 926 4411
rect 1250 4408 1302 4411
rect 1706 4408 1726 4411
rect 1730 4408 2070 4411
rect 2418 4408 2558 4411
rect 2594 4408 3262 4411
rect 4506 4408 4870 4411
rect 328 4403 330 4407
rect 334 4403 337 4407
rect 342 4403 344 4407
rect 550 4402 553 4408
rect 726 4402 729 4408
rect 1352 4403 1354 4407
rect 1358 4403 1361 4407
rect 1366 4403 1368 4407
rect 2384 4403 2386 4407
rect 2390 4403 2393 4407
rect 2398 4403 2400 4407
rect 3400 4403 3402 4407
rect 3406 4403 3409 4407
rect 3414 4403 3416 4407
rect 3710 4402 3713 4408
rect 4424 4403 4426 4407
rect 4430 4403 4433 4407
rect 4438 4403 4440 4407
rect 418 4398 494 4401
rect 610 4398 702 4401
rect 802 4398 918 4401
rect 1010 4398 1230 4401
rect 1394 4398 1414 4401
rect 1418 4398 1846 4401
rect 2114 4398 2158 4401
rect 2162 4398 2262 4401
rect 2578 4398 3046 4401
rect 3050 4398 3070 4401
rect 3090 4398 3134 4401
rect 3834 4398 4166 4401
rect 4346 4398 4350 4401
rect 4594 4398 4846 4401
rect 82 4388 142 4391
rect 218 4388 230 4391
rect 282 4388 950 4391
rect 954 4388 982 4391
rect 1098 4388 1310 4391
rect 2434 4388 2446 4391
rect 2450 4388 2494 4391
rect 2498 4388 2710 4391
rect 2762 4388 3150 4391
rect 3490 4388 3614 4391
rect 3666 4388 3694 4391
rect 4386 4388 4702 4391
rect 4770 4388 4798 4391
rect 50 4378 174 4381
rect 202 4378 214 4381
rect 370 4378 494 4381
rect 526 4378 558 4381
rect 626 4378 726 4381
rect 730 4378 1134 4381
rect 1218 4378 1598 4381
rect 2154 4378 2374 4381
rect 2394 4378 2446 4381
rect 2458 4378 2566 4381
rect 2570 4378 2670 4381
rect 2722 4378 2870 4381
rect 2986 4378 3126 4381
rect 3450 4378 3622 4381
rect 3770 4378 3782 4381
rect 3882 4378 4094 4381
rect 4634 4378 4654 4381
rect 526 4372 529 4378
rect 1926 4372 1929 4378
rect 106 4368 246 4371
rect 250 4368 278 4371
rect 282 4368 302 4371
rect 306 4368 318 4371
rect 394 4368 398 4371
rect 402 4368 526 4371
rect 706 4368 798 4371
rect 806 4368 918 4371
rect 978 4368 1014 4371
rect 1034 4368 1078 4371
rect 1082 4368 1326 4371
rect 1754 4368 1894 4371
rect 1898 4368 1918 4371
rect 1954 4368 2070 4371
rect 2074 4368 2182 4371
rect 2186 4368 2326 4371
rect 2418 4368 2422 4371
rect 2482 4368 2534 4371
rect 2570 4368 2582 4371
rect 2590 4368 2662 4371
rect 2802 4368 3022 4371
rect 3382 4371 3385 4378
rect 5038 4372 5041 4378
rect 3382 4368 3414 4371
rect 3666 4368 3942 4371
rect 4298 4368 4406 4371
rect 4650 4368 4782 4371
rect 5050 4368 5062 4371
rect 638 4362 641 4368
rect 806 4362 809 4368
rect 82 4358 102 4361
rect 106 4358 126 4361
rect 146 4358 342 4361
rect 362 4358 374 4361
rect 578 4358 606 4361
rect 610 4358 622 4361
rect 666 4358 742 4361
rect 1186 4358 1190 4361
rect 1258 4358 1326 4361
rect 1330 4358 1470 4361
rect 1474 4358 1478 4361
rect 1602 4358 1614 4361
rect 1622 4361 1625 4368
rect 1622 4358 1726 4361
rect 1770 4358 1830 4361
rect 1942 4361 1945 4368
rect 1938 4358 1945 4361
rect 2090 4358 2150 4361
rect 2330 4358 2446 4361
rect 2590 4361 2593 4368
rect 2482 4358 2593 4361
rect 2686 4361 2689 4368
rect 2774 4362 2777 4368
rect 2686 4358 2694 4361
rect 3442 4358 3518 4361
rect 3558 4361 3561 4368
rect 4086 4362 4089 4368
rect 4134 4362 4137 4368
rect 3554 4358 3561 4361
rect 3690 4358 3838 4361
rect 3850 4358 3862 4361
rect 3898 4358 3902 4361
rect 4010 4358 4030 4361
rect 4178 4358 4206 4361
rect 4210 4358 4214 4361
rect 4458 4358 4638 4361
rect 4650 4358 4654 4361
rect 4858 4358 4878 4361
rect 4882 4358 4894 4361
rect 5034 4358 5062 4361
rect 5122 4358 5142 4361
rect 5154 4358 5177 4361
rect 26 4348 102 4351
rect 162 4348 198 4351
rect 258 4348 270 4351
rect 274 4348 302 4351
rect 338 4348 366 4351
rect 386 4348 390 4351
rect 458 4348 462 4351
rect 610 4348 646 4351
rect 746 4348 774 4351
rect 802 4348 806 4351
rect 882 4348 886 4351
rect 970 4348 1006 4351
rect 1026 4348 1046 4351
rect 1154 4348 1158 4351
rect 1194 4348 1262 4351
rect 1410 4348 1486 4351
rect 1546 4348 1566 4351
rect 1618 4348 1657 4351
rect 1682 4348 1718 4351
rect 1722 4348 1766 4351
rect 1990 4351 1993 4358
rect 1862 4348 1993 4351
rect 2106 4348 2190 4351
rect 2222 4351 2225 4358
rect 2222 4348 2238 4351
rect 2242 4348 2342 4351
rect 2370 4348 2414 4351
rect 2418 4348 2502 4351
rect 2606 4351 2609 4358
rect 2530 4348 2609 4351
rect 2638 4351 2641 4358
rect 2638 4348 2713 4351
rect 2730 4348 2734 4351
rect 2754 4348 2766 4351
rect 2834 4348 2838 4351
rect 3014 4351 3017 4358
rect 3070 4351 3073 4358
rect 3014 4348 3073 4351
rect 90 4338 94 4341
rect 406 4341 409 4348
rect 406 4338 462 4341
rect 586 4338 598 4341
rect 690 4338 694 4341
rect 702 4341 705 4348
rect 1654 4342 1657 4348
rect 1862 4342 1865 4348
rect 2422 4342 2425 4348
rect 2518 4342 2521 4348
rect 2710 4342 2713 4348
rect 2798 4342 2801 4348
rect 702 4338 830 4341
rect 938 4338 958 4341
rect 978 4338 1030 4341
rect 1186 4338 1222 4341
rect 1386 4338 1606 4341
rect 2290 4338 2366 4341
rect 2450 4338 2510 4341
rect 2722 4338 2726 4341
rect 2894 4341 2897 4348
rect 3330 4348 3334 4351
rect 3378 4348 3390 4351
rect 3402 4348 3406 4351
rect 3538 4348 3550 4351
rect 3722 4348 3774 4351
rect 3786 4348 3790 4351
rect 3794 4348 3854 4351
rect 3882 4348 3886 4351
rect 3930 4348 3934 4351
rect 3978 4348 4022 4351
rect 4062 4351 4065 4358
rect 4062 4348 4086 4351
rect 4090 4348 4118 4351
rect 4154 4348 4190 4351
rect 4194 4348 4206 4351
rect 4286 4351 4289 4358
rect 5174 4352 5177 4358
rect 4234 4348 4289 4351
rect 4390 4348 4398 4351
rect 4402 4348 4478 4351
rect 4498 4348 4713 4351
rect 4770 4348 4806 4351
rect 4834 4348 4886 4351
rect 4890 4348 4918 4351
rect 5106 4348 5118 4351
rect 2858 4338 3057 4341
rect 3106 4338 3134 4341
rect 3254 4338 3302 4341
rect 3350 4341 3353 4348
rect 3350 4338 3374 4341
rect 3446 4341 3449 4348
rect 4206 4342 4209 4348
rect 4710 4342 4713 4348
rect 3378 4338 3449 4341
rect 3546 4338 3638 4341
rect 3762 4338 3766 4341
rect 3818 4338 3854 4341
rect 3882 4338 4014 4341
rect 4066 4338 4070 4341
rect 4130 4338 4134 4341
rect 4178 4338 4182 4341
rect 4226 4338 4238 4341
rect 4378 4338 4390 4341
rect 4394 4338 4486 4341
rect 4510 4338 4558 4341
rect 4594 4338 4606 4341
rect 4674 4338 4694 4341
rect 4722 4338 4726 4341
rect 4754 4338 4806 4341
rect 4914 4338 5006 4341
rect 5030 4341 5033 4348
rect 5246 4342 5249 4348
rect 5030 4338 5102 4341
rect 5106 4338 5110 4341
rect 566 4332 569 4338
rect 1262 4332 1265 4338
rect 34 4328 150 4331
rect 370 4328 470 4331
rect 490 4328 494 4331
rect 682 4328 694 4331
rect 706 4328 710 4331
rect 802 4328 814 4331
rect 818 4328 974 4331
rect 1034 4328 1110 4331
rect 1138 4328 1246 4331
rect 1330 4328 1446 4331
rect 1538 4328 1542 4331
rect 1558 4328 1582 4331
rect 1602 4328 1734 4331
rect 1738 4328 1878 4331
rect 1962 4328 2054 4331
rect 2170 4328 2574 4331
rect 2758 4331 2761 4338
rect 3054 4332 3057 4338
rect 3254 4332 3257 4338
rect 4510 4332 4513 4338
rect 4622 4332 4625 4338
rect 5198 4332 5201 4338
rect 2758 4328 2798 4331
rect 2874 4328 2878 4331
rect 3426 4328 3510 4331
rect 3514 4328 3518 4331
rect 3546 4328 3694 4331
rect 3802 4328 3822 4331
rect 3834 4328 3838 4331
rect 4002 4328 4054 4331
rect 4114 4328 4126 4331
rect 4250 4328 4350 4331
rect 1558 4322 1561 4328
rect 258 4318 462 4321
rect 466 4318 510 4321
rect 602 4318 734 4321
rect 750 4318 758 4321
rect 762 4318 937 4321
rect 946 4318 958 4321
rect 1450 4318 1454 4321
rect 1762 4318 1782 4321
rect 1818 4318 1902 4321
rect 1906 4318 1990 4321
rect 2018 4318 2046 4321
rect 2150 4321 2153 4328
rect 2150 4318 2238 4321
rect 2494 4318 2502 4321
rect 2506 4318 2734 4321
rect 2822 4321 2825 4328
rect 2778 4318 2825 4321
rect 2834 4318 2934 4321
rect 3042 4318 3118 4321
rect 3242 4318 3254 4321
rect 3282 4318 3286 4321
rect 3290 4318 3366 4321
rect 3386 4318 3390 4321
rect 3498 4318 3953 4321
rect 4250 4318 4358 4321
rect 4362 4318 4422 4321
rect 4450 4318 4518 4321
rect 4522 4318 4622 4321
rect 4774 4321 4777 4328
rect 4774 4318 4790 4321
rect 5046 4321 5049 4328
rect 4914 4318 5049 4321
rect 5074 4318 5246 4321
rect 5250 4318 5278 4321
rect 218 4308 494 4311
rect 562 4308 590 4311
rect 594 4308 766 4311
rect 934 4311 937 4318
rect 934 4308 1054 4311
rect 1594 4308 1726 4311
rect 1818 4308 1846 4311
rect 1978 4308 1990 4311
rect 2002 4308 2150 4311
rect 2234 4308 2262 4311
rect 2490 4308 2550 4311
rect 2698 4308 2726 4311
rect 2994 4308 3270 4311
rect 3274 4308 3526 4311
rect 3770 4308 3830 4311
rect 3842 4308 3870 4311
rect 3950 4311 3953 4318
rect 3950 4308 4046 4311
rect 4410 4308 4542 4311
rect 4618 4308 4870 4311
rect 4874 4308 4926 4311
rect 5178 4308 5182 4311
rect 848 4303 850 4307
rect 854 4303 857 4307
rect 862 4303 864 4307
rect 1872 4303 1874 4307
rect 1878 4303 1881 4307
rect 1886 4303 1888 4307
rect 2888 4303 2890 4307
rect 2894 4303 2897 4307
rect 2902 4303 2904 4307
rect 3920 4303 3922 4307
rect 3926 4303 3929 4307
rect 3934 4303 3936 4307
rect 4936 4303 4938 4307
rect 4942 4303 4945 4307
rect 4950 4303 4952 4307
rect 10 4298 22 4301
rect 122 4298 134 4301
rect 138 4298 166 4301
rect 418 4298 486 4301
rect 666 4298 686 4301
rect 1578 4298 1606 4301
rect 1626 4298 1662 4301
rect 1746 4298 1774 4301
rect 1922 4298 2022 4301
rect 2042 4298 2062 4301
rect 2274 4298 2462 4301
rect 3394 4298 3550 4301
rect 3554 4298 3678 4301
rect 3682 4298 3790 4301
rect 3794 4298 3806 4301
rect 4082 4298 4374 4301
rect 4546 4298 4646 4301
rect 5162 4298 5174 4301
rect 5194 4298 5238 4301
rect 4414 4292 4417 4298
rect 18 4288 22 4291
rect 370 4288 534 4291
rect 666 4288 726 4291
rect 738 4288 774 4291
rect 786 4288 870 4291
rect 1050 4288 1198 4291
rect 1442 4288 2462 4291
rect 2562 4288 2574 4291
rect 2594 4288 2678 4291
rect 2778 4288 2841 4291
rect 2970 4288 2982 4291
rect 3042 4288 3126 4291
rect 3178 4288 3222 4291
rect 3634 4288 3902 4291
rect 3914 4288 3974 4291
rect 3978 4288 4062 4291
rect 4106 4288 4110 4291
rect 4338 4288 4398 4291
rect 4474 4288 4526 4291
rect 4642 4288 4646 4291
rect 4874 4288 4958 4291
rect 5154 4288 5198 4291
rect 2838 4282 2841 4288
rect 186 4278 198 4281
rect 218 4278 222 4281
rect 314 4278 374 4281
rect 386 4278 409 4281
rect 418 4278 462 4281
rect 474 4278 566 4281
rect 594 4278 606 4281
rect 706 4278 742 4281
rect 986 4278 1022 4281
rect 1090 4278 1094 4281
rect 1354 4278 1358 4281
rect 1362 4278 1398 4281
rect 1426 4278 1510 4281
rect 1682 4278 1686 4281
rect 1754 4278 1766 4281
rect 1826 4278 2054 4281
rect 2058 4278 2086 4281
rect 2146 4278 2217 4281
rect 2226 4278 2318 4281
rect 2354 4278 2430 4281
rect 2514 4278 2566 4281
rect 2642 4278 2774 4281
rect 2810 4278 2822 4281
rect 2842 4278 2878 4281
rect 2898 4278 2918 4281
rect 3010 4278 3014 4281
rect 3826 4278 3878 4281
rect 3914 4278 3958 4281
rect 3962 4278 4046 4281
rect 4050 4278 4302 4281
rect 4322 4278 4374 4281
rect 4410 4278 4417 4281
rect 4482 4278 4518 4281
rect 4594 4278 4662 4281
rect 4674 4278 4742 4281
rect 4754 4278 4758 4281
rect 4986 4278 5006 4281
rect 5034 4278 5054 4281
rect 5186 4278 5201 4281
rect 102 4271 105 4278
rect 66 4268 105 4271
rect 250 4268 254 4271
rect 370 4268 390 4271
rect 406 4271 409 4278
rect 406 4268 414 4271
rect 434 4268 446 4271
rect 482 4268 526 4271
rect 546 4268 582 4271
rect 694 4271 697 4278
rect 674 4268 697 4271
rect 714 4268 726 4271
rect 746 4268 758 4271
rect 790 4268 838 4271
rect 866 4268 985 4271
rect 994 4268 1022 4271
rect 1082 4268 1102 4271
rect 1190 4271 1193 4278
rect 1654 4272 1657 4278
rect 2214 4272 2217 4278
rect 1122 4268 1193 4271
rect 1298 4268 1302 4271
rect 1306 4268 1326 4271
rect 1434 4268 1486 4271
rect 1554 4268 1606 4271
rect 1690 4268 1694 4271
rect 1746 4268 1926 4271
rect 1930 4268 2014 4271
rect 2026 4268 2142 4271
rect 2178 4268 2206 4271
rect 2362 4268 2366 4271
rect 2434 4268 2438 4271
rect 2462 4271 2465 4278
rect 2450 4268 2465 4271
rect 2470 4272 2473 4278
rect 2482 4268 2486 4271
rect 2730 4268 2798 4271
rect 2982 4271 2985 4278
rect 3166 4272 3169 4278
rect 2866 4268 2985 4271
rect 3010 4268 3070 4271
rect 3174 4271 3177 4278
rect 4414 4272 4417 4278
rect 3174 4268 3182 4271
rect 3202 4268 3206 4271
rect 3738 4268 3742 4271
rect 4122 4268 4134 4271
rect 4154 4268 4158 4271
rect 4210 4268 4214 4271
rect 4258 4268 4262 4271
rect 4274 4268 4278 4271
rect 4354 4268 4398 4271
rect 4498 4268 4590 4271
rect 4594 4268 4638 4271
rect 4642 4268 4878 4271
rect 4882 4268 4990 4271
rect 4994 4268 5006 4271
rect 5142 4271 5145 4278
rect 5066 4268 5145 4271
rect 5166 4272 5169 4278
rect 5198 4272 5201 4278
rect 590 4262 593 4268
rect 790 4262 793 4268
rect 98 4258 102 4261
rect 226 4258 230 4261
rect 234 4258 246 4261
rect 378 4258 422 4261
rect 438 4258 486 4261
rect 610 4258 614 4261
rect 626 4258 686 4261
rect 722 4258 734 4261
rect 770 4258 774 4261
rect 786 4258 790 4261
rect 810 4258 814 4261
rect 874 4258 878 4261
rect 930 4258 958 4261
rect 962 4258 974 4261
rect 982 4261 985 4268
rect 982 4258 1025 4261
rect 1066 4258 1142 4261
rect 1146 4258 1166 4261
rect 1298 4258 1382 4261
rect 1410 4258 1446 4261
rect 1542 4261 1545 4268
rect 1514 4258 1545 4261
rect 1742 4261 1745 4268
rect 2814 4262 2817 4268
rect 3270 4262 3273 4268
rect 1658 4258 1745 4261
rect 1754 4258 1822 4261
rect 1826 4258 1830 4261
rect 1834 4258 1934 4261
rect 2066 4258 2105 4261
rect 438 4252 441 4258
rect 1022 4252 1025 4258
rect 2102 4252 2105 4258
rect 2202 4258 2510 4261
rect 2570 4258 2574 4261
rect 2918 4258 3230 4261
rect 3234 4258 3262 4261
rect 3322 4258 3390 4261
rect 3594 4258 3598 4261
rect 3654 4261 3657 4268
rect 3610 4258 3657 4261
rect 3690 4258 3694 4261
rect 3714 4258 3750 4261
rect 3878 4261 3881 4268
rect 3786 4258 3881 4261
rect 4030 4261 4033 4268
rect 4030 4258 4078 4261
rect 4110 4261 4113 4268
rect 5022 4262 5025 4268
rect 5054 4262 5057 4268
rect 4110 4258 4118 4261
rect 4162 4258 4286 4261
rect 4330 4258 4406 4261
rect 4570 4258 4582 4261
rect 4602 4258 4702 4261
rect 4762 4258 4790 4261
rect 4818 4258 4822 4261
rect 4842 4258 4846 4261
rect 4926 4258 5014 4261
rect 5114 4258 5126 4261
rect 5130 4258 5182 4261
rect 2126 4252 2129 4258
rect 2534 4252 2537 4258
rect 18 4248 118 4251
rect 226 4248 302 4251
rect 306 4248 318 4251
rect 362 4248 406 4251
rect 538 4248 638 4251
rect 658 4248 950 4251
rect 954 4248 1014 4251
rect 1042 4248 1366 4251
rect 1370 4248 1670 4251
rect 1738 4248 1750 4251
rect 1758 4248 1777 4251
rect 1786 4248 1814 4251
rect 1842 4248 1926 4251
rect 2162 4248 2190 4251
rect 2210 4248 2254 4251
rect 2282 4248 2438 4251
rect 2714 4248 2817 4251
rect 2918 4251 2921 4258
rect 3558 4252 3561 4258
rect 2834 4248 2921 4251
rect 2930 4248 2937 4251
rect 2954 4248 2958 4251
rect 3018 4248 3030 4251
rect 3154 4248 3246 4251
rect 3522 4248 3526 4251
rect 3670 4248 3702 4251
rect 3706 4248 3790 4251
rect 4074 4248 4110 4251
rect 4210 4248 4214 4251
rect 4234 4248 4262 4251
rect 4282 4248 4294 4251
rect 4422 4251 4425 4258
rect 4926 4252 4929 4258
rect 4370 4248 4425 4251
rect 4554 4248 4566 4251
rect 4802 4248 4806 4251
rect 106 4238 150 4241
rect 386 4238 398 4241
rect 426 4238 566 4241
rect 626 4238 825 4241
rect 834 4238 870 4241
rect 874 4238 950 4241
rect 1282 4238 1422 4241
rect 1694 4241 1697 4248
rect 1506 4238 1697 4241
rect 1758 4242 1761 4248
rect 1774 4242 1777 4248
rect 1966 4242 1969 4248
rect 2814 4242 2817 4248
rect 2934 4242 2937 4248
rect 1866 4238 1958 4241
rect 2002 4238 2198 4241
rect 2210 4238 2382 4241
rect 2386 4238 2486 4241
rect 2498 4238 2782 4241
rect 2858 4238 2910 4241
rect 2922 4238 2926 4241
rect 2954 4238 3166 4241
rect 3170 4238 3454 4241
rect 3630 4241 3633 4248
rect 3490 4238 3633 4241
rect 3670 4242 3673 4248
rect 3798 4241 3801 4248
rect 3786 4238 3801 4241
rect 4098 4238 4734 4241
rect 4858 4238 5046 4241
rect 5146 4238 5206 4241
rect 234 4228 294 4231
rect 298 4228 326 4231
rect 330 4228 406 4231
rect 570 4228 814 4231
rect 822 4231 825 4238
rect 822 4228 1086 4231
rect 1090 4228 1126 4231
rect 1130 4228 1150 4231
rect 1978 4228 2054 4231
rect 2074 4228 2590 4231
rect 2770 4228 2774 4231
rect 2802 4228 2862 4231
rect 2874 4228 3014 4231
rect 3386 4228 3550 4231
rect 3562 4228 4150 4231
rect 4354 4228 4646 4231
rect 4778 4228 5022 4231
rect 5026 4228 5182 4231
rect 242 4218 470 4221
rect 482 4218 710 4221
rect 858 4218 1182 4221
rect 1498 4218 1734 4221
rect 1814 4221 1817 4228
rect 1778 4218 1817 4221
rect 1930 4218 2054 4221
rect 2338 4218 2510 4221
rect 2582 4218 2662 4221
rect 2818 4218 2934 4221
rect 3098 4218 3278 4221
rect 3450 4218 3454 4221
rect 3498 4218 3614 4221
rect 3618 4218 3670 4221
rect 3818 4218 3950 4221
rect 3954 4218 4134 4221
rect 4150 4221 4153 4228
rect 4150 4218 4814 4221
rect 4818 4218 5110 4221
rect 5122 4218 5166 4221
rect 718 4212 721 4218
rect 2582 4212 2585 4218
rect 394 4208 494 4211
rect 554 4208 582 4211
rect 818 4208 878 4211
rect 1482 4208 1502 4211
rect 1746 4208 1966 4211
rect 1994 4208 2190 4211
rect 2706 4208 2862 4211
rect 2866 4208 2982 4211
rect 2986 4208 3022 4211
rect 3802 4208 4006 4211
rect 4018 4208 4094 4211
rect 4186 4208 4222 4211
rect 4482 4208 5030 4211
rect 5162 4208 5190 4211
rect 328 4203 330 4207
rect 334 4203 337 4207
rect 342 4203 344 4207
rect 1352 4203 1354 4207
rect 1358 4203 1361 4207
rect 1366 4203 1368 4207
rect 2384 4203 2386 4207
rect 2390 4203 2393 4207
rect 2398 4203 2400 4207
rect 3400 4203 3402 4207
rect 3406 4203 3409 4207
rect 3414 4203 3416 4207
rect 4424 4203 4426 4207
rect 4430 4203 4433 4207
rect 4438 4203 4440 4207
rect 82 4198 142 4201
rect 474 4198 726 4201
rect 818 4198 886 4201
rect 1770 4198 1814 4201
rect 1994 4198 1998 4201
rect 2050 4198 2238 4201
rect 2450 4198 2470 4201
rect 2754 4198 2854 4201
rect 3026 4198 3286 4201
rect 3290 4198 3302 4201
rect 3762 4198 4182 4201
rect 4186 4198 4398 4201
rect 4530 4198 4766 4201
rect 4842 4198 5198 4201
rect 146 4188 214 4191
rect 218 4188 350 4191
rect 370 4188 558 4191
rect 634 4188 918 4191
rect 1394 4188 1470 4191
rect 1474 4188 1526 4191
rect 1530 4188 1566 4191
rect 1570 4188 1646 4191
rect 1650 4188 1694 4191
rect 1730 4188 1782 4191
rect 1814 4191 1817 4198
rect 1814 4188 1838 4191
rect 1842 4188 1878 4191
rect 1922 4188 2086 4191
rect 2098 4188 2142 4191
rect 2202 4188 2214 4191
rect 2458 4188 2550 4191
rect 2842 4188 3046 4191
rect 3050 4188 3702 4191
rect 3770 4188 3790 4191
rect 3826 4188 4262 4191
rect 4362 4188 4782 4191
rect 4786 4188 4846 4191
rect 5114 4188 5230 4191
rect 146 4178 174 4181
rect 178 4178 262 4181
rect 266 4178 390 4181
rect 538 4178 702 4181
rect 1250 4178 1294 4181
rect 1402 4178 1446 4181
rect 1450 4178 1550 4181
rect 1554 4178 1798 4181
rect 2302 4181 2305 4188
rect 2774 4182 2777 4188
rect 1802 4178 2305 4181
rect 2466 4178 2526 4181
rect 2786 4178 3025 4181
rect 3082 4178 3182 4181
rect 3322 4178 3502 4181
rect 3506 4178 3630 4181
rect 3634 4178 3662 4181
rect 3666 4178 3726 4181
rect 3730 4178 3774 4181
rect 3834 4178 4046 4181
rect 4170 4178 4198 4181
rect 4306 4178 4326 4181
rect 4330 4178 4390 4181
rect 4562 4178 4737 4181
rect 4746 4178 5110 4181
rect 5138 4178 5262 4181
rect 3022 4172 3025 4178
rect 18 4168 22 4171
rect 154 4168 326 4171
rect 330 4168 430 4171
rect 482 4168 598 4171
rect 602 4168 646 4171
rect 682 4168 686 4171
rect 706 4168 710 4171
rect 898 4168 910 4171
rect 914 4168 974 4171
rect 978 4168 1078 4171
rect 1178 4168 1414 4171
rect 1682 4168 1806 4171
rect 1886 4168 1934 4171
rect 2082 4168 2190 4171
rect 2210 4168 2406 4171
rect 2722 4168 2758 4171
rect 2762 4168 2814 4171
rect 3242 4168 3470 4171
rect 3530 4168 3614 4171
rect 3642 4168 3982 4171
rect 4070 4171 4073 4178
rect 4734 4172 4737 4178
rect 4070 4168 4102 4171
rect 4194 4168 4206 4171
rect 4322 4168 4350 4171
rect 4370 4168 4566 4171
rect 4650 4168 4670 4171
rect 5074 4168 5190 4171
rect 1206 4162 1209 4168
rect 214 4158 249 4161
rect 290 4158 414 4161
rect 506 4158 510 4161
rect 538 4158 574 4161
rect 634 4158 694 4161
rect 698 4158 726 4161
rect 1226 4158 1286 4161
rect 1466 4158 1478 4161
rect 1486 4161 1489 4168
rect 1830 4162 1833 4168
rect 1886 4162 1889 4168
rect 1486 4158 1574 4161
rect 1658 4158 1734 4161
rect 1906 4158 2030 4161
rect 2074 4158 2102 4161
rect 2598 4161 2601 4168
rect 5278 4162 5281 4168
rect 2586 4158 2601 4161
rect 2746 4158 2782 4161
rect 2806 4158 2814 4161
rect 2818 4158 2878 4161
rect 3042 4158 3046 4161
rect 3114 4158 3150 4161
rect 3322 4158 3478 4161
rect 3498 4158 3510 4161
rect 3522 4158 3622 4161
rect 3738 4158 3785 4161
rect 3794 4158 3806 4161
rect 3906 4158 4150 4161
rect 4186 4158 4214 4161
rect 4346 4158 4350 4161
rect 4698 4158 4710 4161
rect 4890 4158 4894 4161
rect 5154 4158 5222 4161
rect 214 4152 217 4158
rect 246 4152 249 4158
rect 1174 4152 1177 4158
rect 114 4148 134 4151
rect 170 4148 214 4151
rect 314 4148 374 4151
rect 498 4148 534 4151
rect 618 4148 654 4151
rect 674 4148 758 4151
rect 770 4148 830 4151
rect 834 4148 838 4151
rect 1122 4148 1166 4151
rect 1290 4148 1382 4151
rect 1386 4148 1502 4151
rect 1734 4151 1737 4158
rect 1722 4148 1737 4151
rect 1930 4148 1969 4151
rect 390 4141 393 4148
rect 1854 4142 1857 4148
rect 1966 4142 1969 4148
rect 2170 4148 2174 4151
rect 2194 4148 2198 4151
rect 2314 4148 2350 4151
rect 2354 4148 2438 4151
rect 2458 4148 2558 4151
rect 2650 4148 2814 4151
rect 2818 4148 3134 4151
rect 3138 4148 3286 4151
rect 3406 4148 3478 4151
rect 3662 4151 3665 4158
rect 3514 4148 3561 4151
rect 3662 4148 3742 4151
rect 3782 4151 3785 4158
rect 3782 4148 3862 4151
rect 3962 4148 4030 4151
rect 4034 4148 4086 4151
rect 4098 4148 4126 4151
rect 4194 4148 4230 4151
rect 4234 4148 4246 4151
rect 4250 4148 4470 4151
rect 4518 4151 4521 4158
rect 4518 4148 4606 4151
rect 4642 4148 4702 4151
rect 4706 4148 4710 4151
rect 4762 4148 4790 4151
rect 4874 4148 4990 4151
rect 5082 4148 5158 4151
rect 5214 4148 5238 4151
rect 2134 4142 2137 4148
rect 2246 4142 2249 4148
rect 2614 4142 2617 4148
rect 98 4138 393 4141
rect 506 4138 510 4141
rect 522 4138 582 4141
rect 586 4138 622 4141
rect 690 4138 750 4141
rect 906 4138 918 4141
rect 1210 4138 1222 4141
rect 1258 4138 1313 4141
rect 1442 4138 1454 4141
rect 1586 4138 1758 4141
rect 1874 4138 1878 4141
rect 1906 4138 1910 4141
rect 2114 4138 2121 4141
rect 2194 4138 2206 4141
rect 2362 4138 2430 4141
rect 2622 4141 2625 4148
rect 3406 4142 3409 4148
rect 3558 4142 3561 4148
rect 4734 4142 4737 4148
rect 2622 4138 2694 4141
rect 2786 4138 2790 4141
rect 2826 4138 3022 4141
rect 3042 4138 3086 4141
rect 3106 4138 3110 4141
rect 3154 4138 3238 4141
rect 3250 4138 3334 4141
rect 3458 4138 3545 4141
rect 3746 4138 3790 4141
rect 3858 4138 3982 4141
rect 3986 4138 4158 4141
rect 4162 4138 4166 4141
rect 4178 4138 4302 4141
rect 4330 4138 4358 4141
rect 4394 4138 4430 4141
rect 4490 4138 4598 4141
rect 4602 4138 4614 4141
rect 4634 4138 4638 4141
rect 4682 4138 4694 4141
rect 4858 4138 4878 4141
rect 4898 4138 4910 4141
rect 4930 4138 5150 4141
rect 5174 4141 5177 4148
rect 5154 4138 5177 4141
rect 5214 4142 5217 4148
rect 478 4132 481 4138
rect 1310 4132 1313 4138
rect 122 4128 206 4131
rect 210 4128 270 4131
rect 282 4128 350 4131
rect 506 4128 526 4131
rect 634 4128 638 4131
rect 650 4128 822 4131
rect 1234 4128 1294 4131
rect 1338 4128 1390 4131
rect 1570 4128 1606 4131
rect 1698 4128 1822 4131
rect 2046 4131 2049 4138
rect 3278 4132 3281 4138
rect 2046 4128 2078 4131
rect 2114 4128 2118 4131
rect 2322 4128 2326 4131
rect 2330 4128 2510 4131
rect 2562 4128 2646 4131
rect 2722 4128 2726 4131
rect 2730 4128 2870 4131
rect 3010 4128 3078 4131
rect 3082 4128 3254 4131
rect 3290 4128 3326 4131
rect 3358 4131 3361 4138
rect 3542 4132 3545 4138
rect 3358 4128 3446 4131
rect 3570 4128 3686 4131
rect 4042 4128 4046 4131
rect 4066 4128 4398 4131
rect 4402 4128 4606 4131
rect 4714 4128 4742 4131
rect 4842 4128 4902 4131
rect 5098 4128 5110 4131
rect 5246 4131 5249 4138
rect 5114 4128 5249 4131
rect 542 4122 545 4128
rect 550 4122 553 4128
rect 170 4118 366 4121
rect 386 4118 534 4121
rect 570 4118 790 4121
rect 802 4118 950 4121
rect 1178 4118 1238 4121
rect 1242 4118 1278 4121
rect 1314 4118 1326 4121
rect 1362 4118 1382 4121
rect 1534 4121 1537 4128
rect 1426 4118 1537 4121
rect 1626 4118 1742 4121
rect 1818 4118 1822 4121
rect 1826 4118 1902 4121
rect 1954 4118 2086 4121
rect 2402 4118 2486 4121
rect 2570 4118 2630 4121
rect 2642 4118 2678 4121
rect 2682 4118 2734 4121
rect 2746 4118 2766 4121
rect 2770 4118 2934 4121
rect 2938 4118 3190 4121
rect 3458 4118 3782 4121
rect 3786 4118 3902 4121
rect 3914 4118 4062 4121
rect 4258 4118 4278 4121
rect 4282 4118 4310 4121
rect 4314 4118 4382 4121
rect 4522 4118 4662 4121
rect 4714 4118 4726 4121
rect 5050 4118 5198 4121
rect 74 4108 86 4111
rect 138 4108 158 4111
rect 522 4108 622 4111
rect 642 4108 694 4111
rect 1010 4108 1286 4111
rect 1290 4108 1462 4111
rect 1538 4108 1630 4111
rect 1690 4108 1830 4111
rect 1922 4108 1974 4111
rect 1978 4108 2342 4111
rect 2370 4108 2534 4111
rect 2538 4108 2582 4111
rect 2674 4108 2798 4111
rect 2802 4108 2814 4111
rect 3026 4108 3198 4111
rect 3210 4108 3470 4111
rect 3474 4108 3494 4111
rect 3498 4108 3518 4111
rect 3626 4108 3758 4111
rect 4042 4108 4102 4111
rect 4210 4108 4278 4111
rect 4346 4108 4374 4111
rect 4402 4108 4494 4111
rect 4714 4108 4822 4111
rect 5186 4108 5198 4111
rect 848 4103 850 4107
rect 854 4103 857 4107
rect 862 4103 864 4107
rect 1872 4103 1874 4107
rect 1878 4103 1881 4107
rect 1886 4103 1888 4107
rect 2888 4103 2890 4107
rect 2894 4103 2897 4107
rect 2902 4103 2904 4107
rect 3920 4103 3922 4107
rect 3926 4103 3929 4107
rect 3934 4103 3936 4107
rect 4936 4103 4938 4107
rect 4942 4103 4945 4107
rect 4950 4103 4952 4107
rect 138 4098 254 4101
rect 322 4098 438 4101
rect 546 4098 710 4101
rect 1178 4098 1566 4101
rect 1650 4098 1734 4101
rect 2034 4098 2166 4101
rect 2174 4098 2366 4101
rect 2434 4098 2526 4101
rect 2554 4098 2574 4101
rect 2618 4098 2622 4101
rect 2626 4098 2686 4101
rect 2690 4098 2774 4101
rect 3202 4098 3310 4101
rect 3490 4098 3494 4101
rect 3642 4098 3790 4101
rect 3794 4098 3846 4101
rect 4066 4098 4262 4101
rect 4290 4098 4510 4101
rect 4634 4098 4654 4101
rect 4730 4098 4750 4101
rect 5130 4098 5142 4101
rect 5146 4098 5222 4101
rect 202 4088 206 4091
rect 466 4088 566 4091
rect 578 4088 606 4091
rect 610 4088 678 4091
rect 770 4088 870 4091
rect 1098 4088 1246 4091
rect 1298 4088 1390 4091
rect 1710 4088 1758 4091
rect 1850 4088 1926 4091
rect 1938 4088 1998 4091
rect 2174 4091 2177 4098
rect 2002 4088 2177 4091
rect 2634 4088 2830 4091
rect 2834 4088 2846 4091
rect 2850 4088 2918 4091
rect 2938 4088 2998 4091
rect 3122 4088 3126 4091
rect 3442 4088 3646 4091
rect 3722 4088 3766 4091
rect 3770 4088 3814 4091
rect 3886 4088 4030 4091
rect 4034 4088 4046 4091
rect 4070 4088 4222 4091
rect 4362 4088 4366 4091
rect 4970 4088 5134 4091
rect 5170 4088 5182 4091
rect 210 4078 230 4081
rect 234 4078 358 4081
rect 390 4081 393 4088
rect 1710 4082 1713 4088
rect 390 4078 414 4081
rect 546 4078 558 4081
rect 562 4078 630 4081
rect 842 4078 982 4081
rect 1050 4078 1342 4081
rect 1362 4078 1430 4081
rect 1482 4078 1606 4081
rect 1722 4078 1726 4081
rect 1746 4078 1758 4081
rect 1778 4078 1782 4081
rect 1842 4078 1918 4081
rect 1938 4078 1942 4081
rect 1954 4078 2038 4081
rect 2106 4078 2230 4081
rect 2242 4078 2334 4081
rect 2378 4078 2406 4081
rect 2506 4078 2598 4081
rect 2802 4078 2926 4081
rect 3010 4078 3118 4081
rect 3186 4078 3222 4081
rect 3270 4081 3273 4088
rect 3234 4078 3273 4081
rect 3278 4081 3281 4088
rect 3886 4082 3889 4088
rect 4070 4082 4073 4088
rect 3278 4078 3302 4081
rect 3346 4078 3350 4081
rect 3458 4078 3606 4081
rect 3610 4078 3638 4081
rect 3714 4078 3718 4081
rect 3898 4078 3902 4081
rect 3914 4078 4006 4081
rect 4010 4078 4054 4081
rect 4338 4078 4374 4081
rect 5186 4078 5190 4081
rect 726 4072 729 4078
rect 1190 4072 1193 4078
rect 2454 4072 2457 4078
rect 162 4068 182 4071
rect 258 4068 345 4071
rect 362 4068 582 4071
rect 682 4068 702 4071
rect 946 4068 998 4071
rect 1378 4068 1398 4071
rect 1538 4068 1550 4071
rect 1554 4068 2126 4071
rect 2138 4068 2454 4071
rect 2462 4071 2465 4078
rect 4230 4072 4233 4078
rect 2462 4068 2558 4071
rect 2562 4068 2598 4071
rect 2698 4068 2702 4071
rect 2706 4068 2782 4071
rect 3018 4068 3022 4071
rect 3050 4068 3054 4071
rect 3194 4068 4054 4071
rect 4114 4068 4198 4071
rect 4242 4068 4262 4071
rect 4290 4068 4294 4071
rect 4330 4068 4390 4071
rect 4530 4068 4614 4071
rect 4618 4068 4646 4071
rect 4710 4071 4713 4078
rect 4806 4071 4809 4078
rect 4918 4071 4921 4078
rect 5046 4072 5049 4078
rect 4710 4068 5006 4071
rect 5262 4068 5270 4071
rect 342 4062 345 4068
rect 1502 4062 1505 4068
rect 74 4058 198 4061
rect 290 4058 302 4061
rect 346 4058 414 4061
rect 418 4058 422 4061
rect 434 4058 454 4061
rect 458 4058 478 4061
rect 486 4058 518 4061
rect 538 4058 550 4061
rect 562 4058 566 4061
rect 578 4058 614 4061
rect 650 4058 670 4061
rect 698 4058 814 4061
rect 882 4058 910 4061
rect 914 4058 950 4061
rect 1154 4058 1166 4061
rect 1306 4058 1326 4061
rect 1602 4058 1654 4061
rect 1714 4058 1718 4061
rect 1754 4058 1798 4061
rect 1806 4058 1830 4061
rect 1850 4058 1950 4061
rect 1962 4058 1966 4061
rect 1986 4058 2014 4061
rect 2082 4058 2150 4061
rect 2242 4058 2302 4061
rect 2426 4058 2446 4061
rect 2498 4058 2590 4061
rect 2610 4058 2718 4061
rect 2722 4058 2830 4061
rect 2894 4061 2897 4068
rect 3094 4062 3097 4068
rect 2894 4058 2950 4061
rect 2954 4058 2966 4061
rect 2970 4058 3006 4061
rect 3074 4058 3094 4061
rect 3106 4058 3214 4061
rect 3218 4058 3262 4061
rect 3394 4059 3430 4061
rect 4086 4062 4089 4068
rect 4414 4062 4417 4068
rect 3394 4058 3433 4059
rect 3442 4058 3470 4061
rect 3474 4058 3502 4061
rect 3634 4058 3638 4061
rect 3714 4058 3742 4061
rect 3826 4058 3990 4061
rect 4050 4058 4078 4061
rect 4170 4058 4206 4061
rect 4258 4058 4294 4061
rect 4486 4058 4566 4061
rect 4674 4058 4886 4061
rect 5050 4058 5166 4061
rect 5262 4061 5265 4068
rect 5170 4058 5265 4061
rect 94 4048 102 4051
rect 154 4048 158 4051
rect 258 4048 278 4051
rect 302 4048 374 4051
rect 486 4051 489 4058
rect 418 4048 489 4051
rect 498 4048 718 4051
rect 838 4051 841 4058
rect 838 4048 878 4051
rect 902 4048 934 4051
rect 1114 4048 1158 4051
rect 1394 4048 1398 4051
rect 1502 4048 1662 4051
rect 1806 4051 1809 4058
rect 3774 4052 3777 4058
rect 4486 4052 4489 4058
rect 5166 4052 5169 4058
rect 1794 4048 1809 4051
rect 1834 4048 1846 4051
rect 1922 4048 2046 4051
rect 2058 4048 2302 4051
rect 2306 4048 2318 4051
rect 2346 4048 2574 4051
rect 2698 4048 2766 4051
rect 2822 4048 2862 4051
rect 2874 4048 2894 4051
rect 3026 4048 3158 4051
rect 3202 4048 3254 4051
rect 3594 4048 3633 4051
rect 3714 4048 3718 4051
rect 4074 4048 4078 4051
rect 4154 4048 4238 4051
rect 4274 4048 4286 4051
rect 4362 4048 4366 4051
rect 4386 4048 4454 4051
rect 5018 4048 5057 4051
rect 94 4042 97 4048
rect 106 4038 110 4041
rect 254 4041 257 4048
rect 194 4038 257 4041
rect 302 4041 305 4048
rect 902 4042 905 4048
rect 1446 4042 1449 4048
rect 1502 4042 1505 4048
rect 274 4038 305 4041
rect 314 4038 438 4041
rect 442 4038 470 4041
rect 474 4038 486 4041
rect 546 4038 638 4041
rect 666 4038 686 4041
rect 938 4038 990 4041
rect 1034 4038 1222 4041
rect 1522 4038 1574 4041
rect 1674 4038 1678 4041
rect 1862 4041 1865 4048
rect 2822 4042 2825 4048
rect 3310 4042 3313 4048
rect 3630 4042 3633 4048
rect 5054 4042 5057 4048
rect 1810 4038 1865 4041
rect 1982 4038 1990 4041
rect 1994 4038 2078 4041
rect 2090 4038 2102 4041
rect 2386 4038 2470 4041
rect 2474 4038 2734 4041
rect 3094 4038 3134 4041
rect 3154 4038 3246 4041
rect 3650 4038 3726 4041
rect 3730 4038 3910 4041
rect 3914 4038 3950 4041
rect 4010 4038 4174 4041
rect 4242 4038 4246 4041
rect 4466 4038 4854 4041
rect 5154 4038 5230 4041
rect 1294 4032 1297 4038
rect 2142 4032 2145 4038
rect 3094 4032 3097 4038
rect 50 4028 454 4031
rect 458 4028 510 4031
rect 570 4028 665 4031
rect 1538 4028 1686 4031
rect 1922 4028 2054 4031
rect 2834 4028 2854 4031
rect 2866 4028 2870 4031
rect 3338 4028 3526 4031
rect 3546 4028 3654 4031
rect 3730 4028 3854 4031
rect 3978 4028 4182 4031
rect 4338 4028 4830 4031
rect 4962 4028 5078 4031
rect 5138 4028 5193 4031
rect 662 4022 665 4028
rect 234 4018 398 4021
rect 410 4018 510 4021
rect 1514 4018 1662 4021
rect 1746 4018 2206 4021
rect 2414 4021 2417 4028
rect 5190 4022 5193 4028
rect 2218 4018 2417 4021
rect 2514 4018 2550 4021
rect 2778 4018 2822 4021
rect 2826 4018 2990 4021
rect 3122 4018 3494 4021
rect 3514 4018 3550 4021
rect 3602 4018 3678 4021
rect 3706 4018 4158 4021
rect 4162 4018 4294 4021
rect 4298 4018 4494 4021
rect 4746 4018 5182 4021
rect 66 4008 254 4011
rect 442 4008 494 4011
rect 506 4008 694 4011
rect 842 4008 1302 4011
rect 1378 4008 1590 4011
rect 1834 4008 1854 4011
rect 1858 4008 2078 4011
rect 2122 4008 2326 4011
rect 2514 4008 2734 4011
rect 2882 4008 3038 4011
rect 3042 4008 3358 4011
rect 3426 4008 3486 4011
rect 3490 4008 4054 4011
rect 4090 4008 4358 4011
rect 4850 4008 5094 4011
rect 5194 4008 5198 4011
rect 328 4003 330 4007
rect 334 4003 337 4007
rect 342 4003 344 4007
rect 1352 4003 1354 4007
rect 1358 4003 1361 4007
rect 1366 4003 1368 4007
rect 2384 4003 2386 4007
rect 2390 4003 2393 4007
rect 2398 4003 2400 4007
rect 3400 4003 3402 4007
rect 3406 4003 3409 4007
rect 3414 4003 3416 4007
rect 4424 4003 4426 4007
rect 4430 4003 4433 4007
rect 4438 4003 4440 4007
rect 90 3998 134 4001
rect 178 3998 238 4001
rect 290 3998 318 4001
rect 354 3998 638 4001
rect 1082 3998 1286 4001
rect 1810 3998 1838 4001
rect 1850 3998 1854 4001
rect 1858 3998 1974 4001
rect 2082 3998 2206 4001
rect 3306 3998 3374 4001
rect 3474 3998 4246 4001
rect 4354 3998 4358 4001
rect 5110 3992 5113 3998
rect 26 3988 142 3991
rect 330 3988 406 3991
rect 418 3988 518 3991
rect 606 3988 614 3991
rect 618 3988 646 3991
rect 1002 3988 1150 3991
rect 1282 3988 1310 3991
rect 1314 3988 1702 3991
rect 1714 3988 1942 3991
rect 1970 3988 2006 3991
rect 2010 3988 2094 3991
rect 2314 3988 2478 3991
rect 3226 3988 3342 3991
rect 3378 3988 3526 3991
rect 3530 3988 3574 3991
rect 3618 3988 3622 3991
rect 3802 3988 4094 3991
rect 4346 3988 4654 3991
rect 4658 3988 4822 3991
rect 5130 3988 5134 3991
rect 82 3978 86 3981
rect 90 3978 174 3981
rect 206 3981 209 3988
rect 206 3978 222 3981
rect 378 3978 494 3981
rect 498 3978 526 3981
rect 594 3978 598 3981
rect 626 3978 702 3981
rect 730 3978 854 3981
rect 1350 3978 1462 3981
rect 1506 3978 1694 3981
rect 1698 3978 1750 3981
rect 1766 3978 1926 3981
rect 1962 3978 2134 3981
rect 2378 3978 2582 3981
rect 3010 3978 3102 3981
rect 3146 3978 3214 3981
rect 3434 3978 4046 3981
rect 4306 3978 4726 3981
rect 4730 3978 4870 3981
rect 582 3972 585 3978
rect 10 3968 38 3971
rect 42 3968 350 3971
rect 370 3968 414 3971
rect 454 3968 462 3971
rect 466 3968 558 3971
rect 562 3968 574 3971
rect 586 3968 678 3971
rect 706 3968 734 3971
rect 1062 3971 1065 3978
rect 1050 3968 1065 3971
rect 1286 3971 1289 3978
rect 1226 3968 1289 3971
rect 1350 3972 1353 3978
rect 1666 3968 1694 3971
rect 1766 3971 1769 3978
rect 1706 3968 1769 3971
rect 1778 3968 2126 3971
rect 2138 3968 2198 3971
rect 2334 3971 2337 3978
rect 2298 3968 2337 3971
rect 2426 3968 2494 3971
rect 2650 3968 2750 3971
rect 2754 3968 2846 3971
rect 2942 3971 2945 3978
rect 2942 3968 3249 3971
rect 3326 3971 3329 3978
rect 3290 3968 3329 3971
rect 3562 3968 3574 3971
rect 3682 3968 3830 3971
rect 4042 3968 4118 3971
rect 4374 3968 4518 3971
rect 4754 3968 4758 3971
rect 4794 3968 4825 3971
rect 42 3958 126 3961
rect 146 3958 150 3961
rect 202 3958 230 3961
rect 282 3958 294 3961
rect 314 3958 318 3961
rect 322 3958 358 3961
rect 450 3958 462 3961
rect 550 3958 958 3961
rect 962 3958 1094 3961
rect 1114 3958 1374 3961
rect 1378 3958 1502 3961
rect 1658 3958 2118 3961
rect 2138 3958 2190 3961
rect 2222 3961 2225 3968
rect 2222 3958 2321 3961
rect 2330 3958 2334 3961
rect 2534 3961 2537 3968
rect 2490 3958 2537 3961
rect 2626 3958 2710 3961
rect 2770 3958 2830 3961
rect 2954 3958 3150 3961
rect 3246 3961 3249 3968
rect 3246 3958 3390 3961
rect 3394 3958 3430 3961
rect 3622 3961 3625 3968
rect 4374 3962 4377 3968
rect 4822 3962 4825 3968
rect 5014 3968 5102 3971
rect 3610 3958 3625 3961
rect 3718 3958 3726 3961
rect 3730 3958 3782 3961
rect 3866 3958 3966 3961
rect 4130 3958 4254 3961
rect 4346 3958 4350 3961
rect 4490 3958 4494 3961
rect 4730 3958 4806 3961
rect 4826 3958 4854 3961
rect 4914 3958 4918 3961
rect 4998 3961 5001 3968
rect 4994 3958 5001 3961
rect 5014 3962 5017 3968
rect 5022 3958 5038 3961
rect 5122 3958 5142 3961
rect 5162 3958 5174 3961
rect 550 3952 553 3958
rect 158 3948 222 3951
rect 306 3948 374 3951
rect 394 3948 502 3951
rect 506 3948 550 3951
rect 562 3948 582 3951
rect 906 3948 982 3951
rect 1010 3948 1054 3951
rect 1130 3948 1230 3951
rect 1290 3948 1294 3951
rect 1338 3948 1414 3951
rect 1418 3948 1486 3951
rect 1490 3948 1510 3951
rect 1666 3948 1670 3951
rect 1674 3948 1758 3951
rect 1802 3948 1870 3951
rect 1898 3948 1902 3951
rect 2010 3948 2014 3951
rect 2042 3948 2046 3951
rect 2126 3951 2129 3958
rect 2090 3948 2129 3951
rect 2138 3948 2158 3951
rect 2170 3948 2174 3951
rect 2186 3948 2230 3951
rect 2318 3951 2321 3958
rect 3182 3952 3185 3958
rect 3502 3952 3505 3958
rect 3638 3952 3641 3958
rect 2318 3948 2398 3951
rect 2442 3948 2694 3951
rect 2786 3948 2806 3951
rect 2810 3948 2838 3951
rect 2858 3948 2862 3951
rect 2882 3948 2918 3951
rect 3074 3948 3086 3951
rect 3130 3948 3158 3951
rect 3378 3948 3382 3951
rect 3490 3948 3494 3951
rect 3510 3948 3518 3951
rect 3522 3948 3614 3951
rect 3650 3948 3718 3951
rect 3722 3948 3726 3951
rect 3794 3948 3910 3951
rect 3914 3948 3934 3951
rect 3954 3948 3966 3951
rect 4078 3948 4086 3951
rect 4110 3951 4113 3958
rect 4110 3948 4222 3951
rect 4274 3948 4286 3951
rect 4446 3948 4478 3951
rect 4506 3948 4510 3951
rect 4610 3948 4614 3951
rect 4746 3948 4806 3951
rect 4890 3948 4894 3951
rect 4914 3948 4950 3951
rect 4986 3948 4990 3951
rect 5002 3948 5006 3951
rect 5022 3951 5025 3958
rect 5018 3948 5025 3951
rect 5050 3948 5054 3951
rect 62 3941 65 3948
rect 158 3942 161 3948
rect 390 3942 393 3948
rect 734 3942 737 3948
rect 62 3938 70 3941
rect 258 3938 286 3941
rect 378 3938 382 3941
rect 410 3938 430 3941
rect 474 3938 574 3941
rect 578 3938 606 3941
rect 754 3938 774 3941
rect 798 3941 801 3948
rect 1790 3942 1793 3948
rect 1942 3942 1945 3948
rect 2430 3942 2433 3948
rect 2878 3942 2881 3948
rect 778 3938 838 3941
rect 970 3938 1030 3941
rect 1034 3938 1374 3941
rect 1402 3938 1542 3941
rect 1602 3938 1686 3941
rect 1810 3938 1934 3941
rect 2018 3938 2022 3941
rect 2034 3938 2038 3941
rect 2058 3938 2206 3941
rect 2330 3938 2334 3941
rect 2506 3938 2534 3941
rect 2858 3938 2873 3941
rect 3050 3938 3110 3941
rect 3318 3941 3321 3948
rect 4022 3942 4025 3948
rect 4078 3942 4081 3948
rect 4446 3942 4449 3948
rect 3138 3938 3321 3941
rect 3386 3938 3390 3941
rect 3402 3938 3526 3941
rect 3530 3938 3566 3941
rect 3610 3938 3614 3941
rect 3642 3938 3654 3941
rect 3698 3938 3734 3941
rect 3922 3938 3990 3941
rect 4122 3938 4150 3941
rect 4274 3938 4310 3941
rect 4518 3941 4521 3948
rect 5122 3948 5158 3951
rect 4518 3938 4734 3941
rect 4810 3938 4894 3941
rect 4898 3938 4921 3941
rect 54 3931 57 3938
rect 198 3932 201 3938
rect 1750 3932 1753 3938
rect 54 3928 110 3931
rect 410 3928 454 3931
rect 458 3928 486 3931
rect 514 3928 646 3931
rect 754 3928 809 3931
rect 1018 3928 1054 3931
rect 1242 3928 1270 3931
rect 1274 3928 1278 3931
rect 1418 3928 1470 3931
rect 1490 3928 1510 3931
rect 1554 3928 1574 3931
rect 1674 3928 1742 3931
rect 1794 3928 1814 3931
rect 1818 3928 1822 3931
rect 1986 3928 1990 3931
rect 2090 3928 2182 3931
rect 2194 3928 2198 3931
rect 2246 3931 2249 3938
rect 2438 3932 2441 3938
rect 2246 3928 2358 3931
rect 2474 3928 2518 3931
rect 2582 3931 2585 3938
rect 2582 3928 2638 3931
rect 2798 3931 2801 3938
rect 2706 3928 2801 3931
rect 2870 3932 2873 3938
rect 2874 3928 3054 3931
rect 3234 3928 3286 3931
rect 3474 3928 3678 3931
rect 3730 3928 3734 3931
rect 3990 3931 3993 3938
rect 4918 3932 4921 3938
rect 5050 3938 5078 3941
rect 5170 3938 5190 3941
rect 4990 3932 4993 3938
rect 4998 3932 5001 3938
rect 3866 3928 3961 3931
rect 3990 3928 4014 3931
rect 4066 3928 4070 3931
rect 4122 3928 4302 3931
rect 4306 3928 4390 3931
rect 4554 3928 4606 3931
rect 4650 3928 4846 3931
rect 5150 3931 5153 3938
rect 5022 3928 5153 3931
rect 5270 3932 5273 3938
rect 6 3921 9 3928
rect 806 3922 809 3928
rect 1662 3922 1665 3928
rect 2230 3922 2233 3928
rect 3958 3922 3961 3928
rect 4958 3922 4961 3928
rect 5022 3922 5025 3928
rect 6 3918 62 3921
rect 226 3918 446 3921
rect 450 3918 478 3921
rect 530 3918 638 3921
rect 658 3918 758 3921
rect 826 3918 870 3921
rect 962 3918 990 3921
rect 994 3918 1078 3921
rect 1114 3918 1134 3921
rect 1138 3918 1526 3921
rect 1722 3918 1918 3921
rect 2330 3918 2558 3921
rect 2570 3918 3198 3921
rect 3218 3918 3318 3921
rect 3458 3918 3494 3921
rect 3546 3918 3574 3921
rect 3658 3918 3750 3921
rect 4106 3918 4238 3921
rect 4306 3918 4326 3921
rect 4730 3918 4790 3921
rect 4794 3918 4958 3921
rect 66 3908 198 3911
rect 306 3908 326 3911
rect 434 3908 542 3911
rect 570 3908 686 3911
rect 690 3908 838 3911
rect 922 3908 1022 3911
rect 1026 3908 1142 3911
rect 1154 3908 1174 3911
rect 1218 3908 1222 3911
rect 1250 3908 1390 3911
rect 1738 3908 1806 3911
rect 2330 3908 2566 3911
rect 2594 3908 2638 3911
rect 2642 3908 2718 3911
rect 2730 3908 2742 3911
rect 2930 3908 3126 3911
rect 3198 3911 3201 3918
rect 3582 3912 3585 3918
rect 3198 3908 3462 3911
rect 3466 3908 3566 3911
rect 3978 3908 4126 3911
rect 4138 3908 4142 3911
rect 4170 3908 4230 3911
rect 4234 3908 4446 3911
rect 4538 3908 4542 3911
rect 4626 3908 4894 3911
rect 848 3903 850 3907
rect 854 3903 857 3907
rect 862 3903 864 3907
rect 1872 3903 1874 3907
rect 1878 3903 1881 3907
rect 1886 3903 1888 3907
rect 2888 3903 2890 3907
rect 2894 3903 2897 3907
rect 2902 3903 2904 3907
rect 3920 3903 3922 3907
rect 3926 3903 3929 3907
rect 3934 3903 3936 3907
rect 4502 3902 4505 3908
rect 4936 3903 4938 3907
rect 4942 3903 4945 3907
rect 4950 3903 4952 3907
rect 58 3898 182 3901
rect 514 3898 790 3901
rect 794 3898 841 3901
rect 874 3898 990 3901
rect 1210 3898 1334 3901
rect 1442 3898 1454 3901
rect 1458 3898 1718 3901
rect 1754 3898 1790 3901
rect 1794 3898 1822 3901
rect 2366 3898 2574 3901
rect 2578 3898 2830 3901
rect 2978 3898 3262 3901
rect 3322 3898 3366 3901
rect 3378 3898 3382 3901
rect 3578 3898 3590 3901
rect 3618 3898 3670 3901
rect 3674 3898 3694 3901
rect 3946 3898 4030 3901
rect 4338 3898 4398 3901
rect 4538 3898 4590 3901
rect 5002 3898 5118 3901
rect 154 3888 166 3891
rect 170 3888 174 3891
rect 378 3888 550 3891
rect 634 3888 766 3891
rect 838 3891 841 3898
rect 838 3888 918 3891
rect 938 3888 969 3891
rect 1178 3888 1830 3891
rect 1890 3888 2134 3891
rect 2170 3888 2286 3891
rect 2322 3888 2334 3891
rect 2366 3891 2369 3898
rect 2338 3888 2369 3891
rect 2386 3888 2510 3891
rect 2514 3888 2614 3891
rect 2626 3888 2662 3891
rect 2826 3888 2974 3891
rect 3234 3888 3382 3891
rect 3398 3888 3406 3891
rect 3410 3888 3534 3891
rect 3586 3888 3622 3891
rect 3650 3888 3686 3891
rect 3690 3888 4593 3891
rect 966 3882 969 3888
rect 4590 3882 4593 3888
rect 4894 3888 4990 3891
rect 5042 3888 5142 3891
rect 5146 3888 5174 3891
rect 4894 3882 4897 3888
rect 122 3878 126 3881
rect 162 3878 230 3881
rect 354 3878 438 3881
rect 442 3878 486 3881
rect 490 3878 534 3881
rect 602 3878 710 3881
rect 874 3878 958 3881
rect 970 3878 974 3881
rect 1058 3878 1158 3881
rect 1178 3878 1182 3881
rect 1202 3878 1222 3881
rect 1234 3878 1238 3881
rect 1354 3878 1382 3881
rect 1426 3878 1486 3881
rect 1602 3878 1630 3881
rect 1634 3878 1662 3881
rect 1714 3878 1774 3881
rect 1778 3878 1782 3881
rect 2002 3878 2070 3881
rect 2226 3878 2278 3881
rect 2418 3878 2422 3881
rect 2442 3878 2486 3881
rect 2554 3878 2649 3881
rect 2746 3878 2838 3881
rect 2914 3878 2918 3881
rect 2922 3878 3094 3881
rect 3122 3878 3214 3881
rect 3282 3878 3542 3881
rect 3570 3878 3646 3881
rect 3650 3878 3686 3881
rect 3698 3878 3726 3881
rect 3874 3878 3966 3881
rect 3970 3878 3998 3881
rect 4034 3878 4302 3881
rect 4314 3878 4414 3881
rect 4426 3878 4454 3881
rect 4498 3878 4510 3881
rect 4594 3878 4609 3881
rect 5038 3881 5041 3888
rect 4922 3878 5041 3881
rect 18 3868 86 3871
rect 90 3868 190 3871
rect 194 3868 286 3871
rect 290 3868 366 3871
rect 574 3871 577 3878
rect 506 3868 577 3871
rect 762 3868 849 3871
rect 914 3868 934 3871
rect 938 3868 982 3871
rect 986 3868 1302 3871
rect 1322 3868 1326 3871
rect 1334 3871 1337 3878
rect 1814 3872 1817 3878
rect 2102 3872 2105 3878
rect 2646 3872 2649 3878
rect 1334 3868 1550 3871
rect 1826 3868 1830 3871
rect 1842 3868 1894 3871
rect 1922 3868 1926 3871
rect 2050 3868 2054 3871
rect 2138 3868 2150 3871
rect 2154 3868 2350 3871
rect 2354 3868 2406 3871
rect 2450 3868 2502 3871
rect 2506 3868 2574 3871
rect 2666 3868 2670 3871
rect 2682 3868 2686 3871
rect 2738 3868 2742 3871
rect 2846 3871 2849 3878
rect 2878 3871 2881 3878
rect 4606 3872 4609 3878
rect 5174 3872 5177 3878
rect 2846 3868 2881 3871
rect 2914 3868 2950 3871
rect 3122 3868 3126 3871
rect 3178 3868 3350 3871
rect 3354 3868 3430 3871
rect 3442 3868 3494 3871
rect 3498 3868 3526 3871
rect 3682 3868 3694 3871
rect 3802 3868 3862 3871
rect 3922 3868 4198 3871
rect 4202 3868 4206 3871
rect 4274 3868 4550 3871
rect 4554 3868 4574 3871
rect 4842 3868 4862 3871
rect 4866 3868 4998 3871
rect 846 3862 849 3868
rect 122 3858 126 3861
rect 130 3858 262 3861
rect 362 3858 382 3861
rect 938 3858 942 3861
rect 1002 3858 1006 3861
rect 1066 3858 1070 3861
rect 1186 3858 1209 3861
rect 1226 3858 1262 3861
rect 1306 3858 1310 3861
rect 1314 3858 1366 3861
rect 1378 3858 1382 3861
rect 1402 3858 1462 3861
rect 1554 3858 1630 3861
rect 1698 3858 1726 3861
rect 1758 3861 1761 3868
rect 2086 3862 2089 3868
rect 1746 3858 1761 3861
rect 1810 3858 1894 3861
rect 1906 3858 1942 3861
rect 2010 3858 2014 3861
rect 2106 3858 2150 3861
rect 2254 3858 2270 3861
rect 2414 3861 2417 3868
rect 2386 3858 2417 3861
rect 2574 3861 2577 3868
rect 2574 3858 2598 3861
rect 2674 3858 2838 3861
rect 2850 3858 2854 3861
rect 2878 3861 2881 3868
rect 5030 3862 5033 3868
rect 2878 3858 2918 3861
rect 2978 3858 3046 3861
rect 3074 3858 3134 3861
rect 3154 3858 3222 3861
rect 3306 3858 3310 3861
rect 3362 3858 3630 3861
rect 3634 3858 3646 3861
rect 3746 3858 3854 3861
rect 4114 3858 4126 3861
rect 4162 3858 4246 3861
rect 4338 3858 4342 3861
rect 4394 3858 4430 3861
rect 4458 3858 4462 3861
rect 4466 3858 4486 3861
rect 4754 3858 4790 3861
rect 5118 3861 5121 3868
rect 5118 3858 5150 3861
rect 5170 3858 5174 3861
rect 5194 3858 5198 3861
rect 5250 3858 5254 3861
rect 114 3848 206 3851
rect 218 3848 222 3851
rect 266 3848 374 3851
rect 418 3848 446 3851
rect 450 3848 494 3851
rect 498 3848 518 3851
rect 522 3848 702 3851
rect 934 3851 937 3858
rect 706 3848 937 3851
rect 1046 3851 1049 3858
rect 1086 3852 1089 3858
rect 1094 3852 1097 3858
rect 1206 3852 1209 3858
rect 2038 3852 2041 3858
rect 2254 3852 2257 3858
rect 3070 3852 3073 3858
rect 3718 3852 3721 3858
rect 3886 3852 3889 3858
rect 1010 3848 1049 3851
rect 1058 3848 1078 3851
rect 1258 3848 1398 3851
rect 1610 3848 1646 3851
rect 1650 3848 1798 3851
rect 1834 3848 1838 3851
rect 1930 3848 1950 3851
rect 1954 3848 1990 3851
rect 2066 3848 2070 3851
rect 2082 3848 2110 3851
rect 2154 3848 2214 3851
rect 2266 3848 2302 3851
rect 2306 3848 2342 3851
rect 2346 3848 2358 3851
rect 2378 3848 2574 3851
rect 2630 3848 2649 3851
rect 2810 3848 2862 3851
rect 2926 3848 2934 3851
rect 3106 3848 3182 3851
rect 3378 3848 3382 3851
rect 3498 3848 3542 3851
rect 3586 3848 3590 3851
rect 3810 3848 3814 3851
rect 3862 3848 3870 3851
rect 4122 3848 4222 3851
rect 4298 3848 4318 3851
rect 4370 3848 4374 3851
rect 4386 3848 4526 3851
rect 4846 3851 4849 3858
rect 4894 3852 4897 3858
rect 4982 3852 4985 3858
rect 4846 3848 4870 3851
rect 4874 3848 4886 3851
rect 5042 3848 5166 3851
rect 2630 3842 2633 3848
rect 2646 3842 2649 3848
rect 2926 3842 2929 3848
rect 3862 3842 3865 3848
rect 26 3838 38 3841
rect 42 3838 78 3841
rect 82 3838 94 3841
rect 106 3838 126 3841
rect 138 3838 262 3841
rect 314 3838 374 3841
rect 378 3838 446 3841
rect 474 3838 478 3841
rect 1034 3838 1038 3841
rect 1042 3838 1878 3841
rect 1882 3838 2006 3841
rect 2250 3838 2446 3841
rect 2490 3838 2566 3841
rect 2714 3838 2870 3841
rect 3098 3838 3294 3841
rect 3298 3838 3446 3841
rect 3498 3838 3734 3841
rect 3754 3838 3846 3841
rect 3978 3838 4894 3841
rect 5138 3838 5150 3841
rect 5154 3838 5222 3841
rect 74 3828 102 3831
rect 130 3828 238 3831
rect 242 3828 278 3831
rect 282 3828 350 3831
rect 354 3828 382 3831
rect 466 3828 702 3831
rect 1018 3828 1422 3831
rect 1498 3828 1678 3831
rect 1834 3828 1854 3831
rect 2098 3828 2438 3831
rect 3038 3831 3041 3838
rect 3038 3828 3182 3831
rect 3218 3828 3366 3831
rect 3370 3828 3462 3831
rect 3706 3828 3782 3831
rect 3786 3828 3806 3831
rect 4018 3828 4094 3831
rect 4098 3828 4158 3831
rect 4282 3828 4374 3831
rect 4378 3828 4494 3831
rect 4498 3828 4678 3831
rect 4682 3828 4734 3831
rect 4754 3828 4865 3831
rect 102 3822 105 3828
rect 226 3818 310 3821
rect 370 3818 390 3821
rect 474 3818 478 3821
rect 1222 3818 1230 3821
rect 1446 3821 1449 3828
rect 4862 3822 4865 3828
rect 1234 3818 1449 3821
rect 1458 3818 1638 3821
rect 1642 3818 1942 3821
rect 1946 3818 2126 3821
rect 2346 3818 2670 3821
rect 2722 3818 3070 3821
rect 3274 3818 3598 3821
rect 3602 3818 3686 3821
rect 4066 3818 4110 3821
rect 4114 3818 4230 3821
rect 4258 3818 4854 3821
rect 4998 3821 5001 3828
rect 4874 3818 5001 3821
rect 5126 3812 5129 3818
rect 74 3808 126 3811
rect 282 3808 318 3811
rect 1474 3808 1646 3811
rect 1770 3808 1966 3811
rect 2114 3808 2294 3811
rect 2506 3808 2582 3811
rect 3282 3808 3342 3811
rect 3466 3808 3710 3811
rect 4002 3808 4302 3811
rect 4826 3808 4910 3811
rect 328 3803 330 3807
rect 334 3803 337 3807
rect 342 3803 344 3807
rect 1352 3803 1354 3807
rect 1358 3803 1361 3807
rect 1366 3803 1368 3807
rect 1694 3802 1697 3808
rect 2384 3803 2386 3807
rect 2390 3803 2393 3807
rect 2398 3803 2400 3807
rect 3086 3802 3089 3808
rect 3400 3803 3402 3807
rect 3406 3803 3409 3807
rect 3414 3803 3416 3807
rect 4424 3803 4426 3807
rect 4430 3803 4433 3807
rect 4438 3803 4440 3807
rect 210 3798 310 3801
rect 1018 3798 1022 3801
rect 1106 3798 1174 3801
rect 1450 3798 1534 3801
rect 1546 3798 1694 3801
rect 1914 3798 2094 3801
rect 2178 3798 2366 3801
rect 2506 3798 2510 3801
rect 3506 3798 3526 3801
rect 3858 3798 3958 3801
rect 3962 3798 4006 3801
rect 4010 3798 4342 3801
rect 4346 3798 4358 3801
rect 4722 3798 4958 3801
rect 4978 3798 5014 3801
rect 5114 3798 5118 3801
rect 250 3788 422 3791
rect 1218 3788 1446 3791
rect 1458 3788 1574 3791
rect 1586 3788 1790 3791
rect 2034 3788 2182 3791
rect 2402 3788 2766 3791
rect 2770 3788 2878 3791
rect 2986 3788 3086 3791
rect 3154 3788 3206 3791
rect 3634 3788 3662 3791
rect 3858 3788 3982 3791
rect 4114 3788 4134 3791
rect 4370 3788 4510 3791
rect 4794 3788 4822 3791
rect 4858 3788 5054 3791
rect 5110 3788 5150 3791
rect -26 3781 -22 3782
rect -26 3778 30 3781
rect 34 3778 118 3781
rect 122 3778 158 3781
rect 162 3778 278 3781
rect 1146 3778 1374 3781
rect 1378 3778 1502 3781
rect 1562 3778 1702 3781
rect 1914 3778 2022 3781
rect 2114 3778 2158 3781
rect 2394 3778 2806 3781
rect 2810 3778 3094 3781
rect 3138 3778 3262 3781
rect 3266 3778 3398 3781
rect 3442 3778 3446 3781
rect 3450 3778 3526 3781
rect 3730 3778 3750 3781
rect 3898 3778 3926 3781
rect 3930 3778 3950 3781
rect 3986 3778 4038 3781
rect 4174 3781 4177 3788
rect 5110 3782 5113 3788
rect 4138 3778 4177 3781
rect 4202 3778 4542 3781
rect 4654 3778 4990 3781
rect 5058 3778 5094 3781
rect 42 3768 46 3771
rect 66 3768 78 3771
rect 90 3768 102 3771
rect 106 3768 113 3771
rect 130 3768 134 3771
rect 410 3768 446 3771
rect 642 3768 646 3771
rect 1162 3768 1206 3771
rect 1242 3768 1414 3771
rect 1426 3768 1438 3771
rect 1478 3768 1486 3771
rect 1490 3768 1518 3771
rect 1854 3771 1857 3778
rect 4654 3772 4657 3778
rect 1818 3768 1857 3771
rect 1938 3768 2126 3771
rect 2362 3768 2702 3771
rect 2798 3768 2806 3771
rect 2810 3768 2822 3771
rect 2842 3768 3046 3771
rect 3122 3768 3758 3771
rect 3778 3768 4174 3771
rect 4178 3768 4382 3771
rect 4386 3768 4398 3771
rect 4418 3768 4542 3771
rect 4634 3768 4654 3771
rect 4706 3768 4742 3771
rect 4914 3768 4942 3771
rect 4998 3771 5001 3778
rect 4946 3768 5001 3771
rect 5082 3768 5110 3771
rect 5114 3768 5118 3771
rect -26 3761 -22 3762
rect -26 3758 86 3761
rect 90 3758 134 3761
rect 254 3761 257 3768
rect 3030 3762 3033 3768
rect 210 3758 257 3761
rect 282 3758 310 3761
rect 314 3758 1150 3761
rect 1154 3758 1886 3761
rect 1994 3758 2222 3761
rect 2306 3758 2310 3761
rect 2338 3758 2438 3761
rect 2442 3758 2478 3761
rect 2482 3758 2526 3761
rect 2634 3758 2670 3761
rect 2698 3758 3022 3761
rect 3042 3758 3046 3761
rect 3146 3758 3150 3761
rect 3174 3758 3190 3761
rect 3230 3758 3262 3761
rect 3290 3758 3462 3761
rect 3474 3758 3478 3761
rect 3562 3758 3718 3761
rect 3834 3758 3910 3761
rect 3994 3758 3998 3761
rect 4010 3758 4022 3761
rect 4058 3758 4270 3761
rect 4330 3758 4334 3761
rect 4362 3758 4406 3761
rect 4546 3758 4614 3761
rect 4626 3758 4630 3761
rect 4798 3761 4801 3768
rect 4730 3758 4801 3761
rect 4842 3758 4926 3761
rect 4994 3758 5110 3761
rect 5158 3761 5161 3768
rect 5138 3758 5161 3761
rect 1934 3752 1937 3758
rect 50 3748 54 3751
rect 82 3748 86 3751
rect 98 3748 102 3751
rect 234 3748 358 3751
rect 402 3748 414 3751
rect 786 3748 846 3751
rect 854 3748 886 3751
rect 934 3748 977 3751
rect 1162 3748 1222 3751
rect 1306 3748 1470 3751
rect 1506 3748 1510 3751
rect 1602 3748 1606 3751
rect 1730 3748 1734 3751
rect 1754 3748 1878 3751
rect 1958 3751 1961 3758
rect 3174 3752 3177 3758
rect 3230 3752 3233 3758
rect 1958 3748 1982 3751
rect 2122 3748 2142 3751
rect 2162 3748 2361 3751
rect 2410 3748 2502 3751
rect 2626 3748 2662 3751
rect 2698 3748 2721 3751
rect 2730 3748 2742 3751
rect 2786 3748 2790 3751
rect 2834 3748 2918 3751
rect 2954 3748 2982 3751
rect 3010 3748 3174 3751
rect 3218 3748 3222 3751
rect 3394 3748 3486 3751
rect 3610 3748 3662 3751
rect 3718 3751 3721 3758
rect 3718 3748 3894 3751
rect 3898 3748 4070 3751
rect 4210 3748 4374 3751
rect 4410 3748 4462 3751
rect 4498 3748 4545 3751
rect 4626 3748 4630 3751
rect 4750 3748 4766 3751
rect 4850 3748 4865 3751
rect 4906 3748 4918 3751
rect 4922 3748 4926 3751
rect 4994 3748 5126 3751
rect 5130 3748 5270 3751
rect 5274 3748 5294 3751
rect 106 3738 110 3741
rect 154 3738 217 3741
rect 266 3738 294 3741
rect 298 3738 318 3741
rect 394 3738 510 3741
rect 550 3741 553 3748
rect 566 3741 569 3748
rect 662 3741 665 3748
rect 758 3741 761 3748
rect 550 3738 761 3741
rect 854 3741 857 3748
rect 934 3742 937 3748
rect 974 3742 977 3748
rect 1614 3742 1617 3748
rect 794 3738 857 3741
rect 882 3738 910 3741
rect 1098 3738 1166 3741
rect 1194 3738 1230 3741
rect 1250 3738 1254 3741
rect 1314 3738 1390 3741
rect 1418 3738 1478 3741
rect 1482 3738 1582 3741
rect 1642 3738 1646 3741
rect 1670 3741 1673 3748
rect 1670 3738 1686 3741
rect 1698 3738 1742 3741
rect 1746 3738 1902 3741
rect 1954 3738 1966 3741
rect 1982 3738 1990 3741
rect 1994 3738 2038 3741
rect 2086 3741 2089 3748
rect 2358 3742 2361 3748
rect 2082 3738 2089 3741
rect 2114 3738 2246 3741
rect 2290 3738 2318 3741
rect 2442 3738 2446 3741
rect 2498 3738 2502 3741
rect 2506 3738 2558 3741
rect 2586 3738 2638 3741
rect 2642 3738 2686 3741
rect 2706 3738 2710 3741
rect 2718 3741 2721 3748
rect 3366 3742 3369 3748
rect 3382 3742 3385 3748
rect 4542 3742 4545 3748
rect 4750 3742 4753 3748
rect 4862 3742 4865 3748
rect 4982 3742 4985 3748
rect 2718 3738 2782 3741
rect 2786 3738 2798 3741
rect 2842 3738 3286 3741
rect 3330 3738 3358 3741
rect 3418 3738 3462 3741
rect 3466 3738 3526 3741
rect 3530 3738 4030 3741
rect 4106 3738 4374 3741
rect 4578 3738 4662 3741
rect 4762 3738 4838 3741
rect 5114 3738 5129 3741
rect 214 3732 217 3738
rect 878 3732 881 3738
rect 2486 3732 2489 3738
rect 5126 3732 5129 3738
rect 5182 3738 5190 3741
rect 5182 3732 5185 3738
rect 138 3728 198 3731
rect 218 3728 294 3731
rect 298 3728 398 3731
rect 434 3728 590 3731
rect 650 3728 678 3731
rect 922 3728 926 3731
rect 1122 3728 1302 3731
rect 1490 3728 1550 3731
rect 1630 3728 1638 3731
rect 1642 3728 1646 3731
rect 1738 3728 1934 3731
rect 1946 3728 1958 3731
rect 2026 3728 2126 3731
rect 2154 3728 2158 3731
rect 2282 3728 2310 3731
rect 2314 3728 2326 3731
rect 2346 3728 2350 3731
rect 2418 3728 2422 3731
rect 2666 3728 2782 3731
rect 2794 3728 2822 3731
rect 2826 3728 2862 3731
rect 2882 3728 2942 3731
rect 3002 3728 3134 3731
rect 3162 3728 3182 3731
rect 3274 3728 3294 3731
rect 3338 3728 3454 3731
rect 3514 3728 3726 3731
rect 3730 3728 3734 3731
rect 3770 3728 3918 3731
rect 3994 3728 3998 3731
rect 4338 3728 4350 3731
rect 4358 3728 4390 3731
rect 4650 3728 4678 3731
rect 4850 3728 4862 3731
rect 4866 3728 4918 3731
rect 4978 3728 5038 3731
rect 5222 3731 5225 3738
rect 5222 3728 5294 3731
rect 194 3718 462 3721
rect 850 3718 894 3721
rect 1486 3721 1489 3728
rect 1186 3718 1489 3721
rect 1554 3718 1662 3721
rect 1666 3718 1846 3721
rect 1850 3718 1950 3721
rect 2138 3718 2270 3721
rect 2338 3718 2814 3721
rect 2818 3718 2862 3721
rect 2974 3721 2977 3728
rect 3982 3722 3985 3728
rect 2946 3718 2977 3721
rect 2986 3718 3198 3721
rect 3202 3718 3974 3721
rect 4166 3721 4169 3728
rect 4166 3718 4182 3721
rect 4310 3721 4313 3728
rect 4358 3722 4361 3728
rect 4310 3718 4326 3721
rect 4418 3718 4502 3721
rect 4794 3718 4958 3721
rect 4978 3718 5014 3721
rect 5134 3721 5137 3728
rect 5134 3718 5142 3721
rect 5166 3712 5169 3718
rect 202 3708 326 3711
rect 330 3708 486 3711
rect 602 3708 686 3711
rect 890 3708 1110 3711
rect 1194 3708 1710 3711
rect 1954 3708 1990 3711
rect 2018 3708 2206 3711
rect 2214 3708 2494 3711
rect 2522 3708 2590 3711
rect 2658 3708 2694 3711
rect 2714 3708 2718 3711
rect 2930 3708 2966 3711
rect 2978 3708 3110 3711
rect 3210 3708 3494 3711
rect 3498 3708 3534 3711
rect 3546 3708 3550 3711
rect 3714 3708 3734 3711
rect 3898 3708 3902 3711
rect 3978 3708 3998 3711
rect 4010 3708 4014 3711
rect 4250 3708 4774 3711
rect 848 3703 850 3707
rect 854 3703 857 3707
rect 862 3703 864 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1886 3703 1888 3707
rect 42 3698 62 3701
rect 66 3698 142 3701
rect 146 3698 206 3701
rect 410 3698 446 3701
rect 930 3698 1110 3701
rect 1258 3698 1286 3701
rect 1290 3698 1398 3701
rect 1490 3698 1686 3701
rect 1898 3698 2030 3701
rect 2042 3698 2070 3701
rect 2082 3698 2094 3701
rect 2106 3698 2110 3701
rect 2214 3701 2217 3708
rect 2888 3703 2890 3707
rect 2894 3703 2897 3707
rect 2902 3703 2904 3707
rect 3920 3703 3922 3707
rect 3926 3703 3929 3707
rect 3934 3703 3936 3707
rect 4936 3703 4938 3707
rect 4942 3703 4945 3707
rect 4950 3703 4952 3707
rect 2122 3698 2217 3701
rect 2258 3698 2262 3701
rect 2378 3698 2462 3701
rect 2466 3698 2542 3701
rect 2554 3698 2566 3701
rect 2586 3698 2606 3701
rect 2658 3698 2726 3701
rect 2746 3698 2782 3701
rect 2818 3698 2846 3701
rect 2922 3698 2982 3701
rect 3002 3698 3254 3701
rect 3458 3698 3526 3701
rect 3762 3698 3782 3701
rect 3954 3698 4038 3701
rect 4194 3698 4206 3701
rect 4234 3698 4414 3701
rect 5130 3698 5134 3701
rect 5162 3698 5174 3701
rect 5250 3698 5294 3701
rect 482 3688 566 3691
rect 850 3688 958 3691
rect 962 3688 1030 3691
rect 1142 3688 1150 3691
rect 1154 3688 1353 3691
rect 1362 3688 1502 3691
rect 1602 3688 1662 3691
rect 1666 3688 1814 3691
rect 2002 3688 2110 3691
rect 2226 3688 2286 3691
rect 2402 3688 2414 3691
rect 2418 3688 2630 3691
rect 2650 3688 2654 3691
rect 2798 3688 2806 3691
rect 2810 3688 2966 3691
rect 3042 3688 3086 3691
rect 3090 3688 3097 3691
rect 3106 3688 3334 3691
rect 3378 3688 3502 3691
rect 3522 3688 3574 3691
rect 3602 3688 3790 3691
rect 3842 3688 3942 3691
rect 3970 3688 4006 3691
rect 4138 3688 4166 3691
rect 4218 3688 4358 3691
rect 4362 3688 4366 3691
rect 4450 3688 4534 3691
rect 4666 3688 4678 3691
rect 4682 3688 4710 3691
rect 4842 3688 4950 3691
rect 4962 3688 4990 3691
rect 5106 3688 5150 3691
rect 1350 3682 1353 3688
rect -26 3681 -22 3682
rect -26 3678 14 3681
rect 130 3678 190 3681
rect 194 3678 206 3681
rect 210 3678 398 3681
rect 402 3678 454 3681
rect 530 3678 590 3681
rect 674 3678 718 3681
rect 722 3678 742 3681
rect 750 3678 758 3681
rect 762 3678 878 3681
rect 962 3678 982 3681
rect 1018 3678 1110 3681
rect 1114 3678 1158 3681
rect 1250 3678 1310 3681
rect 1378 3678 1430 3681
rect 1570 3678 1718 3681
rect 1834 3678 1838 3681
rect 1918 3681 1921 3688
rect 2974 3682 2977 3688
rect 1866 3678 1921 3681
rect 1938 3678 2190 3681
rect 2210 3678 2414 3681
rect 2418 3678 2430 3681
rect 2442 3678 2526 3681
rect 2562 3678 2790 3681
rect 2794 3678 2814 3681
rect 2842 3678 2846 3681
rect 2994 3678 3022 3681
rect 3342 3681 3345 3688
rect 3034 3678 3502 3681
rect 3898 3678 4222 3681
rect 4266 3678 4318 3681
rect 4406 3681 4409 3688
rect 4406 3678 4542 3681
rect 4590 3681 4593 3688
rect 5278 3682 5281 3688
rect 4590 3678 5118 3681
rect 5122 3678 5142 3681
rect 5178 3678 5206 3681
rect 106 3668 118 3671
rect 178 3668 206 3671
rect 210 3668 246 3671
rect 250 3668 270 3671
rect 434 3668 446 3671
rect 450 3668 734 3671
rect 738 3668 774 3671
rect 850 3668 966 3671
rect 970 3668 998 3671
rect 1114 3668 1118 3671
rect 1210 3668 1214 3671
rect 1242 3668 1246 3671
rect 1274 3668 1302 3671
rect 1314 3668 1454 3671
rect 1478 3671 1481 3678
rect 1478 3668 1486 3671
rect 1490 3668 1502 3671
rect 1586 3668 1590 3671
rect 1750 3671 1753 3678
rect 1750 3668 1782 3671
rect 1786 3668 1894 3671
rect 1930 3668 2102 3671
rect 2106 3668 2158 3671
rect 2250 3668 2297 3671
rect 2418 3668 2598 3671
rect 2738 3668 2966 3671
rect 3018 3668 3030 3671
rect 3050 3668 3118 3671
rect 3138 3668 3166 3671
rect 3242 3668 3246 3671
rect 3274 3668 3278 3671
rect 3346 3668 3350 3671
rect 3426 3668 3454 3671
rect 3514 3668 3550 3671
rect 3578 3668 3638 3671
rect 3658 3668 3662 3671
rect 3778 3668 4158 3671
rect 4162 3668 4166 3671
rect 4194 3668 4302 3671
rect 4306 3668 4326 3671
rect 4330 3668 4358 3671
rect 4770 3668 4958 3671
rect 4962 3668 5182 3671
rect -26 3661 -22 3662
rect 6 3661 9 3668
rect -26 3658 38 3661
rect 66 3658 86 3661
rect 90 3658 166 3661
rect 170 3658 198 3661
rect 202 3658 254 3661
rect 394 3658 510 3661
rect 586 3658 606 3661
rect 610 3658 630 3661
rect 642 3658 654 3661
rect 702 3658 710 3661
rect 726 3658 750 3661
rect 762 3659 822 3661
rect 2294 3662 2297 3668
rect 3046 3662 3049 3668
rect 4630 3662 4633 3668
rect 762 3658 825 3659
rect 922 3658 974 3661
rect 978 3658 1406 3661
rect 1426 3658 1478 3661
rect 1482 3658 1510 3661
rect 1514 3658 1574 3661
rect 1594 3658 1614 3661
rect 1618 3658 1854 3661
rect 1994 3658 2022 3661
rect 2058 3658 2062 3661
rect 2114 3658 2150 3661
rect 2330 3658 2438 3661
rect 2450 3658 2486 3661
rect 2494 3658 2585 3661
rect 2634 3658 2686 3661
rect 2714 3658 2721 3661
rect 2762 3658 2769 3661
rect 2850 3658 2881 3661
rect 702 3652 705 3658
rect 726 3652 729 3658
rect 2494 3652 2497 3658
rect 18 3648 54 3651
rect 58 3648 78 3651
rect 82 3648 110 3651
rect 114 3648 150 3651
rect 514 3648 590 3651
rect 626 3648 630 3651
rect 946 3648 1006 3651
rect 1178 3648 1182 3651
rect 1242 3648 1246 3651
rect 1314 3648 1318 3651
rect 1378 3648 1438 3651
rect 1582 3648 1609 3651
rect 910 3641 913 3648
rect 1550 3642 1553 3648
rect 1582 3642 1585 3648
rect 1606 3642 1609 3648
rect 1622 3648 1726 3651
rect 1802 3648 1822 3651
rect 1826 3648 1902 3651
rect 1930 3648 2137 3651
rect 2234 3648 2422 3651
rect 2442 3648 2446 3651
rect 2538 3648 2574 3651
rect 2582 3651 2585 3658
rect 2766 3652 2769 3658
rect 2878 3652 2881 3658
rect 2946 3658 2950 3661
rect 2962 3658 2982 3661
rect 3034 3658 3038 3661
rect 3090 3658 3158 3661
rect 3242 3658 3310 3661
rect 3338 3658 3350 3661
rect 3370 3658 3470 3661
rect 3610 3658 3646 3661
rect 3706 3658 3838 3661
rect 3842 3658 4006 3661
rect 4010 3658 4054 3661
rect 4090 3658 4094 3661
rect 4098 3658 4182 3661
rect 4210 3658 4246 3661
rect 4314 3658 4342 3661
rect 4354 3658 4366 3661
rect 4394 3658 4398 3661
rect 4402 3658 4566 3661
rect 4778 3658 4830 3661
rect 4858 3658 4878 3661
rect 5034 3658 5038 3661
rect 5042 3658 5126 3661
rect 5202 3658 5294 3661
rect 2934 3652 2937 3658
rect 3214 3652 3217 3658
rect 3558 3652 3561 3658
rect 4278 3652 4281 3658
rect 4606 3652 4609 3658
rect 4910 3652 4913 3658
rect 2582 3648 2654 3651
rect 2702 3648 2753 3651
rect 2778 3648 2798 3651
rect 2906 3648 2929 3651
rect 2946 3648 2950 3651
rect 2978 3648 3206 3651
rect 3322 3648 3390 3651
rect 3618 3648 3774 3651
rect 3842 3648 4246 3651
rect 4250 3648 4254 3651
rect 4450 3648 4478 3651
rect 4666 3648 4774 3651
rect 4994 3648 5038 3651
rect 5082 3648 5110 3651
rect 5134 3648 5142 3651
rect 5146 3648 5206 3651
rect 1622 3642 1625 3648
rect 778 3638 950 3641
rect 970 3638 1094 3641
rect 1098 3638 1126 3641
rect 1130 3638 1150 3641
rect 1154 3638 1222 3641
rect 1226 3638 1494 3641
rect 1634 3638 1638 3641
rect 1902 3641 1905 3648
rect 1654 3638 1833 3641
rect 1902 3638 2126 3641
rect 2134 3641 2137 3648
rect 2702 3642 2705 3648
rect 2750 3642 2753 3648
rect 2846 3642 2849 3648
rect 2854 3642 2857 3648
rect 2926 3642 2929 3648
rect 2134 3638 2526 3641
rect 2642 3638 2678 3641
rect 2986 3638 3054 3641
rect 3194 3638 3318 3641
rect 3426 3638 3518 3641
rect 3530 3638 3534 3641
rect 3590 3641 3593 3648
rect 3590 3638 3782 3641
rect 3786 3638 3798 3641
rect 3906 3638 3966 3641
rect 3978 3638 4102 3641
rect 4158 3638 4166 3641
rect 4170 3638 4198 3641
rect 4210 3638 4254 3641
rect 4378 3638 4670 3641
rect 4674 3638 4686 3641
rect 4698 3638 4814 3641
rect 4890 3638 5030 3641
rect 5110 3638 5118 3641
rect 5122 3638 5142 3641
rect 5242 3638 5270 3641
rect 1654 3632 1657 3638
rect 666 3628 1126 3631
rect 1146 3628 1174 3631
rect 1186 3628 1366 3631
rect 1370 3628 1630 3631
rect 1666 3628 1694 3631
rect 1794 3628 1798 3631
rect 1830 3631 1833 3638
rect 1830 3628 2086 3631
rect 2274 3628 2342 3631
rect 2442 3628 2590 3631
rect 2610 3628 2662 3631
rect 2666 3628 2710 3631
rect 2714 3628 2718 3631
rect 2722 3628 2782 3631
rect 2786 3628 2918 3631
rect 2978 3628 3177 3631
rect 3330 3628 3622 3631
rect 3674 3628 3742 3631
rect 3914 3628 3990 3631
rect 4046 3628 4142 3631
rect 4226 3628 4270 3631
rect 4314 3628 4646 3631
rect 4930 3628 5054 3631
rect 266 3618 294 3621
rect 786 3618 806 3621
rect 990 3618 998 3621
rect 1002 3618 1046 3621
rect 1106 3618 1278 3621
rect 1418 3618 2102 3621
rect 2106 3618 2614 3621
rect 2618 3618 3166 3621
rect 3174 3621 3177 3628
rect 4046 3622 4049 3628
rect 3174 3618 3422 3621
rect 3482 3618 3598 3621
rect 4090 3618 4094 3621
rect 4886 3621 4889 3628
rect 4178 3618 4889 3621
rect 5050 3618 5150 3621
rect 294 3612 297 3618
rect 466 3608 590 3611
rect 594 3608 646 3611
rect 1170 3608 1334 3611
rect 1466 3608 1886 3611
rect 1978 3608 2358 3611
rect 2426 3608 2606 3611
rect 2730 3608 2734 3611
rect 2762 3608 2766 3611
rect 2818 3608 2934 3611
rect 3218 3608 3222 3611
rect 3642 3608 3822 3611
rect 3826 3608 4078 3611
rect 4138 3608 4414 3611
rect 4466 3608 4782 3611
rect 4786 3608 4982 3611
rect 328 3603 330 3607
rect 334 3603 337 3607
rect 342 3603 344 3607
rect 1352 3603 1354 3607
rect 1358 3603 1361 3607
rect 1366 3603 1368 3607
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2398 3603 2400 3607
rect 3400 3603 3402 3607
rect 3406 3603 3409 3607
rect 3414 3603 3416 3607
rect 4424 3603 4426 3607
rect 4430 3603 4433 3607
rect 4438 3603 4440 3607
rect 378 3598 926 3601
rect 930 3598 974 3601
rect 1058 3598 1190 3601
rect 1374 3598 1486 3601
rect 1634 3598 1686 3601
rect 2234 3598 2342 3601
rect 2538 3598 2686 3601
rect 2690 3598 2862 3601
rect 2874 3598 3246 3601
rect 3250 3598 3390 3601
rect 3426 3598 3590 3601
rect 3826 3598 4126 3601
rect 4634 3598 5166 3601
rect 514 3588 678 3591
rect 682 3588 798 3591
rect 826 3588 918 3591
rect 962 3588 1038 3591
rect 1162 3588 1214 3591
rect 1218 3588 1270 3591
rect 1374 3591 1377 3598
rect 1838 3592 1841 3598
rect 1346 3588 1377 3591
rect 1474 3588 1662 3591
rect 1738 3588 1790 3591
rect 2114 3588 2286 3591
rect 2330 3588 2454 3591
rect 2578 3588 2606 3591
rect 2746 3588 3054 3591
rect 3058 3588 3158 3591
rect 3194 3588 3326 3591
rect 3458 3588 3542 3591
rect 3554 3588 3574 3591
rect 3594 3588 3694 3591
rect 3994 3588 4310 3591
rect 4450 3588 4614 3591
rect 106 3578 206 3581
rect 210 3578 502 3581
rect 506 3578 630 3581
rect 634 3578 734 3581
rect 738 3578 870 3581
rect 874 3578 1014 3581
rect 1018 3578 1342 3581
rect 1346 3578 1670 3581
rect 1834 3578 2174 3581
rect 2178 3578 2254 3581
rect 2510 3581 2513 3588
rect 5006 3582 5009 3588
rect 2510 3578 2582 3581
rect 2586 3578 2598 3581
rect 2674 3578 2790 3581
rect 2842 3578 2878 3581
rect 3282 3578 3814 3581
rect 3990 3578 4054 3581
rect 4106 3578 4190 3581
rect 4570 3578 4646 3581
rect 370 3568 462 3571
rect 498 3568 542 3571
rect 770 3568 793 3571
rect 1018 3568 1094 3571
rect 1106 3568 1193 3571
rect 1450 3568 1502 3571
rect 1766 3571 1769 3578
rect 2478 3572 2481 3578
rect 1626 3568 1769 3571
rect 1842 3568 1998 3571
rect 2242 3568 2361 3571
rect 2506 3568 2542 3571
rect 2578 3568 2638 3571
rect 2830 3571 2833 3578
rect 2818 3568 2833 3571
rect 2850 3568 2966 3571
rect 2970 3568 3030 3571
rect 3058 3568 3118 3571
rect 3174 3571 3177 3578
rect 3990 3572 3993 3578
rect 3174 3568 3190 3571
rect 3434 3568 3678 3571
rect 4002 3568 4006 3571
rect 4186 3568 4345 3571
rect 4558 3571 4561 3578
rect 4402 3568 4561 3571
rect 4570 3568 4582 3571
rect 114 3558 150 3561
rect 162 3558 302 3561
rect 386 3558 406 3561
rect 426 3558 486 3561
rect 566 3561 569 3568
rect 790 3562 793 3568
rect 1190 3562 1193 3568
rect 566 3558 782 3561
rect 794 3558 822 3561
rect 1002 3558 1174 3561
rect 1218 3558 1230 3561
rect 1234 3558 1422 3561
rect 1530 3558 1670 3561
rect 1786 3558 1790 3561
rect 1986 3558 2030 3561
rect 2034 3558 2054 3561
rect 2138 3558 2166 3561
rect 2250 3558 2254 3561
rect 2282 3558 2326 3561
rect 2358 3561 2361 3568
rect 4014 3562 4017 3568
rect 2358 3558 2550 3561
rect 2578 3558 2598 3561
rect 2650 3558 2686 3561
rect 2730 3558 2830 3561
rect 2866 3558 2950 3561
rect 2954 3558 2974 3561
rect 3002 3558 3294 3561
rect 3466 3558 3470 3561
rect 3506 3558 3542 3561
rect 3706 3558 3710 3561
rect 3730 3558 3734 3561
rect 3754 3558 3758 3561
rect 3962 3558 3990 3561
rect 4022 3561 4025 3568
rect 4062 3562 4065 3568
rect 4022 3558 4030 3561
rect 4226 3558 4278 3561
rect 4330 3558 4334 3561
rect 4342 3561 4345 3568
rect 4342 3558 4494 3561
rect 4514 3558 4526 3561
rect 4534 3558 4582 3561
rect 4602 3558 4686 3561
rect 5006 3561 5009 3568
rect 5006 3558 5094 3561
rect 5162 3558 5174 3561
rect 5242 3558 5246 3561
rect 5274 3558 5286 3561
rect 70 3548 118 3551
rect 422 3551 425 3558
rect 830 3552 833 3558
rect 138 3548 425 3551
rect 442 3548 518 3551
rect 546 3548 606 3551
rect 626 3548 630 3551
rect 642 3548 662 3551
rect 714 3548 798 3551
rect 974 3551 977 3558
rect 1478 3552 1481 3558
rect 1526 3552 1529 3558
rect 898 3548 977 3551
rect 1050 3548 1054 3551
rect 1098 3548 1158 3551
rect 1242 3548 1478 3551
rect 1490 3548 1502 3551
rect 1538 3548 1574 3551
rect 1586 3548 1590 3551
rect 1606 3548 1614 3551
rect 1642 3548 1646 3551
rect 1658 3548 1662 3551
rect 1698 3548 1702 3551
rect 1770 3548 1774 3551
rect 1794 3548 1814 3551
rect 1826 3548 1854 3551
rect 1858 3548 1966 3551
rect 1978 3548 1998 3551
rect 2002 3548 2030 3551
rect 2066 3548 2094 3551
rect 2098 3548 2166 3551
rect 2226 3548 2254 3551
rect 2274 3548 2310 3551
rect 2350 3551 2353 3558
rect 2346 3548 2353 3551
rect 2362 3548 2510 3551
rect 2650 3548 2742 3551
rect 2826 3548 2902 3551
rect 70 3542 73 3548
rect 162 3538 262 3541
rect 314 3538 326 3541
rect 514 3538 526 3541
rect 530 3538 638 3541
rect 642 3538 830 3541
rect 834 3538 846 3541
rect 858 3538 862 3541
rect 890 3538 902 3541
rect 1018 3538 1022 3541
rect 1042 3538 1193 3541
rect 1274 3538 1278 3541
rect 1282 3538 1350 3541
rect 1354 3538 1446 3541
rect 1490 3538 1750 3541
rect 1770 3538 1790 3541
rect 1906 3538 1990 3541
rect 2018 3538 2062 3541
rect 2106 3538 2142 3541
rect 2206 3541 2209 3548
rect 2510 3542 2513 3548
rect 2590 3542 2593 3548
rect 3026 3548 3046 3551
rect 3122 3548 3182 3551
rect 3250 3548 3318 3551
rect 3326 3551 3329 3558
rect 3494 3552 3497 3558
rect 3326 3548 3358 3551
rect 3410 3548 3494 3551
rect 3530 3548 3534 3551
rect 3642 3548 3694 3551
rect 3698 3548 3774 3551
rect 3886 3551 3889 3558
rect 4158 3552 4161 3558
rect 4534 3552 4537 3558
rect 3818 3548 3889 3551
rect 3954 3548 4022 3551
rect 4066 3548 4070 3551
rect 4098 3548 4110 3551
rect 4178 3548 4190 3551
rect 4314 3548 4350 3551
rect 4402 3548 4478 3551
rect 4482 3548 4526 3551
rect 4554 3548 4606 3551
rect 4658 3548 4662 3551
rect 4666 3548 4734 3551
rect 4794 3548 4862 3551
rect 4970 3548 4974 3551
rect 5026 3548 5150 3551
rect 5154 3548 5281 3551
rect 2178 3538 2209 3541
rect 2326 3538 2406 3541
rect 2682 3538 2710 3541
rect 2818 3538 2878 3541
rect 2882 3538 2910 3541
rect 2962 3538 2966 3541
rect 3026 3538 3038 3541
rect 3042 3538 3150 3541
rect 3170 3538 3190 3541
rect 3194 3538 3230 3541
rect 3258 3538 3286 3541
rect 3290 3538 3478 3541
rect 3498 3538 3502 3541
rect 3534 3538 3542 3541
rect 3546 3538 3606 3541
rect 3658 3538 4206 3541
rect 4222 3541 4225 3548
rect 4366 3542 4369 3548
rect 4638 3542 4641 3548
rect 4926 3542 4929 3548
rect 5278 3542 5281 3548
rect 5294 3542 5297 3548
rect 4222 3538 4358 3541
rect 4386 3538 4414 3541
rect 4474 3538 4614 3541
rect 4642 3538 4734 3541
rect 4818 3538 4822 3541
rect 4930 3538 5161 3541
rect 5178 3538 5198 3541
rect 90 3528 174 3531
rect 210 3528 318 3531
rect 390 3531 393 3538
rect 390 3528 462 3531
rect 482 3528 550 3531
rect 562 3528 566 3531
rect 594 3528 766 3531
rect 774 3528 910 3531
rect 1178 3528 1182 3531
rect 1190 3531 1193 3538
rect 2150 3532 2153 3538
rect 2326 3532 2329 3538
rect 5158 3532 5161 3538
rect 1190 3528 1294 3531
rect 1394 3528 1454 3531
rect 1498 3528 1566 3531
rect 1578 3528 1590 3531
rect 1626 3528 1630 3531
rect 1690 3528 1750 3531
rect 1754 3528 1758 3531
rect 1874 3528 2030 3531
rect 2042 3528 2049 3531
rect 2058 3528 2110 3531
rect 2354 3528 2358 3531
rect 2778 3528 2854 3531
rect 2866 3528 3254 3531
rect 3258 3528 3382 3531
rect 3442 3528 3446 3531
rect 3698 3528 3718 3531
rect 3722 3528 3806 3531
rect 3946 3528 3974 3531
rect 4026 3528 4030 3531
rect 4050 3528 4070 3531
rect 4194 3528 4214 3531
rect 4290 3528 4318 3531
rect 4386 3528 4390 3531
rect 4482 3528 4494 3531
rect 4506 3528 4942 3531
rect 4978 3528 5006 3531
rect 5010 3528 5038 3531
rect 5282 3528 5294 3531
rect 18 3518 102 3521
rect 266 3518 342 3521
rect 658 3518 662 3521
rect 774 3521 777 3528
rect 770 3518 777 3521
rect 874 3518 1038 3521
rect 1290 3518 1454 3521
rect 1538 3518 1545 3521
rect 1562 3518 1574 3521
rect 1870 3521 1873 3528
rect 1578 3518 1873 3521
rect 2046 3522 2049 3528
rect 2870 3522 2873 3528
rect 3678 3522 3681 3528
rect 4158 3522 4161 3528
rect 2090 3518 2126 3521
rect 2194 3518 2206 3521
rect 2306 3518 2374 3521
rect 2450 3518 2534 3521
rect 3002 3518 3094 3521
rect 3162 3518 3198 3521
rect 3210 3518 3214 3521
rect 3226 3518 3310 3521
rect 3322 3518 3430 3521
rect 3434 3518 3441 3521
rect 3450 3518 3670 3521
rect 3690 3518 3766 3521
rect 3994 3518 4094 3521
rect 4334 3521 4337 3528
rect 4210 3518 4337 3521
rect 4346 3518 4398 3521
rect 4498 3518 4574 3521
rect 4578 3518 4910 3521
rect 4914 3518 5046 3521
rect 5050 3518 5134 3521
rect 5194 3518 5198 3521
rect 5250 3518 5302 3521
rect 226 3508 638 3511
rect 906 3508 1006 3511
rect 1282 3508 1310 3511
rect 1338 3508 1366 3511
rect 1434 3508 1438 3511
rect 1450 3508 1542 3511
rect 1562 3508 1606 3511
rect 1618 3508 1622 3511
rect 1754 3508 1774 3511
rect 1778 3508 1806 3511
rect 1810 3508 1830 3511
rect 2034 3508 2086 3511
rect 2090 3508 2278 3511
rect 2330 3508 2334 3511
rect 2834 3508 2862 3511
rect 2914 3508 3262 3511
rect 3314 3508 3430 3511
rect 3686 3511 3689 3518
rect 3434 3508 3689 3511
rect 3970 3508 4214 3511
rect 4298 3508 4318 3511
rect 4322 3508 4510 3511
rect 4562 3508 4702 3511
rect 4850 3508 4910 3511
rect 5234 3508 5246 3511
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 862 3503 864 3507
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1886 3503 1888 3507
rect 2888 3503 2890 3507
rect 2894 3503 2897 3507
rect 2902 3503 2904 3507
rect 3920 3503 3922 3507
rect 3926 3503 3929 3507
rect 3934 3503 3936 3507
rect 4936 3503 4938 3507
rect 4942 3503 4945 3507
rect 4950 3503 4952 3507
rect 250 3498 390 3501
rect 394 3498 454 3501
rect 882 3498 966 3501
rect 1074 3498 1577 3501
rect 1586 3498 1710 3501
rect 1922 3498 2062 3501
rect 2218 3498 2230 3501
rect 2298 3498 2334 3501
rect 2338 3498 2766 3501
rect 2794 3498 2881 3501
rect 3210 3498 3214 3501
rect 3218 3498 3278 3501
rect 3282 3498 3502 3501
rect 3522 3498 3606 3501
rect 3610 3498 3630 3501
rect 3962 3498 4118 3501
rect 4146 3498 4310 3501
rect 4474 3498 4518 3501
rect 4522 3498 4590 3501
rect 4594 3498 4646 3501
rect 4978 3498 5214 3501
rect 330 3488 398 3491
rect 450 3488 542 3491
rect 826 3488 870 3491
rect 946 3488 1062 3491
rect 1094 3488 1190 3491
rect 1194 3488 1302 3491
rect 1338 3488 1414 3491
rect 1426 3488 1470 3491
rect 1502 3488 1510 3491
rect 1514 3488 1526 3491
rect 1574 3491 1577 3498
rect 1574 3488 1598 3491
rect 1610 3488 1718 3491
rect 1722 3488 1750 3491
rect 1906 3488 2006 3491
rect 2146 3488 2318 3491
rect 2322 3488 2342 3491
rect 2370 3488 2374 3491
rect 2402 3488 2462 3491
rect 2522 3488 2646 3491
rect 2650 3488 2726 3491
rect 2878 3491 2881 3498
rect 4742 3492 4745 3498
rect 2754 3488 2841 3491
rect 2878 3488 2950 3491
rect 3210 3488 3409 3491
rect 3434 3488 3486 3491
rect 3546 3488 3574 3491
rect 3666 3488 3718 3491
rect 4022 3488 4054 3491
rect 4130 3488 4206 3491
rect 4242 3488 4334 3491
rect 4338 3488 4345 3491
rect 4410 3488 4678 3491
rect 4698 3488 4710 3491
rect 4994 3488 5030 3491
rect 5034 3488 5038 3491
rect 5042 3488 5286 3491
rect 1094 3482 1097 3488
rect 2838 3482 2841 3488
rect 290 3478 510 3481
rect 762 3478 774 3481
rect 778 3478 814 3481
rect 826 3478 886 3481
rect 922 3478 966 3481
rect 1258 3478 1342 3481
rect 1346 3478 1438 3481
rect 1442 3478 1590 3481
rect 1658 3478 1774 3481
rect 1858 3478 2134 3481
rect 2202 3478 2217 3481
rect 2330 3478 2350 3481
rect 2354 3478 2414 3481
rect 2630 3478 2638 3481
rect 2642 3478 2686 3481
rect 2818 3478 2822 3481
rect 2978 3478 3078 3481
rect 3242 3478 3278 3481
rect 3290 3478 3398 3481
rect 3406 3481 3409 3488
rect 3406 3478 3558 3481
rect 3570 3478 3694 3481
rect 3762 3478 3774 3481
rect 3862 3481 3865 3488
rect 4022 3482 4025 3488
rect 3862 3478 3950 3481
rect 4178 3478 4270 3481
rect 4274 3478 4366 3481
rect 4370 3478 4454 3481
rect 4586 3478 4766 3481
rect 4926 3481 4929 3488
rect 4926 3478 5038 3481
rect 5042 3478 5078 3481
rect 5242 3478 5286 3481
rect 2214 3472 2217 3478
rect 3174 3472 3177 3478
rect 3998 3472 4001 3478
rect 58 3468 134 3471
rect 138 3468 166 3471
rect 210 3468 278 3471
rect 306 3468 446 3471
rect 454 3468 529 3471
rect 666 3468 694 3471
rect 898 3468 910 3471
rect 914 3468 982 3471
rect 986 3468 990 3471
rect 994 3468 1198 3471
rect 1202 3468 1206 3471
rect 1274 3468 1278 3471
rect 1410 3468 1470 3471
rect 1474 3468 1518 3471
rect 1522 3468 1534 3471
rect 1570 3468 1582 3471
rect 1594 3468 1678 3471
rect -26 3461 -22 3462
rect 6 3461 9 3468
rect -26 3458 30 3461
rect 274 3458 294 3461
rect 454 3461 457 3468
rect 526 3462 529 3468
rect 1790 3462 1793 3471
rect 1802 3468 1870 3471
rect 1874 3468 1918 3471
rect 1978 3468 2038 3471
rect 2186 3468 2206 3471
rect 2346 3468 2678 3471
rect 2690 3468 2798 3471
rect 2802 3468 2966 3471
rect 2970 3468 2982 3471
rect 2994 3468 3006 3471
rect 3186 3468 3550 3471
rect 3570 3468 3574 3471
rect 3730 3468 3774 3471
rect 4042 3468 4046 3471
rect 4050 3468 4070 3471
rect 4074 3468 4246 3471
rect 4250 3468 4278 3471
rect 4282 3468 4470 3471
rect 4722 3468 4814 3471
rect 4954 3468 4998 3471
rect 5018 3468 5086 3471
rect 5186 3468 5230 3471
rect 394 3458 457 3461
rect 506 3458 510 3461
rect 602 3458 638 3461
rect 642 3458 830 3461
rect 914 3458 918 3461
rect 954 3458 1009 3461
rect 1154 3458 1238 3461
rect 1282 3458 1286 3461
rect 1458 3458 1462 3461
rect 1514 3458 1590 3461
rect 1602 3458 1718 3461
rect 1722 3458 1742 3461
rect 1754 3458 1774 3461
rect 1810 3458 1814 3461
rect 1906 3459 1958 3461
rect 1906 3458 1961 3459
rect 1986 3458 2174 3461
rect 2206 3461 2209 3468
rect 2206 3458 2510 3461
rect 2570 3458 2638 3461
rect 2834 3458 3006 3461
rect 3138 3458 3142 3461
rect 3202 3458 3206 3461
rect 3282 3459 3326 3461
rect 4654 3462 4657 3468
rect 3282 3458 3329 3459
rect 3490 3458 3510 3461
rect 3514 3458 3542 3461
rect 3562 3458 3582 3461
rect 3626 3458 3702 3461
rect 3754 3458 3758 3461
rect 3802 3458 3822 3461
rect 3922 3458 4014 3461
rect 4066 3458 4142 3461
rect 4314 3458 4494 3461
rect 4522 3458 4598 3461
rect 4602 3458 4606 3461
rect 4618 3458 4654 3461
rect 4682 3458 4686 3461
rect 4690 3458 4694 3461
rect 4730 3458 4766 3461
rect 4846 3461 4849 3468
rect 4802 3458 4849 3461
rect 5142 3461 5145 3468
rect 5130 3458 5145 3461
rect 5186 3458 5238 3461
rect 1006 3452 1009 3458
rect 1494 3452 1497 3458
rect 1846 3452 1849 3458
rect 2702 3452 2705 3458
rect 266 3448 310 3451
rect 314 3448 494 3451
rect 554 3448 574 3451
rect 714 3448 862 3451
rect 1202 3448 1238 3451
rect 1242 3448 1270 3451
rect 1290 3448 1342 3451
rect 1534 3448 1550 3451
rect 1582 3448 1590 3451
rect 1594 3448 1646 3451
rect 1854 3448 2350 3451
rect 2354 3448 2550 3451
rect 2754 3448 2822 3451
rect 2826 3448 2950 3451
rect 3146 3448 3150 3451
rect 3234 3448 3302 3451
rect 3306 3448 3998 3451
rect 4002 3448 4006 3451
rect 4130 3448 4230 3451
rect 4490 3448 4601 3451
rect 4682 3448 4689 3451
rect 4770 3448 4870 3451
rect 4962 3448 4982 3451
rect 5026 3448 5038 3451
rect 5130 3448 5246 3451
rect 1518 3442 1521 3448
rect 1534 3442 1537 3448
rect 522 3438 710 3441
rect 714 3438 870 3441
rect 930 3438 942 3441
rect 1082 3438 1086 3441
rect 1202 3438 1486 3441
rect 1854 3441 1857 3448
rect 4598 3442 4601 3448
rect 4686 3442 4689 3448
rect 1770 3438 1857 3441
rect 2018 3438 2038 3441
rect 2190 3438 2198 3441
rect 2202 3438 2286 3441
rect 2378 3438 2502 3441
rect 2662 3438 2670 3441
rect 2674 3438 2750 3441
rect 2818 3438 2846 3441
rect 2850 3438 2886 3441
rect 3090 3438 3246 3441
rect 3250 3438 3542 3441
rect 3766 3438 3774 3441
rect 3778 3438 4086 3441
rect 4090 3438 4214 3441
rect 4634 3438 4654 3441
rect 5098 3438 5126 3441
rect 322 3428 390 3431
rect 394 3428 558 3431
rect 562 3428 574 3431
rect 926 3431 929 3438
rect 5134 3432 5137 3438
rect 578 3428 929 3431
rect 1170 3428 1542 3431
rect 1546 3428 2142 3431
rect 2146 3428 2318 3431
rect 2626 3428 3185 3431
rect 3354 3428 3454 3431
rect 3546 3428 4094 3431
rect 4146 3428 4190 3431
rect 4218 3428 4662 3431
rect 4666 3428 4790 3431
rect 3182 3422 3185 3428
rect 346 3418 398 3421
rect 442 3418 462 3421
rect 610 3418 782 3421
rect 866 3418 1254 3421
rect 1502 3418 1534 3421
rect 2106 3418 2246 3421
rect 2314 3418 2438 3421
rect 2586 3418 2726 3421
rect 2730 3418 2782 3421
rect 2954 3418 3126 3421
rect 3202 3418 3230 3421
rect 3234 3418 3302 3421
rect 3322 3418 3366 3421
rect 3390 3418 3510 3421
rect 3514 3418 3518 3421
rect 3594 3418 4078 3421
rect 4194 3418 4326 3421
rect 4330 3418 4510 3421
rect 4634 3418 4966 3421
rect 5234 3418 5262 3421
rect 1502 3412 1505 3418
rect 458 3408 478 3411
rect 626 3408 694 3411
rect 1594 3408 2166 3411
rect 2250 3408 2366 3411
rect 2514 3408 2710 3411
rect 2714 3408 2790 3411
rect 2930 3408 2974 3411
rect 2978 3408 3038 3411
rect 3066 3408 3174 3411
rect 3390 3411 3393 3418
rect 3298 3408 3393 3411
rect 3450 3408 3590 3411
rect 3594 3408 3598 3411
rect 3714 3408 3982 3411
rect 4474 3408 4830 3411
rect 4986 3408 5014 3411
rect 328 3403 330 3407
rect 334 3403 337 3407
rect 342 3403 344 3407
rect 1352 3403 1354 3407
rect 1358 3403 1361 3407
rect 1366 3403 1368 3407
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2398 3403 2400 3407
rect 3400 3403 3402 3407
rect 3406 3403 3409 3407
rect 3414 3403 3416 3407
rect 4424 3403 4426 3407
rect 4430 3403 4433 3407
rect 4438 3403 4440 3407
rect 602 3398 614 3401
rect 722 3398 806 3401
rect 810 3398 974 3401
rect 978 3398 1094 3401
rect 1426 3398 1750 3401
rect 1754 3398 1854 3401
rect 2034 3398 2158 3401
rect 2162 3398 2326 3401
rect 2426 3398 2446 3401
rect 2682 3398 2694 3401
rect 3218 3398 3246 3401
rect 3762 3398 3902 3401
rect 3906 3398 3982 3401
rect 4474 3398 4702 3401
rect 4706 3398 4910 3401
rect 4986 3398 4990 3401
rect 4994 3398 5030 3401
rect 166 3388 1118 3391
rect 1122 3388 1206 3391
rect 1210 3388 1310 3391
rect 1314 3388 1382 3391
rect 1450 3388 1630 3391
rect 2970 3388 3518 3391
rect 3522 3388 3526 3391
rect 3546 3388 4302 3391
rect 4306 3388 4758 3391
rect 4890 3388 5190 3391
rect 166 3382 169 3388
rect 506 3378 561 3381
rect 746 3378 1134 3381
rect 1266 3378 1294 3381
rect 1298 3378 1422 3381
rect 1498 3378 1526 3381
rect 1770 3378 1790 3381
rect 1810 3378 1822 3381
rect 2114 3378 2302 3381
rect 2306 3378 2622 3381
rect 2698 3378 2806 3381
rect 2882 3378 3414 3381
rect 3770 3378 3846 3381
rect 4066 3378 4110 3381
rect 4506 3378 4518 3381
rect 4546 3378 4550 3381
rect 4570 3378 4662 3381
rect 4738 3378 5006 3381
rect 5050 3378 5102 3381
rect 82 3368 118 3371
rect 350 3371 353 3378
rect 558 3372 561 3378
rect 266 3368 353 3371
rect 778 3368 982 3371
rect 986 3368 1038 3371
rect 1042 3368 1174 3371
rect 1254 3371 1257 3378
rect 1254 3368 1297 3371
rect 1322 3368 1494 3371
rect 1498 3368 1518 3371
rect 1522 3368 1550 3371
rect 1606 3371 1609 3378
rect 1554 3368 1609 3371
rect 1646 3368 1766 3371
rect 1770 3368 1814 3371
rect 2018 3368 2022 3371
rect 2138 3368 2142 3371
rect 2146 3368 2638 3371
rect 2674 3368 2694 3371
rect 2698 3368 2974 3371
rect 2978 3368 3054 3371
rect 3106 3368 3142 3371
rect 3162 3368 3214 3371
rect 3234 3368 3254 3371
rect 3490 3368 3598 3371
rect 4098 3368 4110 3371
rect 4406 3371 4409 3378
rect 4394 3368 4409 3371
rect 4482 3368 4486 3371
rect 4606 3368 4614 3371
rect 4618 3368 4654 3371
rect 4762 3368 4878 3371
rect 4882 3368 4926 3371
rect 4930 3368 4990 3371
rect 4994 3368 5102 3371
rect 5106 3368 5150 3371
rect -26 3361 -22 3362
rect -26 3358 222 3361
rect 374 3361 377 3368
rect 502 3362 505 3368
rect 558 3362 561 3368
rect 322 3358 430 3361
rect 570 3358 590 3361
rect 594 3358 742 3361
rect 750 3361 753 3368
rect 1294 3362 1297 3368
rect 1646 3362 1649 3368
rect 750 3358 878 3361
rect 882 3358 886 3361
rect 994 3358 1014 3361
rect 1146 3358 1150 3361
rect 1202 3358 1278 3361
rect 1298 3358 1326 3361
rect 1466 3358 1486 3361
rect 1490 3358 1502 3361
rect 1546 3358 1574 3361
rect 1586 3358 1598 3361
rect 1666 3358 1710 3361
rect 1770 3358 1774 3361
rect 1802 3358 1830 3361
rect 1922 3358 1934 3361
rect 1962 3358 1982 3361
rect 2030 3361 2033 3368
rect 1986 3358 2033 3361
rect 2058 3358 2134 3361
rect 2170 3358 2630 3361
rect 2734 3358 2742 3361
rect 2746 3358 2798 3361
rect 2938 3358 3046 3361
rect 3070 3361 3073 3368
rect 3070 3358 3166 3361
rect 3358 3361 3361 3368
rect 4486 3362 4489 3368
rect 3282 3358 3361 3361
rect 3426 3358 3430 3361
rect 3466 3358 3550 3361
rect 3570 3358 3574 3361
rect 3586 3358 3694 3361
rect 3738 3358 3782 3361
rect 3834 3358 3854 3361
rect 3874 3358 3958 3361
rect 4314 3358 4462 3361
rect 4498 3358 4518 3361
rect 4522 3358 4662 3361
rect 4722 3358 4726 3361
rect 4730 3358 4854 3361
rect 4898 3358 4942 3361
rect 5130 3358 5198 3361
rect 2670 3352 2673 3358
rect 106 3348 110 3351
rect 114 3348 1958 3351
rect 1962 3348 1966 3351
rect 1970 3348 1998 3351
rect 2002 3348 2166 3351
rect 2258 3348 2318 3351
rect 2442 3348 2470 3351
rect 2474 3348 2518 3351
rect 2618 3348 2662 3351
rect 2706 3348 2726 3351
rect 2730 3348 2758 3351
rect 2906 3348 3006 3351
rect 3010 3348 3038 3351
rect 3090 3348 3126 3351
rect 3282 3348 3286 3351
rect 3354 3348 3438 3351
rect 3442 3348 3486 3351
rect 3634 3348 3702 3351
rect 3858 3348 3902 3351
rect 3914 3348 3950 3351
rect 4098 3348 4126 3351
rect 4242 3348 4254 3351
rect 4258 3348 4366 3351
rect 4370 3348 4566 3351
rect 4642 3348 4742 3351
rect 4746 3348 4758 3351
rect 4786 3348 4798 3351
rect 4834 3348 4870 3351
rect 5118 3348 5206 3351
rect 18 3338 22 3341
rect 26 3338 118 3341
rect 122 3338 134 3341
rect 146 3338 174 3341
rect 522 3338 550 3341
rect 554 3338 630 3341
rect 634 3338 750 3341
rect 802 3338 806 3341
rect 834 3338 838 3341
rect 858 3338 878 3341
rect 890 3338 926 3341
rect 1026 3338 1118 3341
rect 1122 3338 1142 3341
rect 1162 3338 1318 3341
rect 1346 3340 1598 3341
rect 1342 3338 1598 3340
rect 1778 3338 1782 3341
rect 1954 3338 2006 3341
rect 2010 3338 2038 3341
rect 2074 3338 2078 3341
rect 2098 3338 2102 3341
rect 2122 3338 2126 3341
rect 2170 3338 2198 3341
rect 2314 3338 2326 3341
rect 2474 3338 2478 3341
rect 2482 3338 2486 3341
rect 2554 3338 2614 3341
rect 2642 3338 2654 3341
rect 2770 3338 2862 3341
rect 2906 3338 2910 3341
rect 3042 3338 3046 3341
rect 3058 3338 3094 3341
rect 3258 3338 3358 3341
rect 3450 3338 3534 3341
rect 3538 3338 3558 3341
rect 3570 3338 3590 3341
rect 3722 3338 3830 3341
rect 3890 3338 3966 3341
rect 3970 3338 4030 3341
rect 4074 3338 4078 3341
rect 4170 3338 4246 3341
rect 4278 3338 4302 3341
rect 4358 3338 4374 3341
rect 4498 3338 4502 3341
rect 4554 3338 4590 3341
rect 4730 3338 4798 3341
rect 4966 3341 4969 3348
rect 5118 3342 5121 3348
rect 4966 3338 5062 3341
rect 5130 3338 5134 3341
rect 5222 3341 5225 3348
rect 5222 3338 5246 3341
rect 5250 3338 5270 3341
rect 5290 3338 5294 3341
rect 482 3328 558 3331
rect 586 3328 590 3331
rect 634 3328 638 3331
rect 658 3328 670 3331
rect 810 3328 862 3331
rect 890 3328 902 3331
rect 990 3331 993 3338
rect 990 3328 1062 3331
rect 1082 3328 1126 3331
rect 1146 3328 1150 3331
rect 1410 3328 1470 3331
rect 1482 3328 1486 3331
rect 1530 3328 1622 3331
rect 1850 3328 1934 3331
rect 2186 3328 2313 3331
rect 2402 3328 2502 3331
rect 2562 3328 2641 3331
rect 742 3322 745 3328
rect 194 3318 302 3321
rect 402 3318 582 3321
rect 602 3318 646 3321
rect 746 3318 1318 3321
rect 1322 3318 1558 3321
rect 1562 3318 1566 3321
rect 1974 3321 1977 3328
rect 1898 3318 1977 3321
rect 2138 3318 2190 3321
rect 2210 3318 2294 3321
rect 2310 3321 2313 3328
rect 2638 3322 2641 3328
rect 2994 3328 3206 3331
rect 3218 3328 3334 3331
rect 3394 3328 3598 3331
rect 3606 3331 3609 3338
rect 3678 3332 3681 3338
rect 4278 3332 4281 3338
rect 4358 3332 4361 3338
rect 3606 3328 3614 3331
rect 3682 3328 3742 3331
rect 3746 3328 3750 3331
rect 3786 3328 3790 3331
rect 3802 3328 3830 3331
rect 3834 3328 3886 3331
rect 3950 3328 3958 3331
rect 3962 3328 4038 3331
rect 4050 3328 4214 3331
rect 4402 3328 4582 3331
rect 4690 3328 4710 3331
rect 4714 3328 4721 3331
rect 4746 3328 4798 3331
rect 4802 3328 4814 3331
rect 4834 3328 4838 3331
rect 4842 3328 4886 3331
rect 4954 3328 4966 3331
rect 5058 3328 5126 3331
rect 2710 3322 2713 3328
rect 2310 3318 2318 3321
rect 2602 3318 2614 3321
rect 2970 3318 3230 3321
rect 3426 3318 3526 3321
rect 3690 3318 3846 3321
rect 3910 3318 4102 3321
rect 4354 3318 4574 3321
rect 4578 3318 4630 3321
rect 4862 3318 4870 3321
rect 4874 3318 4934 3321
rect 4998 3318 5102 3321
rect 5154 3318 5174 3321
rect 1590 3312 1593 3318
rect 386 3308 518 3311
rect 538 3308 590 3311
rect 634 3308 734 3311
rect 746 3308 806 3311
rect 970 3308 1150 3311
rect 1274 3308 1510 3311
rect 1546 3308 1566 3311
rect 1618 3308 1822 3311
rect 2106 3308 2110 3311
rect 2178 3308 2262 3311
rect 2266 3308 2342 3311
rect 2466 3308 2598 3311
rect 2618 3308 2662 3311
rect 2794 3308 2838 3311
rect 3090 3308 3166 3311
rect 3362 3308 3438 3311
rect 3442 3308 3638 3311
rect 3642 3308 3718 3311
rect 3910 3311 3913 3318
rect 4998 3312 5001 3318
rect 3738 3308 3913 3311
rect 3946 3308 3982 3311
rect 4202 3308 4270 3311
rect 4298 3308 4486 3311
rect 4650 3308 4710 3311
rect 4986 3308 4998 3311
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 862 3303 864 3307
rect 1574 3302 1577 3308
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1886 3303 1888 3307
rect 2742 3302 2745 3308
rect 2888 3303 2890 3307
rect 2894 3303 2897 3307
rect 2902 3303 2904 3307
rect 3920 3303 3922 3307
rect 3926 3303 3929 3307
rect 3934 3303 3936 3307
rect 4936 3303 4938 3307
rect 4942 3303 4945 3307
rect 4950 3303 4952 3307
rect 66 3298 201 3301
rect 346 3298 446 3301
rect 450 3298 590 3301
rect 626 3298 702 3301
rect 2170 3298 2246 3301
rect 18 3288 102 3291
rect 198 3291 201 3298
rect 2254 3292 2257 3298
rect 2270 3292 2273 3301
rect 2442 3298 2510 3301
rect 2570 3298 2638 3301
rect 2642 3298 2734 3301
rect 2818 3298 2870 3301
rect 2930 3298 2942 3301
rect 2970 3298 3102 3301
rect 3170 3298 3270 3301
rect 3378 3298 3646 3301
rect 4098 3298 4478 3301
rect 4658 3298 4790 3301
rect 4818 3298 4838 3301
rect 198 3288 558 3291
rect 562 3288 678 3291
rect 682 3288 774 3291
rect 1394 3288 1494 3291
rect 1502 3288 1526 3291
rect 1562 3288 1582 3291
rect 1650 3288 1726 3291
rect 1762 3288 1894 3291
rect 1922 3288 1942 3291
rect 2034 3288 2137 3291
rect 2202 3288 2238 3291
rect 2286 3288 2294 3291
rect 2298 3288 2382 3291
rect 2570 3288 2670 3291
rect 2682 3288 2793 3291
rect 2834 3288 2838 3291
rect 2874 3288 2950 3291
rect 2962 3288 3014 3291
rect 3066 3288 3294 3291
rect 3338 3288 3366 3291
rect 3370 3288 3454 3291
rect 3506 3288 3670 3291
rect 3674 3288 3710 3291
rect 3722 3288 3886 3291
rect 3890 3288 3910 3291
rect 3994 3288 4014 3291
rect 4186 3288 4198 3291
rect 4338 3288 4358 3291
rect 4482 3288 4518 3291
rect 4530 3288 4886 3291
rect 4970 3288 5070 3291
rect 5074 3288 5158 3291
rect 5186 3288 5198 3291
rect 106 3278 278 3281
rect 450 3278 454 3281
rect 642 3278 694 3281
rect 698 3278 758 3281
rect 770 3278 846 3281
rect 882 3278 886 3281
rect 890 3278 910 3281
rect 1146 3278 1174 3281
rect 1482 3278 1486 3281
rect 1502 3281 1505 3288
rect 2134 3282 2137 3288
rect 1490 3278 1505 3281
rect 1514 3278 1622 3281
rect 1626 3278 1742 3281
rect 1834 3278 1910 3281
rect 2050 3278 2062 3281
rect 2218 3278 2390 3281
rect 2442 3278 2446 3281
rect 2494 3281 2497 3288
rect 2494 3278 2718 3281
rect 2730 3278 2782 3281
rect 2790 3281 2793 3288
rect 2790 3278 2990 3281
rect 3222 3278 3342 3281
rect 3354 3278 3382 3281
rect 3470 3281 3473 3288
rect 3470 3278 3558 3281
rect 3770 3278 3782 3281
rect 3946 3278 4022 3281
rect 4218 3278 4286 3281
rect 4314 3278 4542 3281
rect 4586 3278 4833 3281
rect 4850 3278 4902 3281
rect 4954 3278 5038 3281
rect 2726 3272 2729 3278
rect 194 3268 214 3271
rect 442 3268 534 3271
rect 762 3268 1102 3271
rect 1178 3268 1302 3271
rect 1338 3268 1342 3271
rect 1434 3268 1606 3271
rect 1722 3268 1758 3271
rect 1786 3268 1814 3271
rect 1826 3268 2182 3271
rect 2186 3268 2542 3271
rect 2682 3268 2686 3271
rect 2738 3268 3062 3271
rect 3126 3271 3129 3278
rect 3222 3272 3225 3278
rect 3126 3268 3134 3271
rect 3230 3268 3254 3271
rect 3290 3268 3294 3271
rect 3322 3268 3446 3271
rect 3582 3271 3585 3278
rect 3538 3268 3585 3271
rect 3618 3268 3694 3271
rect 3730 3268 3734 3271
rect 3738 3268 3870 3271
rect 4034 3268 4038 3271
rect 4078 3271 4081 3278
rect 4830 3272 4833 3278
rect 4078 3268 4086 3271
rect 4130 3268 4230 3271
rect 4362 3268 4454 3271
rect 4458 3268 4462 3271
rect 4490 3268 4494 3271
rect 4594 3268 4638 3271
rect 4794 3268 4798 3271
rect 4874 3268 4878 3271
rect 4910 3271 4913 3278
rect 4910 3268 4942 3271
rect 5122 3268 5150 3271
rect 5186 3268 5214 3271
rect 5250 3268 5294 3271
rect 70 3261 73 3268
rect 70 3258 86 3261
rect 198 3258 286 3261
rect 474 3258 478 3261
rect 670 3261 673 3268
rect 734 3262 737 3268
rect 670 3258 734 3261
rect 1002 3258 1086 3261
rect 1166 3261 1169 3268
rect 1166 3258 1209 3261
rect 1290 3258 1518 3261
rect 1522 3258 1526 3261
rect 1530 3258 2030 3261
rect 2034 3258 2038 3261
rect 2042 3258 2358 3261
rect 2362 3258 2470 3261
rect 2474 3258 2478 3261
rect 2482 3258 2494 3261
rect 2506 3258 2518 3261
rect 2706 3258 2742 3261
rect 2762 3258 2886 3261
rect 2890 3258 2934 3261
rect 2938 3258 2942 3261
rect 3230 3261 3233 3268
rect 2994 3258 3233 3261
rect 3242 3258 3270 3261
rect 3274 3258 3430 3261
rect 3502 3261 3505 3268
rect 3474 3258 3505 3261
rect 3530 3258 3558 3261
rect 3562 3258 3686 3261
rect 3690 3258 3942 3261
rect 3990 3261 3993 3268
rect 3990 3258 4022 3261
rect 4050 3258 4062 3261
rect 4082 3258 4158 3261
rect 4334 3261 4337 3268
rect 4210 3258 4337 3261
rect 4342 3261 4345 3268
rect 4510 3262 4513 3268
rect 4342 3258 4414 3261
rect 4482 3258 4486 3261
rect 4530 3258 4534 3261
rect 4578 3258 4582 3261
rect 4586 3258 4598 3261
rect 4618 3259 4734 3261
rect 4618 3258 4737 3259
rect 4818 3258 4838 3261
rect 4922 3258 4934 3261
rect 5210 3258 5254 3261
rect 5270 3258 5294 3261
rect 198 3252 201 3258
rect 918 3252 921 3258
rect 1158 3252 1161 3258
rect 1206 3252 1209 3258
rect 5270 3252 5273 3258
rect 638 3248 657 3251
rect 638 3242 641 3248
rect 654 3242 657 3248
rect 710 3248 838 3251
rect 842 3248 910 3251
rect 994 3248 1078 3251
rect 1106 3248 1126 3251
rect 1294 3248 1326 3251
rect 1450 3248 1454 3251
rect 1482 3248 1502 3251
rect 1530 3248 1534 3251
rect 1570 3248 1582 3251
rect 1594 3248 1606 3251
rect 1618 3248 1670 3251
rect 1706 3248 1846 3251
rect 1962 3248 2033 3251
rect 2042 3248 2246 3251
rect 2286 3248 2305 3251
rect 2482 3248 2486 3251
rect 2530 3248 2758 3251
rect 2810 3248 2830 3251
rect 2834 3248 2838 3251
rect 2858 3248 2990 3251
rect 3254 3248 3326 3251
rect 3338 3248 3814 3251
rect 3818 3248 3862 3251
rect 3922 3248 4025 3251
rect 4218 3248 4262 3251
rect 4266 3248 4313 3251
rect 4322 3248 4406 3251
rect 4410 3248 4534 3251
rect 4538 3248 4542 3251
rect 4590 3248 4598 3251
rect 4602 3248 4662 3251
rect 4842 3248 4846 3251
rect 4874 3248 5102 3251
rect 5154 3248 5166 3251
rect 710 3242 713 3248
rect 1294 3242 1297 3248
rect 674 3238 678 3241
rect 734 3238 774 3241
rect 874 3238 1182 3241
rect 1186 3238 1270 3241
rect 1470 3241 1473 3248
rect 1502 3242 1505 3248
rect 1470 3238 1486 3241
rect 1534 3238 1542 3241
rect 1546 3238 1550 3241
rect 1610 3238 1870 3241
rect 2030 3241 2033 3248
rect 2286 3242 2289 3248
rect 2302 3242 2305 3248
rect 3254 3242 3257 3248
rect 4022 3242 4025 3248
rect 2030 3238 2049 3241
rect 2098 3238 2102 3241
rect 2186 3238 2281 3241
rect 2418 3238 2686 3241
rect 2722 3238 2758 3241
rect 2778 3238 2806 3241
rect 2898 3238 2902 3241
rect 2970 3238 2974 3241
rect 3306 3238 3398 3241
rect 3466 3238 3558 3241
rect 3674 3238 3710 3241
rect 3746 3238 3774 3241
rect 3794 3238 3806 3241
rect 3810 3238 3814 3241
rect 3826 3238 3990 3241
rect 4058 3238 4270 3241
rect 4310 3241 4313 3248
rect 4310 3238 4558 3241
rect 4566 3241 4569 3248
rect 4862 3242 4865 3248
rect 4566 3238 4598 3241
rect 4874 3238 5166 3241
rect 734 3232 737 3238
rect 562 3228 726 3231
rect 842 3228 934 3231
rect 1330 3228 1478 3231
rect 1506 3228 1510 3231
rect 1514 3228 1702 3231
rect 2022 3231 2025 3238
rect 1822 3228 2025 3231
rect 2046 3232 2049 3238
rect 2110 3231 2113 3238
rect 2110 3228 2230 3231
rect 2278 3231 2281 3238
rect 2278 3228 2534 3231
rect 2538 3228 2646 3231
rect 2650 3228 2678 3231
rect 2722 3228 2750 3231
rect 2770 3228 3118 3231
rect 3138 3228 3190 3231
rect 3418 3228 3606 3231
rect 4138 3228 4182 3231
rect 4202 3228 4302 3231
rect 4306 3228 4398 3231
rect 4474 3228 4646 3231
rect 4786 3228 4966 3231
rect 5042 3228 5118 3231
rect 338 3218 414 3221
rect 418 3218 486 3221
rect 494 3221 497 3228
rect 494 3218 750 3221
rect 882 3218 918 3221
rect 970 3218 1022 3221
rect 1270 3221 1273 3228
rect 1822 3222 1825 3228
rect 1270 3218 1310 3221
rect 1514 3218 1710 3221
rect 1874 3218 1998 3221
rect 2010 3218 2070 3221
rect 2106 3218 2294 3221
rect 2298 3218 2374 3221
rect 2674 3218 2710 3221
rect 2858 3218 2910 3221
rect 3106 3218 3422 3221
rect 3858 3218 4470 3221
rect 4562 3218 5086 3221
rect 5090 3218 5118 3221
rect 5162 3218 5174 3221
rect 618 3208 718 3211
rect 874 3208 926 3211
rect 938 3208 1006 3211
rect 1010 3208 1206 3211
rect 1674 3208 1806 3211
rect 1866 3208 2254 3211
rect 2258 3208 2310 3211
rect 2450 3208 2526 3211
rect 2554 3208 2830 3211
rect 3046 3208 3142 3211
rect 3474 3208 4110 3211
rect 4258 3208 4366 3211
rect 4466 3208 4990 3211
rect 4994 3208 5038 3211
rect 5106 3208 5134 3211
rect 328 3203 330 3207
rect 334 3203 337 3207
rect 342 3203 344 3207
rect 1352 3203 1354 3207
rect 1358 3203 1361 3207
rect 1366 3203 1368 3207
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2398 3203 2400 3207
rect 3046 3202 3049 3208
rect 3400 3203 3402 3207
rect 3406 3203 3409 3207
rect 3414 3203 3416 3207
rect 4424 3203 4426 3207
rect 4430 3203 4433 3207
rect 4438 3203 4440 3207
rect 650 3198 686 3201
rect 690 3198 894 3201
rect 906 3198 942 3201
rect 954 3198 1134 3201
rect 1138 3198 1278 3201
rect 1618 3198 1654 3201
rect 1658 3198 1734 3201
rect 1794 3198 2190 3201
rect 2474 3198 2510 3201
rect 2610 3198 2766 3201
rect 2986 3198 3006 3201
rect 3010 3198 3046 3201
rect 3122 3198 3134 3201
rect 3138 3198 3393 3201
rect 3442 3198 3758 3201
rect 4034 3198 4150 3201
rect 4154 3198 4358 3201
rect 4498 3198 4518 3201
rect 4530 3198 4582 3201
rect 4602 3198 4870 3201
rect 5034 3198 5062 3201
rect 114 3188 1262 3191
rect 1278 3191 1281 3198
rect 1278 3188 1590 3191
rect 1706 3188 1782 3191
rect 2014 3188 2062 3191
rect 2786 3188 2894 3191
rect 2898 3188 3078 3191
rect 3082 3188 3382 3191
rect 3390 3191 3393 3198
rect 4990 3192 4993 3198
rect 3390 3188 4110 3191
rect 4114 3188 4118 3191
rect 4146 3188 4166 3191
rect 4186 3188 4326 3191
rect 4330 3188 4374 3191
rect 4386 3188 4689 3191
rect 4794 3188 4806 3191
rect 610 3178 638 3181
rect 642 3178 774 3181
rect 778 3178 870 3181
rect 890 3178 1014 3181
rect 1226 3178 1342 3181
rect 1394 3178 1478 3181
rect 1594 3178 1694 3181
rect 1934 3181 1937 3188
rect 2014 3182 2017 3188
rect 4686 3182 4689 3188
rect 1934 3178 1998 3181
rect 2042 3178 2046 3181
rect 2514 3178 2574 3181
rect 2698 3178 2726 3181
rect 2786 3178 2950 3181
rect 3042 3178 3158 3181
rect 3162 3178 3318 3181
rect 3434 3178 3510 3181
rect 3514 3178 3550 3181
rect 3690 3178 3790 3181
rect 3794 3178 3910 3181
rect 3914 3178 4361 3181
rect 178 3168 326 3171
rect 570 3168 630 3171
rect 634 3168 1094 3171
rect 1130 3168 1374 3171
rect 1382 3171 1385 3178
rect 4358 3172 4361 3178
rect 4530 3178 4550 3181
rect 4554 3178 4582 3181
rect 5166 3181 5169 3188
rect 4810 3178 5169 3181
rect 4518 3172 4521 3178
rect 1382 3168 1398 3171
rect 1458 3168 1478 3171
rect 1482 3168 1574 3171
rect 1638 3168 1734 3171
rect 1778 3168 2070 3171
rect 2082 3168 2142 3171
rect 2234 3168 2302 3171
rect 2490 3168 2638 3171
rect 2958 3168 3006 3171
rect 3126 3168 3222 3171
rect 3610 3168 3742 3171
rect 3746 3168 3998 3171
rect 4138 3168 4142 3171
rect 4346 3168 4350 3171
rect 4362 3168 4494 3171
rect 4534 3168 4542 3171
rect 4546 3168 4558 3171
rect 4570 3168 4854 3171
rect 4858 3168 4897 3171
rect 218 3158 510 3161
rect 586 3158 638 3161
rect 642 3158 710 3161
rect 762 3158 790 3161
rect 874 3158 934 3161
rect 1162 3158 1166 3161
rect 1250 3158 1390 3161
rect 1414 3161 1417 3168
rect 1410 3158 1417 3161
rect 1442 3158 1454 3161
rect 1490 3158 1494 3161
rect 1638 3161 1641 3168
rect 1554 3158 1641 3161
rect 1698 3158 1710 3161
rect 1906 3158 1990 3161
rect 1994 3158 2438 3161
rect 2498 3158 2518 3161
rect 2618 3158 2622 3161
rect 2654 3161 2657 3168
rect 2670 3161 2673 3168
rect 2654 3158 2673 3161
rect 2686 3161 2689 3168
rect 2838 3162 2841 3168
rect 2958 3162 2961 3168
rect 3126 3162 3129 3168
rect 2686 3158 2790 3161
rect 2818 3158 2822 3161
rect 2858 3158 2958 3161
rect 2994 3158 3054 3161
rect 3238 3161 3241 3168
rect 4894 3162 4897 3168
rect 3238 3158 3286 3161
rect 3450 3158 3454 3161
rect 3962 3158 4046 3161
rect 4106 3158 4150 3161
rect 4154 3158 4190 3161
rect 4290 3158 4334 3161
rect 4346 3158 4433 3161
rect 1190 3152 1193 3158
rect 298 3148 302 3151
rect 314 3148 345 3151
rect 18 3138 22 3141
rect 70 3141 73 3148
rect 86 3141 89 3148
rect 182 3141 185 3148
rect 70 3138 185 3141
rect 342 3142 345 3148
rect 610 3148 622 3151
rect 658 3148 670 3151
rect 690 3148 694 3151
rect 698 3148 710 3151
rect 730 3148 790 3151
rect 802 3148 822 3151
rect 826 3148 830 3151
rect 834 3148 894 3151
rect 914 3148 953 3151
rect 422 3141 425 3148
rect 950 3142 953 3148
rect 1090 3148 1174 3151
rect 1238 3148 1289 3151
rect 1426 3148 1542 3151
rect 1626 3148 1630 3151
rect 1666 3148 1670 3151
rect 1698 3148 1742 3151
rect 1806 3151 1809 3158
rect 2486 3152 2489 3158
rect 2550 3152 2553 3158
rect 1806 3148 1838 3151
rect 1846 3148 1942 3151
rect 1970 3148 1985 3151
rect 2098 3148 2110 3151
rect 2154 3148 2222 3151
rect 2262 3148 2270 3151
rect 2434 3148 2481 3151
rect 2570 3148 2654 3151
rect 2794 3148 2934 3151
rect 2970 3148 2998 3151
rect 3142 3151 3145 3158
rect 3198 3152 3201 3158
rect 3894 3152 3897 3158
rect 4430 3152 4433 3158
rect 4562 3158 4606 3161
rect 4698 3158 4726 3161
rect 4818 3158 4822 3161
rect 5058 3158 5078 3161
rect 5098 3158 5110 3161
rect 5142 3161 5145 3168
rect 5142 3158 5238 3161
rect 3034 3148 3145 3151
rect 3154 3148 3182 3151
rect 3254 3148 3358 3151
rect 3482 3148 3662 3151
rect 3666 3148 3678 3151
rect 3730 3148 3734 3151
rect 3794 3148 3806 3151
rect 3850 3148 3862 3151
rect 4066 3148 4086 3151
rect 4130 3148 4134 3151
rect 4162 3148 4182 3151
rect 4418 3148 4422 3151
rect 4438 3151 4441 3158
rect 4534 3152 4537 3158
rect 4886 3152 4889 3158
rect 4438 3148 4446 3151
rect 4522 3148 4526 3151
rect 4578 3148 4582 3151
rect 4594 3148 4638 3151
rect 4730 3148 4758 3151
rect 4866 3148 4870 3151
rect 4910 3151 4913 3158
rect 4910 3148 4934 3151
rect 5002 3148 5118 3151
rect 5126 3151 5129 3158
rect 5122 3148 5129 3151
rect 5194 3148 5222 3151
rect 422 3138 446 3141
rect 506 3138 614 3141
rect 682 3138 718 3141
rect 722 3138 726 3141
rect 738 3138 854 3141
rect 1030 3141 1033 3148
rect 1054 3142 1057 3148
rect 1238 3142 1241 3148
rect 1286 3142 1289 3148
rect 1566 3142 1569 3148
rect 1030 3138 1054 3141
rect 1162 3138 1174 3141
rect 1178 3138 1182 3141
rect 1210 3138 1214 3141
rect 1354 3138 1438 3141
rect 1482 3138 1558 3141
rect 1606 3141 1609 3148
rect 1606 3138 1622 3141
rect 1642 3138 1646 3141
rect 1674 3138 1686 3141
rect 1774 3141 1777 3148
rect 1846 3142 1849 3148
rect 1982 3142 1985 3148
rect 2262 3142 2265 3148
rect 2278 3142 2281 3148
rect 2310 3142 2313 3148
rect 2478 3142 2481 3148
rect 3254 3142 3257 3148
rect 1774 3138 1806 3141
rect 2090 3138 2238 3141
rect 2330 3138 2358 3141
rect 2514 3138 2630 3141
rect 2682 3138 2822 3141
rect 2826 3138 2846 3141
rect 2850 3138 2942 3141
rect 2954 3138 2998 3141
rect 3178 3138 3222 3141
rect 3434 3138 3470 3141
rect 3546 3138 3590 3141
rect 3838 3141 3841 3148
rect 3838 3138 3854 3141
rect 4030 3141 4033 3148
rect 3858 3138 4118 3141
rect 4286 3141 4289 3148
rect 4726 3142 4729 3148
rect 4122 3138 4350 3141
rect 4354 3138 4446 3141
rect 4450 3138 4590 3141
rect 4746 3138 4750 3141
rect 4754 3138 4758 3141
rect 4794 3138 4798 3141
rect 4866 3138 4894 3141
rect 4974 3138 5030 3141
rect 5050 3138 5150 3141
rect 5154 3138 5174 3141
rect 186 3128 198 3131
rect 402 3128 438 3131
rect 594 3128 598 3131
rect 610 3128 798 3131
rect 818 3128 822 3131
rect 850 3128 894 3131
rect 898 3128 966 3131
rect 1018 3128 1078 3131
rect 1102 3131 1105 3138
rect 1462 3132 1465 3138
rect 1478 3132 1481 3138
rect 1102 3128 1126 3131
rect 1146 3128 1254 3131
rect 1402 3128 1406 3131
rect 1494 3128 1526 3131
rect 1602 3128 1630 3131
rect 1654 3131 1657 3138
rect 1654 3128 1782 3131
rect 1802 3128 2086 3131
rect 2122 3128 2350 3131
rect 2482 3128 2486 3131
rect 2654 3131 2657 3138
rect 3110 3132 3113 3138
rect 4974 3132 4977 3138
rect 5198 3132 5201 3138
rect 2538 3128 2569 3131
rect 2654 3128 2726 3131
rect 2842 3128 2854 3131
rect 2906 3128 3054 3131
rect 3170 3128 3446 3131
rect 3530 3128 3654 3131
rect 4018 3128 4070 3131
rect 4186 3128 4262 3131
rect 4370 3128 4382 3131
rect 4410 3128 4414 3131
rect 4474 3128 4518 3131
rect 4570 3128 4646 3131
rect 4874 3128 4974 3131
rect 5018 3128 5038 3131
rect 5082 3128 5110 3131
rect 5206 3131 5209 3138
rect 5206 3128 5230 3131
rect 1494 3122 1497 3128
rect 130 3118 169 3121
rect 218 3118 254 3121
rect 258 3118 566 3121
rect 586 3118 646 3121
rect 650 3118 726 3121
rect 730 3118 734 3121
rect 746 3118 782 3121
rect 802 3118 1246 3121
rect 1450 3118 1462 3121
rect 1542 3121 1545 3128
rect 1542 3118 1926 3121
rect 2018 3118 2022 3121
rect 2298 3118 2326 3121
rect 2346 3118 2550 3121
rect 2554 3118 2558 3121
rect 2566 3121 2569 3128
rect 2566 3118 2662 3121
rect 2666 3118 2686 3121
rect 2786 3118 3150 3121
rect 3170 3118 3430 3121
rect 3518 3121 3521 3128
rect 3518 3118 3534 3121
rect 3802 3118 3910 3121
rect 4338 3118 4366 3121
rect 4398 3121 4401 3128
rect 4398 3118 4422 3121
rect 5054 3121 5057 3128
rect 4650 3118 5057 3121
rect 5178 3118 5294 3121
rect 166 3112 169 3118
rect 4062 3112 4065 3118
rect 4518 3112 4521 3118
rect 234 3108 390 3111
rect 394 3108 478 3111
rect 578 3108 614 3111
rect 682 3108 766 3111
rect 1066 3108 1238 3111
rect 1442 3108 1502 3111
rect 1586 3108 1617 3111
rect 1626 3108 1798 3111
rect 1954 3108 2038 3111
rect 2074 3108 2129 3111
rect 2138 3108 2641 3111
rect 2650 3108 2790 3111
rect 3074 3108 3470 3111
rect 3586 3108 3630 3111
rect 4090 3108 4478 3111
rect 4738 3108 4758 3111
rect 4842 3108 4894 3111
rect 4898 3108 4910 3111
rect 5098 3108 5118 3111
rect 838 3102 841 3108
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 862 3103 864 3107
rect 226 3098 366 3101
rect 378 3098 678 3101
rect 1026 3098 1070 3101
rect 1074 3098 1286 3101
rect 1314 3098 1449 3101
rect 1466 3098 1470 3101
rect 1578 3098 1606 3101
rect 1614 3101 1617 3108
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1886 3103 1888 3107
rect 2126 3102 2129 3108
rect 1614 3098 1822 3101
rect 1898 3098 1934 3101
rect 1938 3098 2022 3101
rect 2290 3098 2486 3101
rect 2570 3098 2598 3101
rect 2638 3101 2641 3108
rect 2888 3103 2890 3107
rect 2894 3103 2897 3107
rect 2902 3103 2904 3107
rect 3920 3103 3922 3107
rect 3926 3103 3929 3107
rect 3934 3103 3936 3107
rect 4936 3103 4938 3107
rect 4942 3103 4945 3107
rect 4950 3103 4952 3107
rect 2638 3098 2878 3101
rect 2922 3098 2942 3101
rect 2982 3098 3006 3101
rect 3178 3098 3206 3101
rect 3394 3098 3662 3101
rect 3946 3098 3982 3101
rect 3986 3098 4238 3101
rect 4242 3098 4270 3101
rect 4274 3098 4310 3101
rect 4466 3098 4470 3101
rect 4474 3098 4502 3101
rect 4714 3098 4758 3101
rect 4762 3098 4838 3101
rect 4858 3098 4918 3101
rect 4970 3098 5110 3101
rect 170 3088 374 3091
rect 498 3088 598 3091
rect 634 3088 750 3091
rect 778 3088 1206 3091
rect 1282 3088 1382 3091
rect 1446 3091 1449 3098
rect 2494 3092 2497 3098
rect 1446 3088 1478 3091
rect 1534 3088 1574 3091
rect 1586 3088 2054 3091
rect 2066 3088 2158 3091
rect 2186 3088 2478 3091
rect 2634 3088 2702 3091
rect 2706 3088 2878 3091
rect 2982 3091 2985 3098
rect 2882 3088 2985 3091
rect 3058 3088 3118 3091
rect 3218 3088 3302 3091
rect 3434 3088 3454 3091
rect 3482 3088 3633 3091
rect 82 3078 270 3081
rect 274 3078 414 3081
rect 418 3078 606 3081
rect 610 3078 662 3081
rect 682 3078 846 3081
rect 850 3078 942 3081
rect 970 3078 1038 3081
rect 1178 3078 1334 3081
rect 1378 3078 1414 3081
rect 1438 3081 1441 3088
rect 1534 3081 1537 3088
rect 3630 3082 3633 3088
rect 3770 3088 3934 3091
rect 4026 3088 4030 3091
rect 4050 3088 4134 3091
rect 4266 3088 4438 3091
rect 4498 3088 4630 3091
rect 4674 3088 4742 3091
rect 4746 3088 4870 3091
rect 4906 3088 4910 3091
rect 5194 3088 5230 3091
rect 5234 3088 5246 3091
rect 1438 3078 1537 3081
rect 1546 3078 1550 3081
rect 1562 3078 1566 3081
rect 1594 3078 1622 3081
rect 1654 3078 1662 3081
rect 1674 3078 1718 3081
rect 1722 3078 1726 3081
rect 1850 3078 1894 3081
rect 1938 3078 1982 3081
rect 2098 3078 2126 3081
rect 2298 3078 2342 3081
rect 2562 3078 2678 3081
rect 2682 3078 2758 3081
rect 2842 3078 2846 3081
rect 2930 3078 3126 3081
rect 3210 3078 3238 3081
rect 3274 3078 3326 3081
rect 3546 3078 3598 3081
rect 3682 3078 3705 3081
rect 3758 3081 3761 3088
rect 3722 3078 3761 3081
rect 3810 3078 3886 3081
rect 3894 3078 4262 3081
rect 4266 3078 4310 3081
rect 4314 3078 4358 3081
rect 4378 3078 4526 3081
rect 4578 3078 5046 3081
rect 5202 3078 5214 3081
rect 1654 3072 1657 3078
rect 3126 3072 3129 3078
rect 3662 3072 3665 3078
rect 10 3068 214 3071
rect 362 3068 406 3071
rect 514 3068 614 3071
rect 618 3068 662 3071
rect 666 3068 670 3071
rect 674 3068 990 3071
rect 1066 3068 1158 3071
rect 1346 3068 1638 3071
rect 1698 3068 1838 3071
rect 1874 3068 1886 3071
rect 2002 3068 2046 3071
rect 2142 3068 2150 3071
rect 2154 3068 2310 3071
rect 2362 3068 2422 3071
rect 2426 3068 2470 3071
rect 2602 3068 2606 3071
rect 2634 3068 3038 3071
rect 3090 3068 3094 3071
rect 3322 3068 3350 3071
rect 3386 3068 3414 3071
rect 3434 3068 3470 3071
rect 3490 3068 3574 3071
rect 3594 3068 3606 3071
rect 3674 3068 3678 3071
rect 3702 3071 3705 3078
rect 3702 3068 3849 3071
rect 3866 3068 3870 3071
rect 3874 3068 3886 3071
rect 3894 3071 3897 3078
rect 3890 3068 3897 3071
rect 3906 3068 3942 3071
rect 3986 3068 4038 3071
rect 4170 3068 4174 3071
rect 4178 3068 4310 3071
rect 4314 3068 4934 3071
rect 4938 3068 4998 3071
rect 5078 3071 5081 3078
rect 5078 3068 5126 3071
rect 90 3058 102 3061
rect 178 3058 198 3061
rect 450 3058 558 3061
rect 562 3058 598 3061
rect 626 3058 662 3061
rect 778 3058 790 3061
rect 810 3059 870 3061
rect 810 3058 873 3059
rect 1010 3058 1038 3061
rect 1138 3058 1166 3061
rect 1182 3061 1185 3068
rect 1326 3062 1329 3068
rect 1182 3058 1198 3061
rect 1226 3058 1230 3061
rect 1334 3061 1337 3068
rect 1334 3058 1398 3061
rect 1418 3058 1438 3061
rect 1450 3058 1454 3061
rect 1474 3058 1486 3061
rect 1490 3058 1598 3061
rect 1650 3058 1838 3061
rect 1866 3058 1870 3061
rect 1918 3061 1921 3068
rect 1882 3058 1921 3061
rect 2058 3058 2070 3061
rect 2082 3058 2110 3061
rect 2126 3061 2129 3068
rect 2126 3058 2262 3061
rect 2310 3061 2313 3068
rect 2558 3062 2561 3068
rect 2310 3058 2454 3061
rect 2514 3058 2518 3061
rect 2594 3058 2598 3061
rect 2618 3058 2638 3061
rect 2658 3058 2782 3061
rect 2786 3058 2830 3061
rect 2842 3058 2862 3061
rect 2866 3058 2886 3061
rect 2930 3058 3022 3061
rect 3062 3061 3065 3068
rect 3694 3062 3697 3068
rect 3846 3062 3849 3068
rect 3026 3058 3065 3061
rect 3082 3058 3246 3061
rect 3250 3058 3334 3061
rect 3338 3058 3622 3061
rect 3626 3058 3630 3061
rect 3642 3058 3646 3061
rect 3746 3058 3750 3061
rect 3914 3058 3958 3061
rect 4026 3058 4030 3061
rect 4034 3058 4038 3061
rect 4154 3058 4198 3061
rect 4234 3058 4257 3061
rect 158 3052 161 3058
rect 198 3052 201 3058
rect 558 3052 561 3058
rect 650 3048 694 3051
rect 1106 3048 1198 3051
rect 1202 3048 1270 3051
rect 1278 3048 1310 3051
rect 1370 3048 1374 3051
rect 1386 3048 1446 3051
rect 1450 3048 1454 3051
rect 1490 3048 1598 3051
rect 1622 3051 1625 3058
rect 4254 3052 4257 3058
rect 4266 3058 4302 3061
rect 4378 3058 4478 3061
rect 4602 3058 4606 3061
rect 4698 3058 4702 3061
rect 4722 3058 4758 3061
rect 4778 3058 4942 3061
rect 4946 3058 4958 3061
rect 5114 3058 5142 3061
rect 4262 3052 4265 3058
rect 1622 3048 1702 3051
rect 1706 3048 1726 3051
rect 1858 3048 1862 3051
rect 1890 3048 1894 3051
rect 1906 3048 2062 3051
rect 2282 3048 2366 3051
rect 2378 3048 2438 3051
rect 2450 3048 2502 3051
rect 2530 3048 2534 3051
rect 2546 3048 2582 3051
rect 2622 3048 2630 3051
rect 2634 3048 2718 3051
rect 2786 3048 2790 3051
rect 2834 3048 2934 3051
rect 2946 3048 3086 3051
rect 3098 3048 3118 3051
rect 3146 3048 3150 3051
rect 3338 3048 3374 3051
rect 3378 3048 3414 3051
rect 3458 3048 3622 3051
rect 3714 3048 3721 3051
rect 818 3038 934 3041
rect 1278 3041 1281 3048
rect 3718 3042 3721 3048
rect 3886 3048 3894 3051
rect 4106 3048 4174 3051
rect 4298 3048 4414 3051
rect 4454 3048 4462 3051
rect 4466 3048 4574 3051
rect 4642 3048 4646 3051
rect 4714 3048 4718 3051
rect 4762 3048 4766 3051
rect 4914 3048 4974 3051
rect 4986 3048 4998 3051
rect 3886 3042 3889 3048
rect 938 3038 1281 3041
rect 1306 3038 1422 3041
rect 1442 3038 1582 3041
rect 1610 3038 1622 3041
rect 1642 3038 1894 3041
rect 2170 3038 2270 3041
rect 2306 3038 2310 3041
rect 2490 3038 2774 3041
rect 2866 3038 2982 3041
rect 2994 3038 3078 3041
rect 3082 3038 3302 3041
rect 3338 3038 3366 3041
rect 3386 3038 3454 3041
rect 4002 3038 4086 3041
rect 4310 3038 4350 3041
rect 4658 3038 4798 3041
rect 4886 3041 4889 3048
rect 4802 3038 4889 3041
rect 4902 3041 4905 3048
rect 4902 3038 4918 3041
rect 562 3028 574 3031
rect 578 3028 1078 3031
rect 1530 3028 1582 3031
rect 1682 3028 1782 3031
rect 1826 3028 1854 3031
rect 1890 3028 2110 3031
rect 2134 3028 2137 3038
rect 4310 3032 4313 3038
rect 2922 3028 3030 3031
rect 3034 3028 3038 3031
rect 3154 3028 3158 3031
rect 3178 3028 3358 3031
rect 3366 3028 3590 3031
rect 3682 3028 3782 3031
rect 3818 3028 4006 3031
rect 4010 3028 4054 3031
rect 4138 3028 4198 3031
rect 4330 3028 4398 3031
rect 4426 3028 4494 3031
rect 4510 3031 4513 3038
rect 4510 3028 4774 3031
rect 4914 3028 4926 3031
rect 4962 3028 5190 3031
rect 306 3018 326 3021
rect 330 3018 614 3021
rect 754 3018 1078 3021
rect 1298 3018 1598 3021
rect 1606 3021 1609 3028
rect 3046 3022 3049 3028
rect 1606 3018 1686 3021
rect 1954 3018 1958 3021
rect 1994 3018 2094 3021
rect 2098 3018 2126 3021
rect 2474 3018 2718 3021
rect 2722 3018 2830 3021
rect 3090 3018 3102 3021
rect 3366 3021 3369 3028
rect 3250 3018 3369 3021
rect 3394 3018 3494 3021
rect 3498 3018 3878 3021
rect 3882 3018 3958 3021
rect 4066 3018 4142 3021
rect 4386 3018 4694 3021
rect 5094 3018 5110 3021
rect 5178 3018 5190 3021
rect 5234 3018 5238 3021
rect 5258 3018 5286 3021
rect 5094 3012 5097 3018
rect 770 3008 926 3011
rect 1426 3008 1478 3011
rect 1482 3008 1742 3011
rect 1826 3008 1910 3011
rect 2202 3008 2350 3011
rect 2570 3008 2654 3011
rect 2842 3008 3070 3011
rect 3202 3008 3358 3011
rect 3474 3008 4190 3011
rect 4194 3008 4222 3011
rect 4394 3008 4406 3011
rect 4482 3008 4518 3011
rect 4586 3008 5014 3011
rect 5026 3008 5033 3011
rect 5106 3008 5230 3011
rect 5234 3008 5278 3011
rect 328 3003 330 3007
rect 334 3003 337 3007
rect 342 3003 344 3007
rect 1352 3003 1354 3007
rect 1358 3003 1361 3007
rect 1366 3003 1368 3007
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2398 3003 2400 3007
rect 3400 3003 3402 3007
rect 3406 3003 3409 3007
rect 3414 3003 3416 3007
rect 4424 3003 4426 3007
rect 4430 3003 4433 3007
rect 4438 3003 4440 3007
rect 666 2998 1142 3001
rect 1290 2998 1294 3001
rect 1394 2998 1614 3001
rect 1618 2998 1654 3001
rect 2074 2998 2182 3001
rect 2274 2998 2366 3001
rect 2666 2998 3014 3001
rect 3034 2998 3174 3001
rect 3274 2998 3286 3001
rect 3290 2998 3302 3001
rect 3562 2998 3598 3001
rect 3738 2998 4022 3001
rect 4170 2998 4198 3001
rect 4562 2998 4782 3001
rect 4890 2998 4966 3001
rect 4970 2998 5022 3001
rect 5030 3001 5033 3008
rect 5030 2998 5102 3001
rect 282 2988 286 2991
rect 410 2988 742 2991
rect 754 2988 774 2991
rect 1210 2988 1270 2991
rect 1274 2988 1462 2991
rect 1634 2988 1702 2991
rect 1798 2988 2078 2991
rect 2082 2988 2238 2991
rect 2242 2988 2246 2991
rect 2250 2988 2334 2991
rect 2338 2988 2454 2991
rect 2470 2991 2473 2998
rect 2466 2988 2473 2991
rect 2570 2988 3062 2991
rect 3258 2988 3390 2991
rect 3442 2988 3478 2991
rect 3710 2988 3718 2991
rect 3722 2988 3742 2991
rect 3890 2988 3894 2991
rect 3898 2988 3926 2991
rect 3930 2988 4318 2991
rect 4322 2988 4454 2991
rect 4458 2988 4582 2991
rect 4690 2988 4913 2991
rect 1798 2982 1801 2988
rect 4910 2982 4913 2988
rect 5130 2988 5134 2991
rect 298 2978 310 2981
rect 458 2978 638 2981
rect 738 2978 1062 2981
rect 1074 2978 1086 2981
rect 1090 2978 1622 2981
rect 1914 2978 1966 2981
rect 2250 2978 2550 2981
rect 2554 2978 3174 2981
rect 3186 2978 3198 2981
rect 3210 2978 3350 2981
rect 3354 2978 3521 2981
rect 3586 2978 3686 2981
rect 3706 2978 3806 2981
rect 4006 2978 4414 2981
rect 4418 2978 4470 2981
rect 4698 2978 4702 2981
rect 4706 2978 4902 2981
rect 4990 2981 4993 2988
rect 4914 2978 4993 2981
rect 3518 2972 3521 2978
rect 4006 2972 4009 2978
rect 5134 2972 5137 2978
rect 170 2968 518 2971
rect 610 2968 654 2971
rect 1322 2968 1342 2971
rect 1522 2968 1534 2971
rect 1650 2968 1678 2971
rect 2482 2968 2502 2971
rect 2678 2968 2686 2971
rect 2690 2968 2766 2971
rect 2818 2968 3142 2971
rect 3202 2968 3230 2971
rect 3314 2968 3414 2971
rect 3570 2968 3758 2971
rect 3802 2968 4006 2971
rect 4158 2968 4214 2971
rect 4378 2968 4390 2971
rect 4394 2968 4446 2971
rect 4474 2968 4486 2971
rect 4666 2968 4734 2971
rect 4738 2968 4966 2971
rect 146 2958 310 2961
rect 758 2961 761 2968
rect 714 2958 761 2961
rect 1274 2958 2006 2961
rect 2054 2961 2057 2968
rect 4158 2962 4161 2968
rect 4334 2962 4337 2968
rect 2054 2958 2318 2961
rect 2346 2958 2478 2961
rect 2482 2958 2518 2961
rect 2522 2958 2574 2961
rect 2650 2958 2670 2961
rect 2674 2958 2710 2961
rect 2994 2958 3030 2961
rect 3162 2958 3198 2961
rect 3514 2958 3702 2961
rect 3770 2958 3798 2961
rect 3930 2958 3974 2961
rect 3994 2958 4022 2961
rect 4058 2958 4078 2961
rect 4402 2958 4406 2961
rect 4418 2958 4422 2961
rect 4482 2958 4486 2961
rect 4514 2958 4681 2961
rect 4706 2958 4822 2961
rect 4874 2958 5094 2961
rect 5098 2958 5182 2961
rect 606 2952 609 2958
rect 610 2948 662 2951
rect 810 2948 814 2951
rect 866 2948 902 2951
rect 942 2951 945 2958
rect 914 2948 1030 2951
rect 1138 2948 1142 2951
rect 1158 2951 1161 2958
rect 1158 2948 1166 2951
rect 1258 2948 1262 2951
rect 1466 2948 1582 2951
rect 1586 2948 1654 2951
rect 1662 2948 1718 2951
rect 1738 2948 1785 2951
rect 1810 2948 1822 2951
rect 1954 2948 1966 2951
rect 2002 2948 2014 2951
rect 2106 2948 2206 2951
rect 2258 2948 2262 2951
rect 2362 2948 2414 2951
rect 2434 2948 2446 2951
rect 2506 2948 2510 2951
rect 2626 2948 2702 2951
rect 2862 2951 2865 2958
rect 2862 2948 2942 2951
rect 2978 2948 2990 2951
rect 3154 2948 3222 2951
rect 3234 2948 3254 2951
rect 3378 2948 3382 2951
rect 3538 2948 3558 2951
rect 3650 2948 3718 2951
rect 3746 2948 3942 2951
rect 3986 2948 4046 2951
rect 4210 2948 4310 2951
rect 4314 2948 4350 2951
rect 4358 2951 4361 2958
rect 4678 2952 4681 2958
rect 4358 2948 4366 2951
rect 4394 2948 4582 2951
rect 4786 2948 4862 2951
rect 4866 2948 4937 2951
rect 4946 2948 5030 2951
rect 5218 2948 5270 2951
rect 5334 2951 5338 2952
rect 5298 2948 5338 2951
rect 126 2941 129 2948
rect 222 2941 225 2948
rect 66 2938 225 2941
rect 318 2941 321 2948
rect 678 2942 681 2948
rect 718 2942 721 2948
rect 1662 2942 1665 2948
rect 1782 2942 1785 2948
rect 2998 2942 3001 2948
rect 318 2938 350 2941
rect 626 2938 638 2941
rect 1098 2938 1102 2941
rect 1146 2938 1190 2941
rect 1258 2938 1262 2941
rect 1338 2938 1358 2941
rect 1410 2938 1422 2941
rect 1578 2938 1638 2941
rect 1818 2938 1822 2941
rect 1842 2938 1974 2941
rect 1978 2938 2070 2941
rect 2178 2938 2214 2941
rect 2258 2938 2342 2941
rect 2490 2938 2534 2941
rect 2562 2938 2566 2941
rect 2570 2938 2582 2941
rect 2618 2938 2654 2941
rect 2658 2938 2702 2941
rect 2754 2938 2758 2941
rect 3034 2938 3198 2941
rect 3202 2938 3246 2941
rect 3354 2938 3366 2941
rect 3390 2938 3393 2948
rect 3982 2942 3985 2948
rect 3482 2938 3534 2941
rect 3634 2938 3958 2941
rect 3962 2938 3982 2941
rect 4026 2938 4078 2941
rect 4082 2938 4174 2941
rect 4194 2938 4198 2941
rect 4306 2938 4494 2941
rect 4498 2938 4502 2941
rect 4514 2938 4518 2941
rect 4530 2938 4566 2941
rect 4734 2941 4737 2948
rect 4934 2942 4937 2948
rect 5150 2942 5153 2948
rect 4666 2938 4737 2941
rect 4834 2938 4846 2941
rect 4874 2938 4878 2941
rect 4938 2938 5038 2941
rect 5154 2938 5166 2941
rect 5258 2938 5286 2941
rect 74 2928 166 2931
rect 250 2928 329 2931
rect 326 2922 329 2928
rect 546 2928 630 2931
rect 690 2928 694 2931
rect 698 2928 878 2931
rect 1054 2931 1057 2938
rect 2486 2932 2489 2938
rect 3430 2932 3433 2938
rect 4526 2932 4529 2938
rect 882 2928 1057 2931
rect 1122 2928 1254 2931
rect 1258 2928 1310 2931
rect 1354 2928 1526 2931
rect 1538 2928 1742 2931
rect 1746 2928 1785 2931
rect 1818 2928 1830 2931
rect 2074 2928 2078 2931
rect 2090 2928 2230 2931
rect 2322 2928 2481 2931
rect 2554 2928 2598 2931
rect 2610 2928 2990 2931
rect 3034 2928 3070 2931
rect 3074 2928 3206 2931
rect 3222 2928 3238 2931
rect 3290 2928 3302 2931
rect 3386 2928 3422 2931
rect 3450 2928 3574 2931
rect 3642 2928 3934 2931
rect 3974 2928 3982 2931
rect 3986 2928 4030 2931
rect 4114 2928 4142 2931
rect 4178 2928 4278 2931
rect 4374 2928 4406 2931
rect 4418 2928 4446 2931
rect 4490 2928 4518 2931
rect 4554 2928 4622 2931
rect 4762 2928 4862 2931
rect 4986 2928 5134 2931
rect 5138 2928 5294 2931
rect 18 2918 102 2921
rect 154 2918 214 2921
rect 398 2921 401 2928
rect 398 2918 502 2921
rect 642 2918 686 2921
rect 698 2918 750 2921
rect 770 2918 870 2921
rect 978 2918 1318 2921
rect 1322 2918 1774 2921
rect 1782 2921 1785 2928
rect 1782 2918 1918 2921
rect 1942 2921 1945 2928
rect 1942 2918 1982 2921
rect 2026 2918 2094 2921
rect 2114 2918 2390 2921
rect 2478 2921 2481 2928
rect 3222 2922 3225 2928
rect 2478 2918 2510 2921
rect 2586 2918 2726 2921
rect 2754 2918 3198 2921
rect 3234 2918 3294 2921
rect 3298 2918 3510 2921
rect 3570 2918 3646 2921
rect 3958 2921 3961 2928
rect 3866 2918 3961 2921
rect 4318 2922 4321 2928
rect 4374 2922 4377 2928
rect 4434 2918 4478 2921
rect 4482 2918 4489 2921
rect 4538 2918 4694 2921
rect 4698 2918 4814 2921
rect 4866 2918 4942 2921
rect 5010 2918 5254 2921
rect 4838 2912 4841 2918
rect 4854 2912 4857 2918
rect 306 2908 374 2911
rect 378 2908 454 2911
rect 538 2908 782 2911
rect 786 2908 814 2911
rect 1018 2908 1038 2911
rect 1046 2908 1262 2911
rect 1378 2908 1766 2911
rect 1914 2908 2118 2911
rect 2122 2908 2198 2911
rect 2354 2908 2534 2911
rect 2642 2908 2678 2911
rect 3058 2908 3246 2911
rect 3250 2908 3326 2911
rect 3362 2908 3838 2911
rect 3842 2908 3902 2911
rect 4306 2908 4414 2911
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 862 2903 864 2907
rect 210 2898 230 2901
rect 234 2898 342 2901
rect 450 2898 646 2901
rect 674 2898 718 2901
rect 914 2898 934 2901
rect 1046 2901 1049 2908
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1886 2903 1888 2907
rect 2888 2903 2890 2907
rect 2894 2903 2897 2907
rect 2902 2903 2904 2907
rect 3920 2903 3922 2907
rect 3926 2903 3929 2907
rect 3934 2903 3936 2907
rect 4936 2903 4938 2907
rect 4942 2903 4945 2907
rect 4950 2903 4952 2907
rect 938 2898 1049 2901
rect 1090 2898 1262 2901
rect 1306 2898 1478 2901
rect 1490 2898 1598 2901
rect 1714 2898 1798 2901
rect 1826 2898 1854 2901
rect 1914 2898 1998 2901
rect 2002 2898 2174 2901
rect 2306 2898 2326 2901
rect 2330 2898 2574 2901
rect 2602 2898 2606 2901
rect 2634 2898 2742 2901
rect 2914 2898 3550 2901
rect 3554 2898 3870 2901
rect 3970 2898 3998 2901
rect 4058 2898 4126 2901
rect 4130 2898 4190 2901
rect 4322 2898 4558 2901
rect 4562 2898 4590 2901
rect 4658 2898 4854 2901
rect 4858 2898 4878 2901
rect 5170 2898 5230 2901
rect 106 2888 297 2891
rect 294 2882 297 2888
rect 494 2888 534 2891
rect 558 2888 566 2891
rect 570 2888 590 2891
rect 598 2888 662 2891
rect 706 2888 806 2891
rect 814 2891 817 2898
rect 814 2888 942 2891
rect 1042 2888 1046 2891
rect 1074 2888 1078 2891
rect 1130 2888 1246 2891
rect 1250 2888 1326 2891
rect 1338 2888 1390 2891
rect 1770 2888 1862 2891
rect 2042 2888 2086 2891
rect 2090 2888 2102 2891
rect 2146 2888 2150 2891
rect 2178 2888 2214 2891
rect 2274 2888 2294 2891
rect 2482 2888 2574 2891
rect 2586 2888 2598 2891
rect 2602 2888 2609 2891
rect 2626 2888 2942 2891
rect 2946 2888 3030 2891
rect 3146 2888 3190 2891
rect 3194 2888 3238 2891
rect 3262 2888 3270 2891
rect 3274 2888 3350 2891
rect 3522 2888 3542 2891
rect 3554 2888 3646 2891
rect 3650 2888 3734 2891
rect 3858 2888 4022 2891
rect 4122 2888 4158 2891
rect 4178 2888 4230 2891
rect 4298 2888 4334 2891
rect 4954 2888 5118 2891
rect 494 2882 497 2888
rect 114 2878 182 2881
rect 298 2878 318 2881
rect 506 2878 574 2881
rect 598 2881 601 2888
rect 578 2878 601 2881
rect 618 2878 622 2881
rect 642 2878 678 2881
rect 682 2878 974 2881
rect 978 2878 998 2881
rect 1002 2878 1422 2881
rect 1442 2878 1510 2881
rect 1582 2881 1585 2888
rect 2342 2882 2345 2888
rect 1582 2878 1590 2881
rect 1754 2878 2038 2881
rect 2146 2878 2182 2881
rect 2186 2878 2278 2881
rect 2434 2878 2526 2881
rect 2562 2878 2638 2881
rect 2658 2878 3134 2881
rect 3138 2878 3654 2881
rect 3690 2878 3782 2881
rect 3906 2878 3990 2881
rect 4098 2878 4174 2881
rect 4178 2878 4286 2881
rect 4298 2878 4337 2881
rect 4538 2878 4566 2881
rect 4598 2881 4601 2888
rect 5166 2882 5169 2888
rect 4570 2878 4601 2881
rect 4802 2878 4862 2881
rect 5026 2878 5078 2881
rect 206 2872 209 2878
rect 1750 2872 1753 2878
rect 4334 2872 4337 2878
rect 114 2868 142 2871
rect 146 2868 158 2871
rect 274 2868 278 2871
rect 362 2868 366 2871
rect 450 2868 502 2871
rect 530 2868 534 2871
rect 586 2868 662 2871
rect 666 2868 734 2871
rect 874 2868 878 2871
rect 970 2868 1038 2871
rect 1138 2868 1190 2871
rect 1290 2868 1294 2871
rect 1306 2868 1310 2871
rect 1410 2868 1454 2871
rect 1626 2868 1702 2871
rect 1762 2868 1782 2871
rect 1802 2868 1894 2871
rect 1978 2868 2030 2871
rect 2074 2868 2254 2871
rect 2306 2868 2430 2871
rect 2858 2868 2966 2871
rect 3010 2868 3014 2871
rect 3098 2868 3174 2871
rect 3202 2868 3206 2871
rect 3322 2868 3334 2871
rect 3338 2868 3366 2871
rect 3498 2868 3526 2871
rect 3546 2868 3558 2871
rect 3594 2868 3782 2871
rect 3786 2868 3910 2871
rect 3914 2868 3998 2871
rect 4002 2868 4153 2871
rect 4158 2868 4166 2871
rect 4170 2868 4222 2871
rect 4546 2868 4574 2871
rect 4678 2868 4750 2871
rect 4890 2868 4990 2871
rect 5062 2868 5142 2871
rect 42 2858 46 2861
rect 146 2858 150 2861
rect 202 2858 350 2861
rect 354 2858 526 2861
rect 530 2858 558 2861
rect 562 2858 1054 2861
rect 1058 2858 1590 2861
rect 1594 2858 1766 2861
rect 1778 2858 2142 2861
rect 2146 2858 2150 2861
rect 2214 2858 2366 2861
rect 2510 2861 2513 2868
rect 2426 2858 2513 2861
rect 2542 2861 2545 2868
rect 2542 2858 2582 2861
rect 2590 2861 2593 2868
rect 2590 2858 2614 2861
rect 2622 2861 2625 2868
rect 2622 2858 2630 2861
rect 2658 2859 2662 2861
rect 2658 2858 2665 2859
rect 2778 2858 2782 2861
rect 2818 2858 2846 2861
rect 2850 2858 2870 2861
rect 2946 2858 3054 2861
rect 3058 2858 3126 2861
rect 3178 2858 3262 2861
rect 3282 2858 3302 2861
rect 3366 2858 3430 2861
rect 3582 2858 3622 2861
rect 3694 2858 3750 2861
rect 3802 2858 3830 2861
rect 3834 2858 3846 2861
rect 3986 2858 4014 2861
rect 4042 2858 4046 2861
rect 4150 2861 4153 2868
rect 4326 2862 4329 2868
rect 4526 2862 4529 2868
rect 4542 2862 4545 2868
rect 4678 2862 4681 2868
rect 4150 2858 4174 2861
rect 4194 2858 4310 2861
rect 4338 2858 4398 2861
rect 4478 2858 4486 2861
rect 4586 2858 4638 2861
rect 4786 2858 4806 2861
rect 4838 2861 4841 2868
rect 5062 2862 5065 2868
rect 5142 2862 5145 2868
rect 4834 2858 4846 2861
rect 4890 2858 4950 2861
rect 90 2848 190 2851
rect 194 2848 206 2851
rect 266 2848 278 2851
rect 370 2848 513 2851
rect 522 2848 534 2851
rect 538 2848 630 2851
rect 634 2848 646 2851
rect 738 2848 742 2851
rect 898 2848 918 2851
rect 930 2848 1078 2851
rect 1082 2848 1086 2851
rect 1098 2848 1102 2851
rect 1114 2848 1118 2851
rect 1290 2848 1294 2851
rect 1306 2848 1310 2851
rect 1394 2848 1438 2851
rect 1562 2848 1566 2851
rect 1698 2848 1734 2851
rect 1774 2848 1782 2851
rect 1786 2848 1830 2851
rect 2058 2848 2070 2851
rect 2082 2848 2110 2851
rect 2118 2848 2182 2851
rect 2186 2848 2190 2851
rect 2214 2851 2217 2858
rect 3366 2852 3369 2858
rect 3542 2852 3545 2858
rect 3582 2852 3585 2858
rect 3694 2852 3697 2858
rect 4478 2852 4481 2858
rect 2194 2848 2217 2851
rect 2250 2848 2294 2851
rect 2370 2848 2518 2851
rect 2858 2848 2926 2851
rect 3074 2848 3126 2851
rect 3146 2848 3190 2851
rect 3194 2848 3225 2851
rect 3266 2848 3318 2851
rect 3562 2848 3574 2851
rect 3834 2848 3846 2851
rect 3850 2848 4030 2851
rect 4050 2848 4238 2851
rect 4250 2848 4478 2851
rect 4794 2848 4798 2851
rect 4834 2848 4961 2851
rect 5210 2848 5214 2851
rect 5226 2848 5230 2851
rect 246 2842 249 2848
rect 510 2842 513 2848
rect 106 2838 198 2841
rect 258 2838 310 2841
rect 314 2838 358 2841
rect 394 2838 398 2841
rect 546 2838 598 2841
rect 618 2838 710 2841
rect 846 2838 854 2841
rect 858 2838 902 2841
rect 930 2838 1150 2841
rect 1154 2838 1158 2841
rect 1162 2838 1382 2841
rect 1386 2838 1438 2841
rect 1570 2838 1942 2841
rect 1978 2838 2065 2841
rect 2118 2841 2121 2848
rect 2766 2842 2769 2848
rect 3222 2842 3225 2848
rect 4958 2842 4961 2848
rect 2074 2838 2121 2841
rect 2138 2838 2310 2841
rect 3330 2838 3366 2841
rect 3466 2838 3622 2841
rect 3626 2838 3782 2841
rect 3858 2838 3998 2841
rect 4122 2838 4510 2841
rect 4514 2838 4718 2841
rect 5090 2838 5214 2841
rect 2062 2832 2065 2838
rect 114 2828 134 2831
rect 386 2828 566 2831
rect 570 2828 598 2831
rect 826 2828 886 2831
rect 890 2828 966 2831
rect 970 2828 1134 2831
rect 1138 2828 1206 2831
rect 1210 2828 1310 2831
rect 1426 2828 1534 2831
rect 1682 2828 1686 2831
rect 2122 2828 2342 2831
rect 2674 2828 2846 2831
rect 3050 2828 3166 2831
rect 3274 2828 3334 2831
rect 3354 2828 4206 2831
rect 4774 2831 4777 2838
rect 4250 2828 4777 2831
rect 4946 2828 5078 2831
rect 5250 2828 5286 2831
rect 186 2818 534 2821
rect 690 2818 1542 2821
rect 1546 2818 1806 2821
rect 1810 2818 2094 2821
rect 2098 2818 2425 2821
rect 2466 2818 2470 2821
rect 2530 2818 2654 2821
rect 2690 2818 2942 2821
rect 3122 2818 3462 2821
rect 3498 2818 3534 2821
rect 3538 2818 3558 2821
rect 3794 2818 4134 2821
rect 4282 2818 4462 2821
rect 4502 2818 4510 2821
rect 4514 2818 4646 2821
rect 5026 2818 5038 2821
rect 5042 2818 5086 2821
rect 5202 2818 5222 2821
rect 394 2808 638 2811
rect 690 2808 694 2811
rect 706 2808 766 2811
rect 770 2808 958 2811
rect 962 2808 1118 2811
rect 1146 2808 1334 2811
rect 1410 2808 1422 2811
rect 1522 2808 1585 2811
rect 1674 2808 1726 2811
rect 1746 2808 1822 2811
rect 1826 2808 1934 2811
rect 1938 2808 2086 2811
rect 2098 2808 2134 2811
rect 2218 2808 2310 2811
rect 2422 2811 2425 2818
rect 5286 2812 5289 2818
rect 2422 2808 2462 2811
rect 2538 2808 3030 2811
rect 3106 2808 3110 2811
rect 3114 2808 3390 2811
rect 3426 2808 3966 2811
rect 3974 2808 4350 2811
rect 4490 2808 5054 2811
rect 328 2803 330 2807
rect 334 2803 337 2807
rect 342 2803 344 2807
rect 474 2798 558 2801
rect 562 2798 630 2801
rect 702 2801 705 2808
rect 1352 2803 1354 2807
rect 1358 2803 1361 2807
rect 1366 2803 1368 2807
rect 634 2798 705 2801
rect 826 2798 894 2801
rect 906 2798 982 2801
rect 1098 2798 1142 2801
rect 1162 2798 1214 2801
rect 1582 2801 1585 2808
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2398 2803 2400 2807
rect 2406 2802 2409 2808
rect 3400 2803 3402 2807
rect 3406 2803 3409 2807
rect 3414 2803 3416 2807
rect 1582 2798 1742 2801
rect 1762 2798 1814 2801
rect 1930 2798 2094 2801
rect 2106 2798 2214 2801
rect 2490 2798 2502 2801
rect 2706 2798 2966 2801
rect 2970 2798 3006 2801
rect 3018 2798 3278 2801
rect 3626 2798 3638 2801
rect 3974 2801 3977 2808
rect 4424 2803 4426 2807
rect 4430 2803 4433 2807
rect 4438 2803 4440 2807
rect 3698 2798 3977 2801
rect 3994 2798 3998 2801
rect 4130 2798 4166 2801
rect 4810 2798 5110 2801
rect 5162 2798 5174 2801
rect 498 2788 574 2791
rect 698 2788 702 2791
rect 722 2788 822 2791
rect 834 2788 1070 2791
rect 1090 2788 1102 2791
rect 1106 2788 1398 2791
rect 1602 2788 1758 2791
rect 1842 2788 2454 2791
rect 2458 2788 2958 2791
rect 2994 2788 3286 2791
rect 3306 2788 3478 2791
rect 4122 2788 4198 2791
rect 4578 2788 4614 2791
rect 4714 2788 4830 2791
rect 5058 2788 5102 2791
rect 5242 2788 5254 2791
rect 1574 2782 1577 2788
rect 3038 2782 3041 2788
rect 346 2778 382 2781
rect 506 2778 582 2781
rect 618 2778 1398 2781
rect 1410 2778 1550 2781
rect 1738 2778 2006 2781
rect 2114 2778 2262 2781
rect 2274 2778 2654 2781
rect 2658 2778 2750 2781
rect 2794 2778 2822 2781
rect 3002 2778 3014 2781
rect 3074 2778 3334 2781
rect 3338 2778 3638 2781
rect 3658 2778 3910 2781
rect 4034 2778 4222 2781
rect 4226 2778 4598 2781
rect 4602 2778 4670 2781
rect 4882 2778 5062 2781
rect 5074 2778 5134 2781
rect 290 2768 1174 2771
rect 1178 2768 1270 2771
rect 1298 2768 1454 2771
rect 1514 2768 1574 2771
rect 1578 2768 1582 2771
rect 1642 2768 1718 2771
rect 2130 2768 2142 2771
rect 2146 2768 2153 2771
rect 2162 2768 2174 2771
rect 2210 2768 2286 2771
rect 2290 2768 2382 2771
rect 2482 2768 2486 2771
rect 2562 2768 2678 2771
rect 2682 2768 2782 2771
rect 2786 2768 2806 2771
rect 2850 2768 2926 2771
rect 3026 2768 3718 2771
rect 3786 2768 4022 2771
rect 4042 2768 4062 2771
rect 4066 2768 4126 2771
rect 4234 2768 4238 2771
rect 4354 2768 4561 2771
rect 4586 2768 4622 2771
rect 4698 2768 4710 2771
rect 4738 2768 4790 2771
rect 4858 2768 4870 2771
rect 4922 2768 4974 2771
rect 4978 2768 5038 2771
rect 5090 2768 5126 2771
rect 514 2758 550 2761
rect 646 2758 654 2761
rect 658 2758 726 2761
rect 858 2758 937 2761
rect 946 2758 950 2761
rect 962 2758 966 2761
rect 970 2758 990 2761
rect 1010 2758 1086 2761
rect 1122 2758 1126 2761
rect 1154 2758 1158 2761
rect 1354 2758 1478 2761
rect 1482 2758 1502 2761
rect 2038 2761 2041 2768
rect 1562 2758 2041 2761
rect 2090 2758 2270 2761
rect 2294 2758 2494 2761
rect 2502 2761 2505 2768
rect 2502 2758 2534 2761
rect 2610 2758 2862 2761
rect 2866 2758 2870 2761
rect 2882 2758 2926 2761
rect 2938 2758 2950 2761
rect 2962 2758 2966 2761
rect 3474 2758 3494 2761
rect 3570 2758 3606 2761
rect 3714 2758 3758 2761
rect 3770 2758 3798 2761
rect 3810 2758 3846 2761
rect 3866 2758 3958 2761
rect 4050 2758 4086 2761
rect 4202 2758 4302 2761
rect 4334 2761 4337 2768
rect 4306 2758 4337 2761
rect 4558 2762 4561 2768
rect 4686 2761 4689 2768
rect 4578 2758 4689 2761
rect 4754 2758 4758 2761
rect 4762 2758 4894 2761
rect 4906 2758 4926 2761
rect 5018 2758 5086 2761
rect 50 2748 118 2751
rect 130 2748 254 2751
rect 290 2748 390 2751
rect 566 2751 569 2758
rect 934 2752 937 2758
rect 530 2748 569 2751
rect 594 2748 598 2751
rect 618 2748 622 2751
rect 642 2748 710 2751
rect 714 2748 718 2751
rect 738 2748 742 2751
rect 818 2748 897 2751
rect 906 2748 929 2751
rect 1074 2748 1134 2751
rect 1190 2751 1193 2758
rect 1154 2748 1193 2751
rect 1442 2748 1462 2751
rect 1466 2748 1502 2751
rect 1542 2751 1545 2758
rect 2294 2752 2297 2758
rect 2494 2752 2497 2758
rect 3166 2752 3169 2758
rect 1542 2748 1558 2751
rect 1570 2748 1662 2751
rect 1722 2748 1950 2751
rect 1962 2748 2134 2751
rect 2146 2748 2150 2751
rect 2242 2748 2246 2751
rect 2514 2748 2550 2751
rect 2642 2748 2750 2751
rect 2754 2748 2777 2751
rect 2794 2748 2798 2751
rect 2882 2748 2918 2751
rect 2954 2748 2958 2751
rect 3074 2748 3102 2751
rect 3106 2748 3150 2751
rect 3210 2748 3238 2751
rect 3242 2748 3262 2751
rect 3302 2751 3305 2758
rect 4110 2752 4113 2758
rect 4174 2752 4177 2758
rect 3302 2748 3390 2751
rect 3426 2748 3510 2751
rect 3522 2748 3894 2751
rect 3898 2748 3950 2751
rect 4026 2748 4046 2751
rect 4090 2748 4094 2751
rect 4098 2748 4102 2751
rect 4186 2748 4310 2751
rect 4314 2748 4390 2751
rect 4442 2748 4478 2751
rect 4594 2748 4766 2751
rect 4786 2748 4790 2751
rect 4906 2748 4910 2751
rect 4922 2748 4926 2751
rect 5026 2748 5166 2751
rect 5170 2748 5198 2751
rect 5218 2748 5238 2751
rect 5334 2751 5338 2752
rect 5282 2748 5338 2751
rect 66 2738 161 2741
rect 270 2741 273 2748
rect 894 2742 897 2748
rect 926 2742 929 2748
rect 1734 2742 1737 2748
rect 2774 2742 2777 2748
rect 226 2738 273 2741
rect 314 2738 406 2741
rect 410 2738 518 2741
rect 522 2738 694 2741
rect 718 2738 734 2741
rect 742 2738 878 2741
rect 1074 2738 1078 2741
rect 1434 2738 1486 2741
rect 1578 2738 1694 2741
rect 1770 2738 1806 2741
rect 1842 2738 1886 2741
rect 2042 2738 2094 2741
rect 2122 2738 2134 2741
rect 2202 2738 2246 2741
rect 2266 2738 2270 2741
rect 2282 2738 2342 2741
rect 2450 2738 2606 2741
rect 2634 2738 2678 2741
rect 2794 2738 3102 2741
rect 3154 2738 3166 2741
rect 3474 2738 3574 2741
rect 3722 2738 4334 2741
rect 4338 2738 4382 2741
rect 4414 2741 4417 2748
rect 4414 2738 4478 2741
rect 4554 2738 4582 2741
rect 4658 2738 4662 2741
rect 5022 2741 5025 2748
rect 4690 2738 5025 2741
rect 5066 2738 5126 2741
rect 5202 2738 5254 2741
rect 158 2732 161 2738
rect 718 2732 721 2738
rect 742 2732 745 2738
rect 1102 2732 1105 2738
rect 1110 2732 1113 2738
rect 458 2728 542 2731
rect 554 2728 630 2731
rect 794 2728 918 2731
rect 1178 2728 1366 2731
rect 1378 2728 1438 2731
rect 1442 2728 1454 2731
rect 1546 2728 1606 2731
rect 1702 2731 1705 2738
rect 1758 2732 1761 2738
rect 1702 2728 1750 2731
rect 1830 2728 1833 2738
rect 2886 2732 2889 2738
rect 3358 2732 3361 2738
rect 1854 2728 1862 2731
rect 1866 2728 1942 2731
rect 1994 2728 2070 2731
rect 2258 2728 2574 2731
rect 2578 2728 2598 2731
rect 2618 2728 2622 2731
rect 2738 2728 2862 2731
rect 2978 2728 3342 2731
rect 3394 2728 3542 2731
rect 3546 2728 3678 2731
rect 3802 2728 3806 2731
rect 3882 2728 3886 2731
rect 3946 2728 3974 2731
rect 4082 2728 4097 2731
rect 4234 2728 4286 2731
rect 4314 2728 4374 2731
rect 4458 2728 4566 2731
rect 4570 2728 4790 2731
rect 4794 2728 4862 2731
rect 4922 2728 4950 2731
rect 4970 2728 5030 2731
rect 5042 2728 5086 2731
rect 306 2718 318 2721
rect 386 2718 798 2721
rect 866 2718 942 2721
rect 1114 2718 1118 2721
rect 1126 2721 1129 2728
rect 1126 2718 1150 2721
rect 1162 2718 1190 2721
rect 1410 2718 1422 2721
rect 1426 2718 1486 2721
rect 1506 2718 1566 2721
rect 1586 2718 1590 2721
rect 1698 2718 1774 2721
rect 1906 2718 1998 2721
rect 2074 2718 2142 2721
rect 2178 2718 2182 2721
rect 2482 2718 2510 2721
rect 2546 2718 2574 2721
rect 2594 2718 2598 2721
rect 2610 2718 2814 2721
rect 2818 2718 3174 2721
rect 3178 2718 3742 2721
rect 3750 2721 3753 2728
rect 4094 2722 4097 2728
rect 3746 2718 3753 2721
rect 3762 2718 3902 2721
rect 4242 2718 4262 2721
rect 4330 2718 4334 2721
rect 4386 2718 4414 2721
rect 4446 2721 4449 2728
rect 4418 2718 4449 2721
rect 4766 2718 4774 2721
rect 4778 2718 4854 2721
rect 4962 2718 5062 2721
rect 5066 2718 5238 2721
rect 2582 2712 2585 2718
rect 4742 2712 4745 2718
rect 186 2708 246 2711
rect 250 2708 318 2711
rect 322 2708 366 2711
rect 370 2708 590 2711
rect 602 2708 790 2711
rect 1058 2708 1174 2711
rect 1202 2708 1254 2711
rect 1258 2708 1401 2711
rect 1426 2708 1430 2711
rect 1538 2708 1590 2711
rect 1602 2708 1654 2711
rect 2034 2708 2190 2711
rect 2226 2708 2518 2711
rect 2594 2708 2742 2711
rect 2810 2708 2878 2711
rect 2922 2708 2966 2711
rect 2970 2708 2998 2711
rect 3138 2708 3446 2711
rect 3482 2708 3502 2711
rect 3690 2708 3742 2711
rect 3978 2708 4062 2711
rect 4082 2708 4270 2711
rect 4274 2708 4302 2711
rect 4410 2708 4470 2711
rect 4642 2708 4670 2711
rect 4866 2708 4870 2711
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 862 2703 864 2707
rect 274 2698 350 2701
rect 354 2698 430 2701
rect 594 2698 606 2701
rect 618 2698 774 2701
rect 906 2698 990 2701
rect 1146 2698 1390 2701
rect 1398 2701 1401 2708
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1886 2703 1888 2707
rect 2888 2703 2890 2707
rect 2894 2703 2897 2707
rect 2902 2703 2904 2707
rect 3920 2703 3922 2707
rect 3926 2703 3929 2707
rect 3934 2703 3936 2707
rect 4918 2702 4921 2708
rect 4936 2703 4938 2707
rect 4942 2703 4945 2707
rect 4950 2703 4952 2707
rect 1398 2698 1734 2701
rect 2050 2698 2070 2701
rect 2174 2698 2246 2701
rect 2362 2698 2478 2701
rect 2482 2698 2550 2701
rect 2562 2698 2582 2701
rect 2618 2698 2638 2701
rect 2682 2698 2854 2701
rect 3034 2698 3150 2701
rect 3154 2698 3238 2701
rect 3250 2698 3590 2701
rect 3626 2698 3822 2701
rect 3826 2698 3854 2701
rect 4002 2698 4126 2701
rect 4146 2698 4278 2701
rect 4330 2698 4894 2701
rect 94 2688 150 2691
rect 482 2688 486 2691
rect 550 2688 558 2691
rect 562 2688 582 2691
rect 634 2688 638 2691
rect 858 2688 926 2691
rect 1070 2688 1118 2691
rect 1154 2688 1166 2691
rect 1274 2688 1334 2691
rect 1482 2688 1526 2691
rect 1530 2688 1574 2691
rect 1650 2688 1654 2691
rect 1666 2688 1753 2691
rect 1786 2688 1838 2691
rect 2174 2691 2177 2698
rect 1938 2688 2177 2691
rect 2330 2688 2606 2691
rect 2754 2688 2838 2691
rect 3034 2688 3326 2691
rect 3666 2688 3686 2691
rect 3722 2688 3766 2691
rect 3890 2688 3950 2691
rect 3954 2688 4118 2691
rect 4122 2688 4134 2691
rect 4138 2688 4398 2691
rect 4466 2688 4470 2691
rect 4530 2688 4582 2691
rect 4626 2688 4686 2691
rect 4786 2688 4910 2691
rect 94 2682 97 2688
rect 1070 2682 1073 2688
rect 1750 2682 1753 2688
rect 2182 2682 2185 2688
rect 202 2678 230 2681
rect 242 2678 254 2681
rect 434 2678 886 2681
rect 938 2678 1025 2681
rect 1082 2678 1126 2681
rect 1130 2678 1518 2681
rect 1522 2678 1710 2681
rect 2002 2678 2030 2681
rect 2042 2678 2046 2681
rect 2066 2678 2110 2681
rect 2242 2678 2286 2681
rect 2670 2681 2673 2688
rect 2990 2682 2993 2688
rect 2522 2678 2673 2681
rect 2690 2678 2766 2681
rect 3158 2678 3214 2681
rect 3218 2678 3254 2681
rect 3314 2678 3454 2681
rect 3494 2681 3497 2688
rect 4278 2682 4281 2688
rect 3458 2678 3497 2681
rect 3510 2678 3518 2681
rect 3522 2678 3670 2681
rect 3674 2678 3798 2681
rect 3866 2678 3894 2681
rect 3954 2678 3966 2681
rect 4042 2678 4150 2681
rect 4194 2678 4198 2681
rect 4410 2678 4550 2681
rect 4758 2681 4761 2688
rect 4586 2678 4761 2681
rect 4906 2678 4998 2681
rect 5082 2678 5086 2681
rect 130 2668 134 2671
rect 270 2671 273 2678
rect 270 2668 350 2671
rect 422 2671 425 2678
rect 1022 2672 1025 2678
rect 3158 2672 3161 2678
rect 422 2668 518 2671
rect 538 2668 590 2671
rect 650 2668 673 2671
rect 714 2668 718 2671
rect 738 2668 758 2671
rect 954 2668 966 2671
rect 1066 2668 1086 2671
rect 1090 2668 1118 2671
rect 1130 2668 1142 2671
rect 1170 2668 1206 2671
rect 1210 2668 1326 2671
rect 1338 2668 1350 2671
rect 1386 2668 1598 2671
rect 1626 2668 1686 2671
rect 1706 2668 1830 2671
rect 1834 2668 1862 2671
rect 1874 2668 1926 2671
rect 2018 2668 2046 2671
rect 2098 2668 2134 2671
rect 2154 2668 2678 2671
rect 2682 2668 2982 2671
rect 2994 2668 3022 2671
rect 3498 2668 3518 2671
rect 3602 2668 3606 2671
rect 3730 2668 3734 2671
rect 3738 2668 3750 2671
rect 3830 2671 3833 2678
rect 4262 2672 4265 2678
rect 4390 2672 4393 2678
rect 3818 2668 3833 2671
rect 3890 2668 3934 2671
rect 3938 2668 3958 2671
rect 3978 2668 4014 2671
rect 4362 2668 4374 2671
rect 4538 2668 4550 2671
rect 4554 2668 4662 2671
rect 4838 2671 4841 2678
rect 4834 2668 4841 2671
rect 4914 2668 4942 2671
rect 110 2662 113 2668
rect 50 2658 86 2661
rect 130 2658 166 2661
rect 218 2658 230 2661
rect 250 2658 254 2661
rect 258 2658 286 2661
rect 422 2661 425 2668
rect 290 2658 425 2661
rect 442 2658 481 2661
rect 578 2658 582 2661
rect 594 2658 662 2661
rect 670 2661 673 2668
rect 726 2661 729 2668
rect 814 2662 817 2668
rect 830 2662 833 2668
rect 670 2658 729 2661
rect 762 2658 766 2661
rect 850 2658 910 2661
rect 914 2658 1086 2661
rect 1098 2658 1102 2661
rect 1106 2658 1134 2661
rect 1138 2658 1302 2661
rect 1410 2658 1414 2661
rect 1450 2659 1510 2661
rect 1450 2658 1513 2659
rect 1610 2658 1694 2661
rect 1762 2658 1782 2661
rect 1794 2658 1814 2661
rect 1842 2658 1998 2661
rect 2058 2658 2062 2661
rect 2082 2658 2102 2661
rect 2114 2658 2118 2661
rect 2170 2658 2182 2661
rect 2234 2658 2238 2661
rect 2266 2658 2702 2661
rect 2706 2658 2718 2661
rect 2898 2658 2990 2661
rect 3010 2658 3078 2661
rect 3158 2661 3161 2668
rect 3138 2658 3161 2661
rect 3266 2658 3294 2661
rect 3318 2661 3321 2668
rect 3298 2658 3321 2661
rect 3538 2658 3542 2661
rect 3562 2658 3590 2661
rect 3614 2661 3617 2668
rect 3594 2658 3617 2661
rect 3642 2658 3646 2661
rect 3654 2658 3657 2668
rect 3790 2662 3793 2668
rect 3666 2658 3670 2661
rect 3674 2658 3782 2661
rect 3834 2658 3862 2661
rect 4134 2661 4137 2668
rect 4214 2662 4217 2668
rect 3874 2658 4105 2661
rect 4134 2658 4166 2661
rect 4342 2661 4345 2668
rect 4314 2658 4345 2661
rect 4350 2662 4353 2668
rect 4534 2662 4537 2668
rect 4878 2662 4881 2668
rect 4354 2658 4366 2661
rect 4458 2658 4462 2661
rect 4506 2658 4510 2661
rect 4634 2658 4678 2661
rect 4770 2658 4774 2661
rect 4882 2658 5014 2661
rect 5090 2658 5142 2661
rect 110 2651 113 2658
rect 478 2652 481 2658
rect 1710 2652 1713 2658
rect 3998 2652 4001 2658
rect 4102 2652 4105 2658
rect 110 2648 430 2651
rect 554 2648 558 2651
rect 610 2648 758 2651
rect 810 2648 838 2651
rect 922 2648 1046 2651
rect 1074 2648 1406 2651
rect 1450 2648 1566 2651
rect 1570 2648 1630 2651
rect 1826 2648 2070 2651
rect 2074 2648 2150 2651
rect 2162 2648 2166 2651
rect 2202 2648 2254 2651
rect 2258 2648 2286 2651
rect 2310 2648 2318 2651
rect 2322 2648 2422 2651
rect 2474 2648 2518 2651
rect 2726 2648 2734 2651
rect 2738 2648 2782 2651
rect 2802 2648 2966 2651
rect 2970 2648 3454 2651
rect 3474 2648 3750 2651
rect 3858 2648 3921 2651
rect 4138 2648 4190 2651
rect 4266 2648 4318 2651
rect 4338 2648 4342 2651
rect 4394 2648 4414 2651
rect 4458 2648 4526 2651
rect 4530 2648 4686 2651
rect 4730 2648 4814 2651
rect 4830 2648 4838 2651
rect 4926 2648 4934 2651
rect 4938 2648 5038 2651
rect 5242 2648 5246 2651
rect 5334 2648 5338 2652
rect 274 2638 382 2641
rect 386 2638 406 2641
rect 450 2638 486 2641
rect 506 2638 550 2641
rect 554 2638 566 2641
rect 714 2638 742 2641
rect 766 2641 769 2648
rect 746 2638 769 2641
rect 906 2638 926 2641
rect 1090 2638 1102 2641
rect 1106 2638 1182 2641
rect 1186 2638 1342 2641
rect 1346 2638 1350 2641
rect 1354 2638 1422 2641
rect 1514 2638 1790 2641
rect 2002 2638 2078 2641
rect 2090 2638 2326 2641
rect 2362 2638 2446 2641
rect 2450 2638 2502 2641
rect 2626 2638 2646 2641
rect 2650 2638 2902 2641
rect 2942 2638 2950 2641
rect 2954 2638 3038 2641
rect 3066 2638 3150 2641
rect 3154 2638 3310 2641
rect 3386 2638 3430 2641
rect 3434 2638 3486 2641
rect 3538 2638 3542 2641
rect 3610 2638 3750 2641
rect 3754 2638 3878 2641
rect 3918 2641 3921 2648
rect 3918 2638 4062 2641
rect 4066 2638 4174 2641
rect 5334 2641 5337 2648
rect 4306 2638 5337 2641
rect 698 2628 718 2631
rect 786 2628 1086 2631
rect 1114 2628 1142 2631
rect 1418 2628 1478 2631
rect 1482 2628 1526 2631
rect 1586 2628 1758 2631
rect 1770 2628 1782 2631
rect 1794 2628 1822 2631
rect 2098 2628 2126 2631
rect 2154 2628 2190 2631
rect 2346 2628 2566 2631
rect 2602 2628 2766 2631
rect 2810 2628 3222 2631
rect 3458 2628 3830 2631
rect 4026 2628 4062 2631
rect 4162 2628 4302 2631
rect 4306 2628 4313 2631
rect 4322 2628 4702 2631
rect 4866 2628 4942 2631
rect 2310 2622 2313 2628
rect 122 2618 134 2621
rect 138 2618 142 2621
rect 146 2618 390 2621
rect 394 2618 614 2621
rect 618 2618 670 2621
rect 794 2618 822 2621
rect 1306 2618 1318 2621
rect 1322 2618 1470 2621
rect 1474 2618 1542 2621
rect 1662 2618 1670 2621
rect 1674 2618 1902 2621
rect 1922 2618 1966 2621
rect 2138 2618 2214 2621
rect 2626 2618 2734 2621
rect 2770 2618 2822 2621
rect 2826 2618 2886 2621
rect 2954 2618 2990 2621
rect 3130 2618 3366 2621
rect 3398 2621 3401 2628
rect 3398 2618 3422 2621
rect 3506 2618 3622 2621
rect 3738 2618 4022 2621
rect 4106 2618 4358 2621
rect 4362 2618 4374 2621
rect 4714 2618 5102 2621
rect 426 2608 614 2611
rect 618 2608 1070 2611
rect 1426 2608 1566 2611
rect 1594 2608 1774 2611
rect 1778 2608 1806 2611
rect 1882 2608 1926 2611
rect 1930 2608 1990 2611
rect 2178 2608 2190 2611
rect 2226 2608 2238 2611
rect 2466 2608 2486 2611
rect 2570 2608 2574 2611
rect 2586 2608 2822 2611
rect 2826 2608 3198 2611
rect 3498 2608 3702 2611
rect 3786 2608 3814 2611
rect 3818 2608 4206 2611
rect 4530 2608 4718 2611
rect 4770 2608 5198 2611
rect 328 2603 330 2607
rect 334 2603 337 2607
rect 342 2603 344 2607
rect 1352 2603 1354 2607
rect 1358 2603 1361 2607
rect 1366 2603 1368 2607
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2398 2603 2400 2607
rect 3400 2603 3402 2607
rect 3406 2603 3409 2607
rect 3414 2603 3416 2607
rect 3750 2602 3753 2608
rect 4424 2603 4426 2607
rect 4430 2603 4433 2607
rect 4438 2603 4440 2607
rect 4470 2602 4473 2608
rect 570 2598 846 2601
rect 1402 2598 1622 2601
rect 1690 2598 1750 2601
rect 1754 2598 1830 2601
rect 2074 2598 2078 2601
rect 2098 2598 2174 2601
rect 2242 2598 2334 2601
rect 2682 2598 2782 2601
rect 2922 2598 3054 2601
rect 3066 2598 3174 2601
rect 3178 2598 3390 2601
rect 3554 2598 3558 2601
rect 3570 2598 3718 2601
rect 4154 2598 4318 2601
rect 4506 2598 4598 2601
rect 4690 2598 4838 2601
rect 4842 2598 4902 2601
rect 4906 2598 4990 2601
rect 162 2588 182 2591
rect 266 2588 294 2591
rect 298 2588 2022 2591
rect 2026 2588 2598 2591
rect 2602 2588 3214 2591
rect 3226 2588 3686 2591
rect 3714 2588 3862 2591
rect 4042 2588 4110 2591
rect 4186 2588 4230 2591
rect 4402 2588 4638 2591
rect 4642 2588 4798 2591
rect 5090 2588 5158 2591
rect 4382 2582 4385 2588
rect 90 2578 134 2581
rect 362 2578 486 2581
rect 722 2578 830 2581
rect 1098 2578 1982 2581
rect 1986 2578 4254 2581
rect 4274 2578 4310 2581
rect 4314 2578 4342 2581
rect 4458 2578 4609 2581
rect 4618 2578 4622 2581
rect 4722 2578 4790 2581
rect 3294 2572 3297 2578
rect 4606 2572 4609 2578
rect 266 2568 297 2571
rect 306 2568 326 2571
rect 362 2568 446 2571
rect 714 2568 734 2571
rect 738 2568 801 2571
rect 110 2561 113 2568
rect 42 2558 113 2561
rect 126 2561 129 2568
rect 150 2561 153 2568
rect 294 2562 297 2568
rect 798 2562 801 2568
rect 842 2568 870 2571
rect 882 2568 926 2571
rect 978 2568 1009 2571
rect 1018 2568 1078 2571
rect 1146 2568 1222 2571
rect 1294 2568 1518 2571
rect 1530 2568 1534 2571
rect 1706 2568 2094 2571
rect 2138 2568 2198 2571
rect 2274 2568 2286 2571
rect 2442 2568 2926 2571
rect 2930 2568 2974 2571
rect 3002 2568 3174 2571
rect 3386 2568 3478 2571
rect 3482 2568 3550 2571
rect 3554 2568 3582 2571
rect 3778 2568 3790 2571
rect 3970 2568 4601 2571
rect 4618 2568 4806 2571
rect 4922 2568 5014 2571
rect 5018 2568 5094 2571
rect 5162 2568 5166 2571
rect 126 2558 153 2561
rect 202 2558 278 2561
rect 370 2558 374 2561
rect 466 2558 470 2561
rect 814 2561 817 2568
rect 830 2561 833 2568
rect 1006 2562 1009 2568
rect 1294 2562 1297 2568
rect 2254 2562 2257 2568
rect 814 2558 833 2561
rect 850 2558 870 2561
rect 914 2558 990 2561
rect 1066 2558 1113 2561
rect 1138 2558 1142 2561
rect 1146 2558 1150 2561
rect 1314 2558 1382 2561
rect 1386 2558 1430 2561
rect 1530 2558 1558 2561
rect 1562 2558 1566 2561
rect 1626 2558 1694 2561
rect 1762 2558 1766 2561
rect 1898 2558 1918 2561
rect 2082 2558 2086 2561
rect 2114 2558 2182 2561
rect 2210 2558 2238 2561
rect 2402 2558 2406 2561
rect 2426 2558 2446 2561
rect 2450 2558 2558 2561
rect 2578 2558 2726 2561
rect 2762 2558 2766 2561
rect 2794 2558 2894 2561
rect 2914 2558 2974 2561
rect 3034 2558 3070 2561
rect 3090 2558 3206 2561
rect 3250 2558 3254 2561
rect 3314 2558 3342 2561
rect 3346 2558 3374 2561
rect 3378 2558 3406 2561
rect 3750 2561 3753 2568
rect 3418 2558 3753 2561
rect 3774 2558 3846 2561
rect 4178 2558 4398 2561
rect 4446 2558 4486 2561
rect 4490 2558 4590 2561
rect 4598 2561 4601 2568
rect 4598 2558 4766 2561
rect 4770 2558 4790 2561
rect 4818 2558 4886 2561
rect 4914 2558 4990 2561
rect 5122 2558 5126 2561
rect 5194 2558 5262 2561
rect 114 2548 118 2551
rect 122 2548 214 2551
rect 274 2548 278 2551
rect 378 2548 406 2551
rect 442 2548 654 2551
rect 666 2548 974 2551
rect 1110 2551 1113 2558
rect 978 2548 1105 2551
rect 1110 2548 1198 2551
rect 1330 2548 1334 2551
rect 1418 2548 1422 2551
rect 1538 2548 1585 2551
rect 1594 2548 1614 2551
rect 1662 2548 1726 2551
rect 1974 2551 1977 2558
rect 1802 2548 1977 2551
rect 2002 2548 2142 2551
rect 2186 2548 2222 2551
rect 2226 2548 2254 2551
rect 2562 2548 2590 2551
rect 2658 2548 2662 2551
rect 2666 2548 2673 2551
rect 2706 2548 2718 2551
rect 2726 2551 2729 2558
rect 3022 2552 3025 2558
rect 2726 2548 2782 2551
rect 2794 2548 2798 2551
rect 2850 2548 2886 2551
rect 2890 2548 2902 2551
rect 2954 2548 2958 2551
rect 2986 2548 3001 2551
rect 3010 2548 3014 2551
rect 3090 2548 3118 2551
rect 3130 2548 3190 2551
rect 3194 2548 3201 2551
rect 3242 2548 3246 2551
rect 3250 2548 3382 2551
rect 3774 2551 3777 2558
rect 3394 2548 3777 2551
rect 3786 2548 3790 2551
rect 3818 2548 3822 2551
rect 3914 2548 3974 2551
rect 4058 2548 4070 2551
rect 4122 2548 4126 2551
rect 4134 2551 4137 2558
rect 4446 2552 4449 2558
rect 4134 2548 4158 2551
rect 4402 2548 4446 2551
rect 4458 2548 4465 2551
rect 4522 2548 4542 2551
rect 4618 2548 4878 2551
rect 4882 2548 4926 2551
rect 4962 2548 5046 2551
rect 5146 2548 5214 2551
rect 5334 2551 5338 2552
rect 5250 2548 5338 2551
rect 1102 2542 1105 2548
rect 162 2538 190 2541
rect 258 2538 350 2541
rect 490 2538 566 2541
rect 770 2538 830 2541
rect 846 2538 1030 2541
rect 1058 2538 1062 2541
rect 1130 2538 1166 2541
rect 1178 2538 1190 2541
rect 1194 2538 1206 2541
rect 1210 2538 1254 2541
rect 1266 2538 1342 2541
rect 1490 2538 1566 2541
rect 1582 2541 1585 2548
rect 1662 2542 1665 2548
rect 2718 2542 2721 2548
rect 1582 2538 1630 2541
rect 1722 2538 1838 2541
rect 1842 2538 1910 2541
rect 2218 2538 2302 2541
rect 2306 2538 2422 2541
rect 2498 2538 2582 2541
rect 2786 2538 2838 2541
rect 2842 2538 2926 2541
rect 2986 2538 2990 2541
rect 2998 2541 3001 2548
rect 3078 2542 3081 2548
rect 3126 2542 3129 2548
rect 4462 2542 4465 2548
rect 2998 2538 3014 2541
rect 3034 2538 3046 2541
rect 3106 2538 3110 2541
rect 3162 2538 3166 2541
rect 3178 2538 3214 2541
rect 3258 2538 3310 2541
rect 3490 2538 3518 2541
rect 3554 2538 3566 2541
rect 3642 2538 3678 2541
rect 3682 2538 3702 2541
rect 3706 2538 3734 2541
rect 3738 2538 3774 2541
rect 3810 2538 3870 2541
rect 3882 2538 3958 2541
rect 4154 2538 4174 2541
rect 4354 2538 4398 2541
rect 4426 2538 4430 2541
rect 4610 2538 4614 2541
rect 4674 2538 4710 2541
rect 4874 2538 4966 2541
rect 4994 2538 5094 2541
rect 5242 2538 5246 2541
rect 106 2528 262 2531
rect 298 2528 318 2531
rect 418 2528 470 2531
rect 554 2528 630 2531
rect 634 2528 750 2531
rect 754 2528 806 2531
rect 846 2531 849 2538
rect 1446 2532 1449 2538
rect 1942 2532 1945 2538
rect 826 2528 849 2531
rect 858 2528 974 2531
rect 978 2528 1217 2531
rect 1258 2528 1334 2531
rect 1338 2528 1366 2531
rect 1554 2528 1590 2531
rect 1778 2528 1894 2531
rect 1906 2528 1918 2531
rect 1930 2528 1942 2531
rect 2210 2528 2262 2531
rect 2266 2528 2382 2531
rect 2682 2528 2742 2531
rect 2746 2528 2750 2531
rect 2802 2528 2990 2531
rect 3010 2528 3030 2531
rect 3098 2528 3102 2531
rect 3118 2528 3134 2531
rect 3154 2528 3198 2531
rect 3266 2528 3406 2531
rect 3482 2528 3486 2531
rect 3506 2528 3542 2531
rect 3598 2531 3601 2538
rect 3594 2528 3678 2531
rect 3682 2528 3750 2531
rect 3754 2528 3774 2531
rect 3778 2528 3854 2531
rect 3874 2528 3926 2531
rect 3978 2528 3982 2531
rect 3986 2528 4126 2531
rect 4186 2528 4278 2531
rect 4294 2531 4297 2538
rect 4294 2528 4326 2531
rect 4346 2528 4350 2531
rect 4466 2528 4486 2531
rect 4782 2531 4785 2538
rect 4570 2528 4785 2531
rect 4930 2528 5030 2531
rect 5034 2528 5046 2531
rect 1214 2522 1217 2528
rect 1630 2522 1633 2528
rect 2102 2522 2105 2528
rect 170 2518 222 2521
rect 226 2518 318 2521
rect 466 2518 486 2521
rect 850 2518 878 2521
rect 1026 2518 1094 2521
rect 1218 2518 1454 2521
rect 1466 2518 1590 2521
rect 1834 2518 2038 2521
rect 2126 2521 2129 2528
rect 3118 2522 3121 2528
rect 2126 2518 2134 2521
rect 2234 2518 2278 2521
rect 2282 2518 2382 2521
rect 2658 2518 2670 2521
rect 2674 2518 2806 2521
rect 2882 2518 2894 2521
rect 2938 2518 3030 2521
rect 3042 2518 3118 2521
rect 3170 2518 3254 2521
rect 3298 2518 3454 2521
rect 3474 2518 3614 2521
rect 3618 2518 3625 2521
rect 3634 2518 3822 2521
rect 3826 2518 4030 2521
rect 4042 2518 4158 2521
rect 4382 2521 4385 2528
rect 4314 2518 4385 2521
rect 4642 2518 4646 2521
rect 4694 2518 4750 2521
rect 4786 2518 4902 2521
rect 4906 2518 4934 2521
rect 4970 2518 5086 2521
rect 5090 2518 5158 2521
rect 5258 2518 5278 2521
rect 138 2508 398 2511
rect 546 2508 686 2511
rect 690 2508 790 2511
rect 962 2508 1078 2511
rect 1082 2508 1142 2511
rect 1146 2508 1462 2511
rect 1466 2508 1558 2511
rect 1562 2508 1678 2511
rect 1898 2508 1918 2511
rect 2098 2508 2230 2511
rect 2290 2508 2342 2511
rect 2354 2508 2510 2511
rect 2674 2508 2726 2511
rect 2738 2508 2782 2511
rect 2810 2508 2878 2511
rect 2922 2508 2942 2511
rect 2954 2508 3190 2511
rect 3202 2508 3238 2511
rect 3274 2508 3326 2511
rect 3370 2508 3614 2511
rect 3770 2508 3782 2511
rect 3818 2508 3830 2511
rect 3906 2508 3910 2511
rect 4694 2511 4697 2518
rect 4098 2508 4377 2511
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 862 2503 864 2507
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1886 2503 1888 2507
rect 154 2498 174 2501
rect 266 2498 422 2501
rect 442 2498 470 2501
rect 1154 2498 1174 2501
rect 1210 2498 1318 2501
rect 1322 2498 1486 2501
rect 1498 2498 1502 2501
rect 1530 2498 1598 2501
rect 2018 2498 2078 2501
rect 2098 2498 2158 2501
rect 2286 2501 2289 2508
rect 2888 2503 2890 2507
rect 2894 2503 2897 2507
rect 2902 2503 2904 2507
rect 3920 2503 3922 2507
rect 3926 2503 3929 2507
rect 3934 2503 3936 2507
rect 2178 2498 2289 2501
rect 2306 2498 2422 2501
rect 2626 2498 2630 2501
rect 2634 2498 2846 2501
rect 2930 2498 3038 2501
rect 3050 2498 3070 2501
rect 3226 2498 3230 2501
rect 3274 2498 3302 2501
rect 3306 2498 3342 2501
rect 3354 2498 3358 2501
rect 3450 2498 3646 2501
rect 3658 2498 3870 2501
rect 4066 2498 4078 2501
rect 4146 2498 4198 2501
rect 4234 2498 4326 2501
rect 4330 2498 4366 2501
rect 4374 2501 4377 2508
rect 4510 2508 4697 2511
rect 4706 2508 4926 2511
rect 4510 2502 4513 2508
rect 4936 2503 4938 2507
rect 4942 2503 4945 2507
rect 4950 2503 4952 2507
rect 5190 2502 5193 2508
rect 4374 2498 4510 2501
rect 4594 2498 4734 2501
rect 4738 2498 4838 2501
rect 4978 2498 5070 2501
rect 5098 2498 5118 2501
rect 1518 2492 1521 2498
rect 314 2488 350 2491
rect 354 2488 478 2491
rect 826 2488 1022 2491
rect 1994 2488 1998 2491
rect 2002 2488 2022 2491
rect 2058 2488 2062 2491
rect 2098 2488 2257 2491
rect 162 2478 182 2481
rect 186 2478 334 2481
rect 562 2478 590 2481
rect 606 2481 609 2488
rect 606 2478 742 2481
rect 1370 2478 1414 2481
rect 1646 2481 1649 2488
rect 2254 2482 2257 2488
rect 2602 2488 2694 2491
rect 2706 2488 2782 2491
rect 2794 2488 2798 2491
rect 2946 2488 3006 2491
rect 3018 2488 3022 2491
rect 3066 2488 3286 2491
rect 3290 2488 3718 2491
rect 3746 2488 4361 2491
rect 4378 2488 4710 2491
rect 4762 2488 4870 2491
rect 4890 2488 5006 2491
rect 5194 2488 5198 2491
rect 2374 2482 2377 2488
rect 2558 2482 2561 2488
rect 1646 2478 1902 2481
rect 1922 2478 2086 2481
rect 2106 2478 2118 2481
rect 2386 2478 2534 2481
rect 2666 2478 2726 2481
rect 2746 2478 2774 2481
rect 3062 2481 3065 2488
rect 4358 2482 4361 2488
rect 2882 2478 3065 2481
rect 3082 2478 3086 2481
rect 3194 2478 3230 2481
rect 3258 2478 3278 2481
rect 3282 2478 3294 2481
rect 3330 2478 3350 2481
rect 3490 2478 3553 2481
rect 3610 2478 3614 2481
rect 3634 2478 3705 2481
rect 98 2468 150 2471
rect 226 2468 310 2471
rect 498 2468 574 2471
rect 578 2468 646 2471
rect 706 2468 718 2471
rect 754 2468 822 2471
rect 826 2468 846 2471
rect 866 2468 918 2471
rect 950 2468 990 2471
rect 1026 2468 1030 2471
rect 1202 2468 1214 2471
rect 1242 2468 1302 2471
rect 1402 2468 1446 2471
rect 1474 2468 1494 2471
rect 1514 2468 1534 2471
rect 1618 2468 1622 2471
rect 1762 2468 1782 2471
rect 1786 2468 1814 2471
rect 1834 2468 1878 2471
rect 1890 2468 1990 2471
rect 2018 2468 2022 2471
rect 2034 2468 2358 2471
rect 2362 2468 2470 2471
rect 2482 2468 2577 2471
rect 122 2458 182 2461
rect 186 2458 278 2461
rect 282 2458 286 2461
rect 322 2458 518 2461
rect 522 2458 542 2461
rect 610 2458 614 2461
rect 674 2458 702 2461
rect 726 2461 729 2468
rect 726 2458 798 2461
rect 834 2458 878 2461
rect 890 2458 934 2461
rect 950 2461 953 2468
rect 950 2458 958 2461
rect 978 2458 982 2461
rect 1010 2458 1054 2461
rect 1062 2461 1065 2468
rect 1062 2458 1134 2461
rect 1202 2458 1214 2461
rect 1218 2458 1326 2461
rect 1410 2458 1526 2461
rect 1546 2458 1550 2461
rect 1578 2458 1582 2461
rect 1606 2461 1609 2468
rect 2574 2462 2577 2468
rect 2754 2468 2758 2471
rect 2786 2468 2801 2471
rect 2834 2468 2846 2471
rect 2882 2468 2958 2471
rect 2962 2468 2990 2471
rect 2994 2468 3038 2471
rect 3042 2468 3118 2471
rect 3170 2468 3185 2471
rect 3202 2468 3206 2471
rect 3274 2468 3286 2471
rect 3338 2468 3342 2471
rect 3374 2471 3377 2478
rect 3550 2472 3553 2478
rect 3702 2472 3705 2478
rect 3898 2478 4102 2481
rect 4130 2478 4142 2481
rect 4194 2478 4326 2481
rect 4466 2478 4494 2481
rect 4698 2478 4774 2481
rect 4794 2478 4934 2481
rect 5042 2478 5078 2481
rect 3362 2468 3377 2471
rect 3382 2468 3494 2471
rect 3514 2468 3518 2471
rect 3586 2468 3654 2471
rect 3658 2468 3686 2471
rect 3710 2471 3713 2478
rect 3710 2468 3726 2471
rect 3834 2468 3838 2471
rect 3882 2468 3934 2471
rect 3938 2468 4054 2471
rect 4114 2468 4126 2471
rect 4130 2468 4198 2471
rect 4218 2468 4246 2471
rect 4250 2468 4270 2471
rect 4282 2468 4294 2471
rect 4354 2468 4358 2471
rect 4382 2471 4385 2478
rect 4382 2468 4390 2471
rect 4418 2468 4422 2471
rect 4434 2468 4478 2471
rect 4514 2468 4518 2471
rect 4626 2468 4649 2471
rect 4658 2468 4678 2471
rect 4690 2468 4798 2471
rect 5154 2468 5209 2471
rect 2694 2462 2697 2468
rect 2710 2462 2713 2468
rect 2718 2462 2721 2468
rect 2798 2462 2801 2468
rect 1606 2458 1638 2461
rect 1794 2458 1798 2461
rect 1802 2458 1830 2461
rect 1842 2458 1846 2461
rect 1890 2458 1894 2461
rect 1938 2458 2057 2461
rect 2082 2458 2110 2461
rect 2114 2458 2118 2461
rect 2138 2458 2158 2461
rect 2226 2458 2238 2461
rect 2338 2458 2350 2461
rect 2414 2458 2446 2461
rect 2458 2458 2462 2461
rect 2466 2458 2510 2461
rect 2730 2458 2750 2461
rect 2862 2461 2865 2468
rect 3182 2462 3185 2468
rect 2862 2458 2937 2461
rect 1934 2452 1937 2458
rect 2054 2452 2057 2458
rect 2126 2452 2129 2458
rect 2286 2452 2289 2458
rect 2414 2452 2417 2458
rect 2542 2452 2545 2458
rect 2846 2452 2849 2458
rect 2934 2452 2937 2458
rect 2942 2458 2958 2461
rect 2970 2458 2974 2461
rect 2982 2458 3014 2461
rect 3066 2458 3078 2461
rect 3082 2458 3166 2461
rect 3190 2458 3302 2461
rect 3330 2458 3334 2461
rect 3382 2461 3385 2468
rect 3542 2462 3545 2468
rect 3354 2458 3385 2461
rect 3402 2458 3526 2461
rect 3578 2458 3622 2461
rect 3890 2458 3894 2461
rect 4010 2458 4030 2461
rect 4034 2458 4078 2461
rect 4090 2458 4094 2461
rect 4114 2458 4190 2461
rect 4290 2458 4294 2461
rect 4322 2458 4374 2461
rect 4438 2458 4446 2461
rect 4450 2458 4470 2461
rect 4634 2458 4638 2461
rect 4646 2461 4649 2468
rect 5206 2462 5209 2468
rect 4646 2458 4694 2461
rect 4770 2458 4942 2461
rect 2942 2452 2945 2458
rect 2982 2452 2985 2458
rect 42 2448 113 2451
rect 122 2448 158 2451
rect 418 2448 446 2451
rect 514 2448 526 2451
rect 530 2448 630 2451
rect 634 2448 646 2451
rect 650 2448 878 2451
rect 930 2448 1070 2451
rect 1242 2448 1257 2451
rect 110 2442 113 2448
rect 894 2442 897 2448
rect 1254 2442 1257 2448
rect 1270 2448 1358 2451
rect 1458 2448 1510 2451
rect 1690 2448 1806 2451
rect 1826 2448 1841 2451
rect 1922 2448 1926 2451
rect 2090 2448 2102 2451
rect 2186 2448 2246 2451
rect 2458 2448 2462 2451
rect 2626 2448 2838 2451
rect 3038 2448 3126 2451
rect 3190 2451 3193 2458
rect 4254 2452 4257 2458
rect 3154 2448 3193 2451
rect 3250 2448 3254 2451
rect 3314 2448 3502 2451
rect 3506 2448 3646 2451
rect 3738 2448 3750 2451
rect 3786 2448 3918 2451
rect 3986 2448 4006 2451
rect 4050 2448 4054 2451
rect 4290 2448 4302 2451
rect 4314 2448 4406 2451
rect 4410 2448 4414 2451
rect 4466 2448 4542 2451
rect 4622 2448 4630 2451
rect 4634 2448 4734 2451
rect 4746 2448 4750 2451
rect 4786 2448 4790 2451
rect 4802 2448 4806 2451
rect 4930 2448 4958 2451
rect 4962 2448 5022 2451
rect 5082 2448 5126 2451
rect 1270 2442 1273 2448
rect 1646 2442 1649 2448
rect 1838 2442 1841 2448
rect 1966 2442 1969 2448
rect 2142 2442 2145 2448
rect 2534 2442 2537 2448
rect 146 2438 150 2441
rect 394 2438 478 2441
rect 658 2438 710 2441
rect 994 2438 1014 2441
rect 1050 2438 1054 2441
rect 1058 2438 1065 2441
rect 1074 2438 1158 2441
rect 1186 2438 1246 2441
rect 1306 2438 1454 2441
rect 1458 2438 1470 2441
rect 1690 2438 1710 2441
rect 2090 2438 2134 2441
rect 2242 2438 2270 2441
rect 2274 2438 2326 2441
rect 2386 2438 2430 2441
rect 3038 2441 3041 2448
rect 2542 2438 3041 2441
rect 3058 2438 3166 2441
rect 3182 2438 3318 2441
rect 3322 2438 3366 2441
rect 3370 2438 3510 2441
rect 3514 2438 3558 2441
rect 3562 2438 3598 2441
rect 3602 2438 3734 2441
rect 3738 2438 3886 2441
rect 3970 2438 4134 2441
rect 4274 2438 4358 2441
rect 4378 2438 4558 2441
rect 4642 2438 4790 2441
rect 4794 2438 4918 2441
rect 4970 2438 5054 2441
rect 5058 2438 5150 2441
rect 250 2428 454 2431
rect 714 2428 758 2431
rect 774 2431 777 2438
rect 774 2428 902 2431
rect 930 2428 934 2431
rect 950 2431 953 2438
rect 950 2428 1230 2431
rect 1346 2428 1438 2431
rect 1458 2428 2358 2431
rect 2374 2431 2377 2438
rect 2542 2431 2545 2438
rect 2374 2428 2545 2431
rect 2550 2428 2558 2431
rect 2562 2428 2686 2431
rect 2734 2428 2742 2431
rect 2746 2428 2814 2431
rect 2830 2428 2838 2431
rect 2842 2428 2878 2431
rect 2898 2428 2902 2431
rect 2962 2428 2990 2431
rect 3182 2431 3185 2438
rect 3154 2428 3185 2431
rect 3194 2428 3230 2431
rect 3250 2428 3582 2431
rect 3650 2428 3662 2431
rect 3698 2428 3742 2431
rect 3866 2428 4062 2431
rect 4066 2428 4073 2431
rect 4098 2428 4246 2431
rect 4266 2428 4294 2431
rect 4458 2428 4710 2431
rect 4714 2428 4894 2431
rect 4898 2428 4910 2431
rect 3062 2422 3065 2428
rect 234 2418 462 2421
rect 466 2418 702 2421
rect 706 2418 1558 2421
rect 1738 2418 1750 2421
rect 1866 2418 1942 2421
rect 2058 2418 2158 2421
rect 2166 2418 2174 2421
rect 2178 2418 3054 2421
rect 3142 2421 3145 2428
rect 3142 2418 3222 2421
rect 3234 2418 3446 2421
rect 3522 2418 3726 2421
rect 3738 2418 4046 2421
rect 4074 2418 4102 2421
rect 4122 2418 4382 2421
rect 4386 2418 4398 2421
rect 4434 2418 4478 2421
rect 4482 2418 5294 2421
rect 282 2408 318 2411
rect 450 2408 670 2411
rect 762 2408 1046 2411
rect 1066 2408 1270 2411
rect 1402 2408 1406 2411
rect 1434 2408 1470 2411
rect 1506 2408 1550 2411
rect 1778 2408 1822 2411
rect 1858 2408 2086 2411
rect 2098 2408 2118 2411
rect 2218 2408 2326 2411
rect 2442 2408 2446 2411
rect 2554 2408 2558 2411
rect 2638 2408 2662 2411
rect 2754 2408 2766 2411
rect 2794 2408 2798 2411
rect 2866 2408 2870 2411
rect 2938 2408 2950 2411
rect 2986 2408 3254 2411
rect 3442 2408 3574 2411
rect 3586 2408 3606 2411
rect 3690 2408 3894 2411
rect 3906 2408 4262 2411
rect 4498 2408 4542 2411
rect 5290 2408 5294 2411
rect 5334 2411 5338 2412
rect 5298 2408 5338 2411
rect 278 2402 281 2408
rect 328 2403 330 2407
rect 334 2403 337 2407
rect 342 2403 344 2407
rect 1352 2403 1354 2407
rect 1358 2403 1361 2407
rect 1366 2403 1368 2407
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2398 2403 2400 2407
rect 578 2398 838 2401
rect 882 2398 1054 2401
rect 1386 2398 1390 2401
rect 1402 2398 1486 2401
rect 1522 2398 1534 2401
rect 1538 2398 1710 2401
rect 1770 2398 1774 2401
rect 1834 2398 1966 2401
rect 1986 2398 2022 2401
rect 2122 2398 2158 2401
rect 2170 2398 2342 2401
rect 2638 2401 2641 2408
rect 3400 2403 3402 2407
rect 3406 2403 3409 2407
rect 3414 2403 3416 2407
rect 4424 2403 4426 2407
rect 4430 2403 4433 2407
rect 4438 2403 4440 2407
rect 2538 2398 2641 2401
rect 2666 2398 2686 2401
rect 2722 2398 2726 2401
rect 2794 2398 3094 2401
rect 3138 2398 3142 2401
rect 3202 2398 3374 2401
rect 3442 2398 3478 2401
rect 3530 2398 3662 2401
rect 3666 2398 3734 2401
rect 3746 2398 3894 2401
rect 3914 2398 4166 2401
rect 4170 2398 4310 2401
rect 4402 2398 4406 2401
rect 4690 2398 5337 2401
rect 594 2388 630 2391
rect 634 2388 734 2391
rect 898 2388 966 2391
rect 1234 2388 1326 2391
rect 1386 2388 1630 2391
rect 1642 2388 2198 2391
rect 2250 2388 2369 2391
rect 2378 2388 2446 2391
rect 2482 2388 2566 2391
rect 2578 2388 2638 2391
rect 2650 2388 3070 2391
rect 3074 2388 3342 2391
rect 3362 2388 3422 2391
rect 3478 2391 3481 2398
rect 5334 2392 5337 2398
rect 3478 2388 3694 2391
rect 3746 2388 3769 2391
rect 3826 2388 4057 2391
rect 4082 2388 4150 2391
rect 4162 2388 4169 2391
rect 378 2378 470 2381
rect 474 2378 694 2381
rect 698 2378 726 2381
rect 730 2378 846 2381
rect 850 2378 998 2381
rect 1002 2378 1022 2381
rect 1026 2378 1318 2381
rect 1322 2378 1390 2381
rect 1394 2378 2134 2381
rect 2162 2378 2182 2381
rect 2314 2378 2358 2381
rect 2366 2381 2369 2388
rect 3766 2382 3769 2388
rect 4054 2382 4057 2388
rect 4166 2382 4169 2388
rect 4346 2388 4502 2391
rect 4506 2388 4534 2391
rect 4618 2388 5030 2391
rect 5034 2388 5078 2391
rect 5106 2388 5126 2391
rect 5138 2388 5262 2391
rect 5334 2388 5338 2392
rect 2366 2378 2622 2381
rect 2626 2378 2750 2381
rect 2754 2378 3030 2381
rect 3034 2378 3166 2381
rect 3314 2378 3318 2381
rect 3370 2378 3414 2381
rect 3478 2378 3590 2381
rect 3738 2378 3758 2381
rect 3794 2378 3806 2381
rect 3922 2378 3982 2381
rect 4294 2381 4297 2388
rect 4258 2378 4297 2381
rect 4354 2378 4574 2381
rect 4690 2378 4710 2381
rect 4786 2378 4886 2381
rect 4898 2378 5062 2381
rect 5162 2378 5302 2381
rect 506 2368 526 2371
rect 834 2368 934 2371
rect 938 2368 945 2371
rect 1130 2368 1182 2371
rect 1186 2368 1558 2371
rect 1566 2368 1614 2371
rect 1618 2368 1846 2371
rect 1882 2368 1886 2371
rect 1930 2368 2166 2371
rect 2226 2368 2230 2371
rect 2258 2368 2270 2371
rect 2282 2368 2329 2371
rect 2418 2368 2494 2371
rect 2618 2368 2734 2371
rect 2738 2368 2790 2371
rect 2794 2368 2846 2371
rect 2850 2368 2918 2371
rect 2922 2368 2974 2371
rect 3034 2368 3134 2371
rect 3478 2371 3481 2378
rect 3258 2368 3481 2371
rect 3490 2368 3494 2371
rect 3506 2368 3510 2371
rect 3530 2368 3542 2371
rect 3602 2368 3614 2371
rect 3650 2368 3790 2371
rect 3866 2368 3878 2371
rect 3970 2368 4022 2371
rect 4190 2368 4206 2371
rect 4242 2368 4406 2371
rect 4562 2368 4654 2371
rect 5058 2368 5270 2371
rect 5334 2371 5338 2372
rect 5290 2368 5338 2371
rect 322 2358 414 2361
rect 542 2361 545 2368
rect 542 2358 574 2361
rect 678 2361 681 2368
rect 666 2358 681 2361
rect 906 2358 1038 2361
rect 1066 2358 1126 2361
rect 1130 2358 1137 2361
rect 1194 2358 1206 2361
rect 1314 2358 1526 2361
rect 1566 2361 1569 2368
rect 1546 2358 1569 2361
rect 1602 2358 1662 2361
rect 1730 2358 1750 2361
rect 1754 2358 1774 2361
rect 1786 2358 1798 2361
rect 1810 2358 1958 2361
rect 1970 2358 2022 2361
rect 2082 2358 2094 2361
rect 2194 2358 2206 2361
rect 2226 2358 2238 2361
rect 2266 2358 2270 2361
rect 2278 2358 2294 2361
rect 2326 2361 2329 2368
rect 2502 2362 2505 2368
rect 4190 2362 4193 2368
rect 2326 2358 2422 2361
rect 2522 2358 2606 2361
rect 2626 2358 2630 2361
rect 2650 2358 2654 2361
rect 2714 2358 2774 2361
rect 2778 2358 2830 2361
rect 2938 2358 2998 2361
rect 3010 2358 3014 2361
rect 3090 2358 3110 2361
rect 3218 2358 3249 2361
rect 3298 2358 3318 2361
rect 3322 2358 3350 2361
rect 3370 2358 3398 2361
rect 3426 2358 3574 2361
rect 3578 2358 3614 2361
rect 3634 2358 3814 2361
rect 3882 2358 3894 2361
rect 3898 2358 3958 2361
rect 3994 2358 4014 2361
rect 4042 2358 4070 2361
rect 4106 2358 4126 2361
rect 4194 2358 4310 2361
rect 4370 2358 4486 2361
rect 4510 2361 4513 2368
rect 4510 2358 4582 2361
rect 4634 2358 4641 2361
rect 4738 2358 4790 2361
rect 4814 2361 4817 2368
rect 4794 2358 4817 2361
rect 5018 2358 5110 2361
rect 5250 2358 5278 2361
rect 158 2351 161 2358
rect 122 2348 161 2351
rect 222 2351 225 2358
rect 210 2348 225 2351
rect 462 2351 465 2358
rect 442 2348 465 2351
rect 498 2348 502 2351
rect 530 2348 534 2351
rect 546 2348 577 2351
rect 618 2348 646 2351
rect 658 2348 662 2351
rect 718 2351 721 2358
rect 706 2348 721 2351
rect 746 2348 750 2351
rect 930 2348 934 2351
rect 1026 2348 1126 2351
rect 1130 2348 1182 2351
rect 1254 2351 1257 2358
rect 1670 2352 1673 2358
rect 2070 2352 2073 2358
rect 1210 2348 1257 2351
rect 1370 2348 1374 2351
rect 1450 2348 1462 2351
rect 1466 2348 1478 2351
rect 1530 2348 1630 2351
rect 1682 2348 1710 2351
rect 1714 2348 1742 2351
rect 1762 2348 1782 2351
rect 1842 2348 1846 2351
rect 1890 2348 1926 2351
rect 1938 2348 2046 2351
rect 2082 2348 2134 2351
rect 2238 2348 2246 2351
rect 2278 2351 2281 2358
rect 2430 2352 2433 2358
rect 3118 2352 3121 2358
rect 2250 2348 2281 2351
rect 2402 2348 2406 2351
rect 2546 2348 2558 2351
rect 2650 2348 2822 2351
rect 2842 2348 2854 2351
rect 2858 2348 2862 2351
rect 2886 2348 2894 2351
rect 2898 2348 3046 2351
rect 3058 2348 3062 2351
rect 3098 2348 3102 2351
rect 3130 2348 3166 2351
rect 3170 2348 3190 2351
rect 3202 2348 3238 2351
rect 3246 2351 3249 2358
rect 3246 2348 3254 2351
rect 3330 2348 3334 2351
rect 3354 2348 3382 2351
rect 3386 2348 3430 2351
rect 3442 2348 3446 2351
rect 3466 2348 3518 2351
rect 3522 2348 3550 2351
rect 3642 2348 3646 2351
rect 3682 2348 3686 2351
rect 3698 2348 3750 2351
rect 3838 2351 3841 2358
rect 4638 2352 4641 2358
rect 4958 2352 4961 2358
rect 3838 2348 3870 2351
rect 3962 2348 3974 2351
rect 3986 2348 3990 2351
rect 4002 2348 4038 2351
rect 4050 2348 4118 2351
rect 4154 2348 4174 2351
rect 4290 2348 4310 2351
rect 4354 2348 4366 2351
rect 4490 2348 4526 2351
rect 4530 2348 4614 2351
rect 4666 2348 4702 2351
rect 4706 2348 4798 2351
rect 4970 2348 4982 2351
rect 5162 2348 5174 2351
rect 5334 2351 5338 2352
rect 5298 2348 5338 2351
rect 574 2342 577 2348
rect 1430 2342 1433 2348
rect 1502 2342 1505 2348
rect 130 2338 134 2341
rect 146 2338 302 2341
rect 458 2338 462 2341
rect 522 2338 526 2341
rect 658 2338 766 2341
rect 934 2338 942 2341
rect 1130 2338 1134 2341
rect 1146 2338 1233 2341
rect 1346 2338 1430 2341
rect 1450 2338 1494 2341
rect 1586 2338 1622 2341
rect 1634 2338 1638 2341
rect 1698 2338 1702 2341
rect 1754 2338 1766 2341
rect 1802 2338 1830 2341
rect 1898 2338 2174 2341
rect 2242 2338 2246 2341
rect 2282 2338 2294 2341
rect 2298 2338 2374 2341
rect 2514 2338 2638 2341
rect 2690 2338 2766 2341
rect 2850 2338 2854 2341
rect 2890 2338 2894 2341
rect 2962 2338 2966 2341
rect 2978 2338 2982 2341
rect 2986 2338 2990 2341
rect 3002 2338 3006 2341
rect 3018 2338 3022 2341
rect 3162 2338 3334 2341
rect 3346 2338 3526 2341
rect 3666 2338 3950 2341
rect 3986 2338 4030 2341
rect 4106 2338 4110 2341
rect 4486 2338 4606 2341
rect 4666 2338 4678 2341
rect 4714 2338 4726 2341
rect 4810 2338 4966 2341
rect 4970 2338 4998 2341
rect 5178 2338 5217 2341
rect 5242 2338 5246 2341
rect 42 2328 174 2331
rect 242 2328 350 2331
rect 482 2328 654 2331
rect 782 2331 785 2338
rect 782 2328 814 2331
rect 910 2331 913 2338
rect 818 2328 913 2331
rect 934 2332 937 2338
rect 1230 2332 1233 2338
rect 2670 2332 2673 2338
rect 986 2328 1110 2331
rect 1114 2328 1166 2331
rect 1386 2328 1462 2331
rect 1570 2328 1606 2331
rect 1618 2328 1758 2331
rect 1826 2328 1974 2331
rect 2042 2328 2110 2331
rect 2114 2328 2126 2331
rect 2286 2328 2318 2331
rect 2338 2328 2454 2331
rect 2490 2328 2518 2331
rect 2546 2328 2574 2331
rect 2594 2328 2662 2331
rect 2706 2328 2806 2331
rect 2814 2331 2817 2338
rect 2814 2328 3134 2331
rect 3170 2328 3198 2331
rect 3218 2328 3222 2331
rect 3266 2328 3294 2331
rect 3330 2328 3390 2331
rect 3402 2328 3758 2331
rect 3762 2328 3814 2331
rect 3890 2328 3926 2331
rect 4074 2328 4198 2331
rect 4202 2328 4222 2331
rect 4486 2331 4489 2338
rect 5214 2332 5217 2338
rect 4322 2328 4489 2331
rect 4682 2328 4718 2331
rect 4818 2328 4902 2331
rect 4994 2328 5046 2331
rect 186 2318 278 2321
rect 702 2321 705 2328
rect 702 2318 838 2321
rect 858 2318 886 2321
rect 890 2318 902 2321
rect 910 2321 913 2328
rect 910 2318 982 2321
rect 1018 2318 1518 2321
rect 1534 2321 1537 2328
rect 2286 2322 2289 2328
rect 4286 2322 4289 2328
rect 1534 2318 1558 2321
rect 1602 2318 1606 2321
rect 1618 2318 1678 2321
rect 1690 2318 1694 2321
rect 1754 2318 1758 2321
rect 1906 2318 1934 2321
rect 1978 2318 2038 2321
rect 2066 2318 2070 2321
rect 2530 2318 2566 2321
rect 2570 2318 2614 2321
rect 2642 2318 3006 2321
rect 3026 2318 3038 2321
rect 3042 2318 3126 2321
rect 3146 2318 3198 2321
rect 3314 2318 3342 2321
rect 3418 2318 3478 2321
rect 3490 2318 3494 2321
rect 3518 2318 3526 2321
rect 3618 2318 3622 2321
rect 3754 2318 3830 2321
rect 3850 2318 4022 2321
rect 4026 2318 4078 2321
rect 4194 2318 4270 2321
rect 4306 2318 4398 2321
rect 4402 2318 4550 2321
rect 4670 2321 4673 2328
rect 4670 2318 4686 2321
rect 4694 2318 4702 2321
rect 4706 2318 4758 2321
rect 4770 2318 4782 2321
rect 4786 2318 4838 2321
rect 4930 2318 5030 2321
rect 2190 2312 2193 2318
rect 2318 2312 2321 2318
rect 3374 2312 3377 2318
rect 3518 2312 3521 2318
rect 274 2308 294 2311
rect 426 2308 470 2311
rect 474 2308 742 2311
rect 978 2308 1398 2311
rect 1506 2308 1614 2311
rect 1666 2308 1862 2311
rect 1898 2308 1974 2311
rect 1994 2308 2038 2311
rect 2042 2308 2150 2311
rect 2202 2308 2230 2311
rect 2378 2308 2494 2311
rect 2498 2308 2534 2311
rect 2610 2308 2622 2311
rect 2666 2308 2822 2311
rect 2922 2308 2926 2311
rect 3018 2308 3062 2311
rect 3194 2308 3286 2311
rect 3290 2308 3350 2311
rect 3410 2308 3430 2311
rect 3450 2308 3502 2311
rect 3586 2308 3638 2311
rect 3778 2308 3790 2311
rect 3794 2308 3910 2311
rect 3986 2308 3990 2311
rect 4002 2308 4022 2311
rect 4778 2308 4846 2311
rect 5130 2308 5214 2311
rect 5226 2308 5254 2311
rect 5258 2308 5270 2311
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 862 2303 864 2307
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1886 2303 1888 2307
rect 2888 2303 2890 2307
rect 2894 2303 2897 2307
rect 2902 2303 2904 2307
rect 2950 2302 2953 2308
rect 3920 2303 3922 2307
rect 3926 2303 3929 2307
rect 3934 2303 3936 2307
rect 4936 2303 4938 2307
rect 4942 2303 4945 2307
rect 4950 2303 4952 2307
rect 290 2298 726 2301
rect 994 2298 1022 2301
rect 1026 2298 1158 2301
rect 1162 2298 1246 2301
rect 1250 2298 1406 2301
rect 1442 2298 1454 2301
rect 1458 2298 1577 2301
rect 1738 2298 1790 2301
rect 1994 2298 2118 2301
rect 2178 2298 2270 2301
rect 2282 2298 2334 2301
rect 2362 2298 2638 2301
rect 2650 2298 2718 2301
rect 2730 2298 2774 2301
rect 2810 2298 2838 2301
rect 3130 2298 3222 2301
rect 3234 2298 3286 2301
rect 3290 2298 3398 2301
rect 3410 2298 3670 2301
rect 3818 2298 3854 2301
rect 3890 2298 3910 2301
rect 3978 2298 3982 2301
rect 4266 2298 4342 2301
rect 4490 2298 4766 2301
rect 4842 2298 4918 2301
rect 5018 2298 5086 2301
rect 154 2288 166 2291
rect 170 2288 206 2291
rect 210 2288 390 2291
rect 410 2288 446 2291
rect 466 2288 550 2291
rect 554 2288 654 2291
rect 714 2288 974 2291
rect 1202 2288 1294 2291
rect 1470 2288 1478 2291
rect 1482 2288 1566 2291
rect 1574 2291 1577 2298
rect 1574 2288 1910 2291
rect 1962 2288 1966 2291
rect 1994 2288 2006 2291
rect 2162 2288 2510 2291
rect 2530 2288 2574 2291
rect 2622 2288 2630 2291
rect 2634 2288 2662 2291
rect 2674 2288 2678 2291
rect 2714 2288 2862 2291
rect 2906 2288 2942 2291
rect 3050 2288 3182 2291
rect 3210 2288 3270 2291
rect 3282 2288 3334 2291
rect 3386 2288 3462 2291
rect 3474 2288 3478 2291
rect 3486 2288 3494 2291
rect 3498 2288 3558 2291
rect 3570 2288 3601 2291
rect 3618 2288 3694 2291
rect 3738 2288 3774 2291
rect 3866 2288 4070 2291
rect 4082 2288 4230 2291
rect 4250 2288 4334 2291
rect 4338 2288 4438 2291
rect 4762 2288 4814 2291
rect 4826 2288 4830 2291
rect 4834 2288 4854 2291
rect 5154 2288 5158 2291
rect 5258 2288 5262 2291
rect 42 2278 126 2281
rect 150 2278 262 2281
rect 290 2278 302 2281
rect 370 2278 758 2281
rect 1106 2278 1198 2281
rect 1266 2278 1270 2281
rect 1282 2278 1342 2281
rect 1370 2278 1374 2281
rect 1394 2278 1406 2281
rect 1410 2278 1414 2281
rect 1534 2278 1630 2281
rect 1658 2278 1774 2281
rect 2054 2281 2057 2288
rect 3598 2282 3601 2288
rect 1914 2278 2057 2281
rect 2066 2278 2118 2281
rect 2274 2278 2742 2281
rect 2794 2278 3526 2281
rect 3530 2278 3534 2281
rect 3682 2278 3750 2281
rect 3786 2278 3998 2281
rect 4234 2278 4238 2281
rect 4474 2278 4502 2281
rect 4546 2278 4558 2281
rect 4686 2281 4689 2288
rect 4686 2278 4750 2281
rect 4766 2278 4982 2281
rect 5022 2281 5025 2288
rect 4986 2278 5025 2281
rect 5106 2278 5174 2281
rect 150 2272 153 2278
rect 122 2268 150 2271
rect 178 2268 214 2271
rect 290 2268 294 2271
rect 402 2268 430 2271
rect 434 2268 446 2271
rect 602 2268 678 2271
rect 798 2271 801 2278
rect 1206 2272 1209 2278
rect 1534 2272 1537 2278
rect 3590 2272 3593 2278
rect 4134 2272 4137 2278
rect 786 2268 801 2271
rect 810 2268 822 2271
rect 826 2268 918 2271
rect 974 2268 990 2271
rect 1002 2268 1006 2271
rect 1090 2268 1137 2271
rect 1218 2268 1286 2271
rect 1290 2268 1518 2271
rect 1554 2268 1558 2271
rect 1562 2268 1678 2271
rect 1682 2268 1694 2271
rect 1730 2268 1862 2271
rect 1962 2268 1998 2271
rect 2010 2268 2046 2271
rect 2074 2268 2158 2271
rect 2226 2268 2246 2271
rect 2258 2268 2278 2271
rect 2338 2268 2430 2271
rect 2434 2268 2446 2271
rect 2482 2268 2486 2271
rect 2570 2268 2574 2271
rect 2650 2268 2686 2271
rect 2722 2268 2846 2271
rect 2858 2268 2886 2271
rect 2970 2268 3014 2271
rect 3018 2268 3110 2271
rect 3114 2268 3126 2271
rect 3138 2268 3158 2271
rect 3210 2268 3214 2271
rect 3218 2268 3246 2271
rect 3258 2268 3262 2271
rect 3314 2268 3318 2271
rect 3370 2270 3425 2271
rect 3370 2268 3422 2270
rect 718 2262 721 2268
rect 138 2258 190 2261
rect 218 2258 222 2261
rect 234 2258 246 2261
rect 282 2258 294 2261
rect 306 2258 358 2261
rect 426 2258 526 2261
rect 674 2258 702 2261
rect 762 2258 766 2261
rect 818 2259 894 2261
rect 974 2262 977 2268
rect 818 2258 897 2259
rect 1046 2261 1049 2268
rect 994 2258 1049 2261
rect 1066 2258 1086 2261
rect 1134 2261 1137 2268
rect 1134 2259 1142 2261
rect 1134 2258 1145 2259
rect 1234 2258 1246 2261
rect 1266 2258 1278 2261
rect 1290 2258 1430 2261
rect 1442 2258 1462 2261
rect 1482 2258 1486 2261
rect 1530 2258 1742 2261
rect 1762 2258 1894 2261
rect 1938 2258 1942 2261
rect 1954 2258 1974 2261
rect 2054 2261 2057 2268
rect 2302 2262 2305 2268
rect 2462 2262 2465 2268
rect 3442 2268 3446 2271
rect 3474 2268 3478 2271
rect 3490 2268 3494 2271
rect 3506 2268 3510 2271
rect 3522 2268 3526 2271
rect 3578 2268 3582 2271
rect 3626 2268 3630 2271
rect 3722 2268 3726 2271
rect 3834 2268 3878 2271
rect 3898 2268 3918 2271
rect 3946 2268 4078 2271
rect 4154 2268 4310 2271
rect 4318 2271 4321 2278
rect 4766 2272 4769 2278
rect 4318 2268 4358 2271
rect 4466 2268 4478 2271
rect 4554 2268 4718 2271
rect 4722 2268 4742 2271
rect 4810 2268 4838 2271
rect 4914 2268 5046 2271
rect 5146 2268 5150 2271
rect 5202 2268 5302 2271
rect 2026 2258 2057 2261
rect 2138 2258 2198 2261
rect 2378 2258 2446 2261
rect 2482 2258 2566 2261
rect 2578 2258 2590 2261
rect 2594 2258 2662 2261
rect 2666 2258 2670 2261
rect 2698 2258 2710 2261
rect 2714 2258 2726 2261
rect 2738 2258 2769 2261
rect 322 2248 326 2251
rect 438 2248 446 2251
rect 450 2248 494 2251
rect 690 2248 790 2251
rect 978 2248 1118 2251
rect 1306 2248 1318 2251
rect 1346 2248 1422 2251
rect 1426 2248 1758 2251
rect 1762 2248 2070 2251
rect 2146 2248 2150 2251
rect 2310 2251 2313 2258
rect 2766 2252 2769 2258
rect 2818 2258 2822 2261
rect 2882 2258 2934 2261
rect 2954 2258 2990 2261
rect 3002 2258 3662 2261
rect 3778 2258 3782 2261
rect 3818 2258 3982 2261
rect 4026 2258 4030 2261
rect 4090 2258 4166 2261
rect 4194 2258 4254 2261
rect 4282 2258 4334 2261
rect 4410 2258 4462 2261
rect 4538 2258 4542 2261
rect 4578 2258 4582 2261
rect 4594 2258 4734 2261
rect 4798 2261 4801 2268
rect 4798 2258 4806 2261
rect 4850 2258 5102 2261
rect 5106 2258 5150 2261
rect 5274 2258 5302 2261
rect 2782 2252 2785 2258
rect 4038 2252 4041 2258
rect 2310 2248 2342 2251
rect 2354 2248 2406 2251
rect 2410 2248 2417 2251
rect 2426 2248 2550 2251
rect 2562 2248 2630 2251
rect 2690 2248 2694 2251
rect 2722 2248 2726 2251
rect 2818 2248 2910 2251
rect 2994 2248 3022 2251
rect 3026 2248 3270 2251
rect 3274 2248 3374 2251
rect 3394 2248 3550 2251
rect 3562 2248 3566 2251
rect 3618 2248 3838 2251
rect 3954 2248 3990 2251
rect 4002 2248 4022 2251
rect 4310 2248 4318 2251
rect 4322 2248 4350 2251
rect 4458 2248 4526 2251
rect 4554 2248 4566 2251
rect 4570 2248 4606 2251
rect 4618 2248 4678 2251
rect 4734 2251 4737 2258
rect 4734 2248 5006 2251
rect 5010 2248 5070 2251
rect 5082 2248 5150 2251
rect 5334 2251 5338 2252
rect 5306 2248 5338 2251
rect 842 2238 958 2241
rect 962 2238 1286 2241
rect 1346 2238 1558 2241
rect 1562 2238 1678 2241
rect 2026 2238 2102 2241
rect 2250 2238 2366 2241
rect 2386 2238 2422 2241
rect 2458 2238 2510 2241
rect 2530 2238 2534 2241
rect 2538 2238 3326 2241
rect 3330 2238 3358 2241
rect 3382 2241 3385 2248
rect 3382 2238 3550 2241
rect 3554 2238 3638 2241
rect 3642 2238 3710 2241
rect 3850 2238 4006 2241
rect 4018 2238 4054 2241
rect 4134 2241 4137 2248
rect 4134 2238 4174 2241
rect 4290 2238 4398 2241
rect 4418 2238 4526 2241
rect 4882 2238 5086 2241
rect 5090 2238 5158 2241
rect 250 2228 382 2231
rect 750 2228 870 2231
rect 970 2228 2318 2231
rect 2362 2228 2414 2231
rect 2506 2228 2638 2231
rect 2698 2228 2718 2231
rect 2746 2228 2750 2231
rect 2778 2228 2830 2231
rect 2834 2228 4358 2231
rect 4442 2228 4734 2231
rect 4738 2228 4758 2231
rect 4930 2228 5238 2231
rect 750 2222 753 2228
rect 530 2218 542 2221
rect 546 2218 574 2221
rect 794 2218 1022 2221
rect 1042 2218 1430 2221
rect 1482 2218 1486 2221
rect 1498 2218 1542 2221
rect 1546 2218 1566 2221
rect 1678 2218 1686 2221
rect 1690 2218 1710 2221
rect 1754 2218 2006 2221
rect 2026 2218 2214 2221
rect 2218 2218 2374 2221
rect 2378 2218 2878 2221
rect 3006 2218 3014 2221
rect 3018 2218 3030 2221
rect 3090 2218 3126 2221
rect 3174 2218 3182 2221
rect 3186 2218 3262 2221
rect 3274 2218 3462 2221
rect 3490 2218 3574 2221
rect 3586 2218 3646 2221
rect 3658 2218 4086 2221
rect 4362 2218 4518 2221
rect 4522 2218 4590 2221
rect 4698 2218 4710 2221
rect 4714 2218 4854 2221
rect 4858 2218 4966 2221
rect 5074 2218 5142 2221
rect 5186 2218 5198 2221
rect 5250 2218 5270 2221
rect 3470 2212 3473 2218
rect 618 2208 974 2211
rect 986 2208 1334 2211
rect 1378 2208 1502 2211
rect 1650 2208 1678 2211
rect 1730 2208 1990 2211
rect 1994 2208 2286 2211
rect 2306 2208 2358 2211
rect 2410 2208 2494 2211
rect 2530 2208 2734 2211
rect 2762 2208 2870 2211
rect 2890 2208 2950 2211
rect 2954 2208 3046 2211
rect 3050 2208 3206 2211
rect 3218 2208 3302 2211
rect 3530 2208 3990 2211
rect 4002 2208 4198 2211
rect 4202 2208 4262 2211
rect 4450 2208 4849 2211
rect 4858 2208 4886 2211
rect 5082 2208 5262 2211
rect 328 2203 330 2207
rect 334 2203 337 2207
rect 342 2203 344 2207
rect 1352 2203 1354 2207
rect 1358 2203 1361 2207
rect 1366 2203 1368 2207
rect 2374 2202 2377 2208
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2398 2203 2400 2207
rect 3400 2203 3402 2207
rect 3406 2203 3409 2207
rect 3414 2203 3416 2207
rect 4424 2203 4426 2207
rect 4430 2203 4433 2207
rect 4438 2203 4440 2207
rect 770 2198 1278 2201
rect 1426 2198 1734 2201
rect 1834 2198 1894 2201
rect 1930 2198 2086 2201
rect 2210 2198 2238 2201
rect 2282 2198 2358 2201
rect 2538 2198 2542 2201
rect 2746 2198 2998 2201
rect 3442 2198 3662 2201
rect 3722 2198 3862 2201
rect 3866 2198 3886 2201
rect 3970 2198 3974 2201
rect 4018 2198 4102 2201
rect 4106 2198 4414 2201
rect 4846 2201 4849 2208
rect 4846 2198 4958 2201
rect 5034 2198 5198 2201
rect 5266 2198 5278 2201
rect 750 2192 753 2198
rect 362 2188 734 2191
rect 754 2188 806 2191
rect 946 2188 1014 2191
rect 1206 2188 1238 2191
rect 1658 2188 1694 2191
rect 1698 2188 1742 2191
rect 1946 2188 1950 2191
rect 1978 2188 2310 2191
rect 2538 2188 2566 2191
rect 2826 2188 2838 2191
rect 2938 2188 3246 2191
rect 3266 2188 3766 2191
rect 3774 2188 3838 2191
rect 3874 2188 3894 2191
rect 3914 2188 3974 2191
rect 4058 2188 4086 2191
rect 4274 2188 4294 2191
rect 4306 2188 4390 2191
rect 4658 2188 5078 2191
rect 1206 2182 1209 2188
rect 3774 2182 3777 2188
rect 5182 2182 5185 2188
rect 186 2178 206 2181
rect 210 2178 222 2181
rect 686 2178 694 2181
rect 698 2178 966 2181
rect 1090 2178 1126 2181
rect 1226 2178 1318 2181
rect 1450 2178 1486 2181
rect 1730 2178 1742 2181
rect 1994 2178 2270 2181
rect 2330 2178 2710 2181
rect 2802 2178 2942 2181
rect 3154 2178 3174 2181
rect 3226 2178 3254 2181
rect 3430 2178 3438 2181
rect 3442 2178 3710 2181
rect 3826 2178 3926 2181
rect 3938 2178 4774 2181
rect 4786 2178 4945 2181
rect 5002 2178 5177 2181
rect 178 2168 206 2171
rect 358 2171 361 2178
rect 1566 2172 1569 2178
rect 1590 2172 1593 2178
rect 358 2168 446 2171
rect 690 2168 774 2171
rect 1050 2168 1246 2171
rect 1482 2168 1558 2171
rect 1682 2168 1686 2171
rect 1706 2168 1718 2171
rect 1746 2168 1750 2171
rect 1842 2168 1910 2171
rect 2106 2168 2182 2171
rect 2238 2168 2262 2171
rect 2322 2168 2334 2171
rect 2338 2168 2438 2171
rect 2554 2168 2574 2171
rect 2610 2168 2614 2171
rect 3142 2171 3145 2178
rect 4942 2172 4945 2178
rect 3142 2168 3278 2171
rect 3282 2168 3390 2171
rect 3394 2168 3470 2171
rect 3474 2168 3534 2171
rect 3538 2168 3598 2171
rect 3602 2168 3630 2171
rect 3722 2168 3822 2171
rect 3826 2168 3950 2171
rect 3962 2168 4462 2171
rect 4946 2168 5014 2171
rect 5082 2168 5094 2171
rect 5174 2171 5177 2178
rect 5286 2172 5289 2178
rect 5098 2168 5137 2171
rect 5174 2168 5254 2171
rect 154 2158 238 2161
rect 306 2158 334 2161
rect 354 2158 662 2161
rect 690 2158 718 2161
rect 722 2158 742 2161
rect 846 2158 854 2161
rect 858 2158 934 2161
rect 1006 2158 1249 2161
rect 1258 2158 1278 2161
rect 1282 2158 1406 2161
rect 1410 2158 1670 2161
rect 1698 2158 1846 2161
rect 1898 2158 1910 2161
rect 1962 2158 1966 2161
rect 2034 2158 2094 2161
rect 2134 2158 2198 2161
rect 2238 2161 2241 2168
rect 2302 2162 2305 2168
rect 2210 2158 2241 2161
rect 2250 2158 2254 2161
rect 2482 2158 2862 2161
rect 3242 2158 3246 2161
rect 3266 2158 3302 2161
rect 3306 2158 3358 2161
rect 3362 2158 3382 2161
rect 3842 2158 4094 2161
rect 4242 2158 4494 2161
rect 4662 2161 4665 2168
rect 5030 2162 5033 2168
rect 5134 2162 5137 2168
rect 4546 2158 4665 2161
rect 4674 2158 4710 2161
rect 4714 2158 4822 2161
rect 4898 2158 4910 2161
rect 4994 2158 5022 2161
rect 5090 2158 5094 2161
rect 122 2148 193 2151
rect 386 2148 854 2151
rect 1006 2151 1009 2158
rect 858 2148 1009 2151
rect 1026 2148 1086 2151
rect 1170 2148 1214 2151
rect 1246 2151 1249 2158
rect 1246 2148 1350 2151
rect 1370 2148 1390 2151
rect 1394 2148 1414 2151
rect 1562 2148 1566 2151
rect 1570 2148 1638 2151
rect 1738 2148 1750 2151
rect 1866 2148 1870 2151
rect 1890 2148 1982 2151
rect 2134 2151 2137 2158
rect 2098 2148 2137 2151
rect 2154 2148 2182 2151
rect 2186 2148 2230 2151
rect 2322 2148 2446 2151
rect 2466 2148 2510 2151
rect 2570 2148 2622 2151
rect 2626 2148 2654 2151
rect 2658 2148 2718 2151
rect 2758 2148 2782 2151
rect 2874 2148 2918 2151
rect 2974 2151 2977 2158
rect 2922 2148 2977 2151
rect 3054 2151 3057 2158
rect 3010 2148 3057 2151
rect 3242 2148 3302 2151
rect 3314 2148 3318 2151
rect 3350 2148 3358 2151
rect 3546 2148 3734 2151
rect 3866 2148 3886 2151
rect 3914 2148 3942 2151
rect 4050 2148 4118 2151
rect 4178 2148 4206 2151
rect 4258 2148 4286 2151
rect 4306 2148 4310 2151
rect 4378 2148 4438 2151
rect 4442 2148 4446 2151
rect 4502 2151 4505 2158
rect 4502 2148 4574 2151
rect 4618 2148 4678 2151
rect 4714 2148 4774 2151
rect 4786 2148 4814 2151
rect 4818 2148 4830 2151
rect 4850 2148 4878 2151
rect 4882 2148 4910 2151
rect 4922 2148 4966 2151
rect 5026 2148 5110 2151
rect 5146 2148 5166 2151
rect 5174 2151 5177 2158
rect 5174 2148 5182 2151
rect 190 2142 193 2148
rect 290 2138 422 2141
rect 490 2138 550 2141
rect 570 2138 662 2141
rect 666 2138 670 2141
rect 790 2138 822 2141
rect 826 2138 862 2141
rect 938 2138 1070 2141
rect 1114 2138 1214 2141
rect 1230 2141 1233 2148
rect 1230 2138 1238 2141
rect 1454 2141 1457 2148
rect 1250 2138 1457 2141
rect 1538 2138 1542 2141
rect 1610 2138 1638 2141
rect 1674 2138 1902 2141
rect 1914 2138 1926 2141
rect 1938 2138 1958 2141
rect 2058 2138 2254 2141
rect 2266 2138 2270 2141
rect 2278 2141 2281 2148
rect 2302 2142 2305 2148
rect 2758 2142 2761 2148
rect 3350 2142 3353 2148
rect 3830 2142 3833 2148
rect 3838 2142 3841 2148
rect 2278 2138 2286 2141
rect 2346 2138 2350 2141
rect 2354 2138 2494 2141
rect 2546 2138 2614 2141
rect 2674 2138 2702 2141
rect 2706 2138 2758 2141
rect 2770 2138 3126 2141
rect 3218 2138 3222 2141
rect 3282 2138 3286 2141
rect 3298 2138 3302 2141
rect 3706 2138 3790 2141
rect 3882 2138 3886 2141
rect 3890 2138 3966 2141
rect 3986 2138 4062 2141
rect 4186 2138 4190 2141
rect 4194 2138 4246 2141
rect 4290 2138 4382 2141
rect 4410 2138 4646 2141
rect 4730 2138 4918 2141
rect 4922 2138 5054 2141
rect 5058 2138 5126 2141
rect 5146 2138 5150 2141
rect 734 2132 737 2138
rect 790 2132 793 2138
rect 114 2128 174 2131
rect 178 2128 286 2131
rect 1010 2128 1145 2131
rect 1274 2128 1374 2131
rect 1402 2128 1430 2131
rect 1434 2128 1518 2131
rect 1602 2128 1606 2131
rect 1666 2128 1694 2131
rect 1714 2128 1758 2131
rect 1762 2128 1838 2131
rect 1946 2128 2030 2131
rect 2274 2128 2334 2131
rect 2370 2128 2470 2131
rect 2474 2128 2558 2131
rect 2786 2128 3182 2131
rect 3186 2128 3214 2131
rect 3494 2131 3497 2138
rect 3338 2128 3497 2131
rect 3594 2128 4254 2131
rect 4258 2128 4454 2131
rect 4458 2128 4462 2131
rect 4474 2128 4534 2131
rect 4602 2128 4750 2131
rect 4770 2128 4998 2131
rect 5050 2128 5118 2131
rect 5190 2131 5193 2138
rect 5186 2128 5193 2131
rect 1142 2122 1145 2128
rect 290 2118 310 2121
rect 362 2118 670 2121
rect 674 2118 750 2121
rect 770 2118 846 2121
rect 850 2118 1030 2121
rect 1274 2118 1342 2121
rect 1394 2118 1526 2121
rect 1546 2118 1574 2121
rect 1578 2118 1654 2121
rect 1718 2118 2294 2121
rect 2442 2118 2473 2121
rect 2538 2118 2558 2121
rect 2754 2118 2758 2121
rect 2946 2118 2966 2121
rect 2970 2118 3062 2121
rect 3074 2118 3078 2121
rect 3170 2118 3174 2121
rect 3202 2118 3238 2121
rect 3258 2118 3710 2121
rect 3826 2118 4006 2121
rect 4018 2118 4030 2121
rect 4034 2118 4142 2121
rect 4146 2118 4342 2121
rect 4346 2118 4526 2121
rect 4530 2118 4622 2121
rect 4682 2118 5110 2121
rect 450 2108 638 2111
rect 802 2108 838 2111
rect 1314 2108 1358 2111
rect 1458 2108 1494 2111
rect 1718 2111 1721 2118
rect 1602 2108 1721 2111
rect 1730 2108 1798 2111
rect 1898 2108 1934 2111
rect 1938 2108 1974 2111
rect 1986 2108 2086 2111
rect 2218 2108 2254 2111
rect 2258 2108 2294 2111
rect 2314 2108 2318 2111
rect 2434 2108 2438 2111
rect 2442 2108 2462 2111
rect 2470 2111 2473 2118
rect 5110 2112 5113 2118
rect 2470 2108 2766 2111
rect 2922 2108 3017 2111
rect 3026 2108 3118 2111
rect 3122 2108 3182 2111
rect 3226 2108 3398 2111
rect 3618 2108 3670 2111
rect 3698 2108 3734 2111
rect 3802 2108 3814 2111
rect 3818 2108 3886 2111
rect 3946 2108 4198 2111
rect 4290 2108 4374 2111
rect 4386 2108 4390 2111
rect 4514 2108 4630 2111
rect 4650 2108 4726 2111
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 862 2103 864 2107
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1886 2103 1888 2107
rect 2888 2103 2890 2107
rect 2894 2103 2897 2107
rect 2902 2103 2904 2107
rect 258 2098 302 2101
rect 306 2098 342 2101
rect 466 2098 542 2101
rect 546 2098 566 2101
rect 578 2098 758 2101
rect 1066 2098 1086 2101
rect 1090 2098 1606 2101
rect 1642 2098 1734 2101
rect 1906 2098 1966 2101
rect 2218 2098 2406 2101
rect 2418 2098 2430 2101
rect 2490 2098 2582 2101
rect 2650 2098 2758 2101
rect 2818 2098 2830 2101
rect 2962 2098 3006 2101
rect 3014 2101 3017 2108
rect 3920 2103 3922 2107
rect 3926 2103 3929 2107
rect 3934 2103 3936 2107
rect 4936 2103 4938 2107
rect 4942 2103 4945 2107
rect 4950 2103 4952 2107
rect 5102 2102 5105 2108
rect 5222 2102 5225 2108
rect 3014 2098 3166 2101
rect 3250 2098 3358 2101
rect 3458 2098 3462 2101
rect 3618 2098 3758 2101
rect 3810 2098 3910 2101
rect 3970 2098 4094 2101
rect 4250 2098 4446 2101
rect 4450 2098 4454 2101
rect 4498 2098 4590 2101
rect 4594 2098 4662 2101
rect 530 2088 542 2091
rect 730 2088 838 2091
rect 882 2088 1022 2091
rect 1066 2088 1158 2091
rect 1162 2088 1334 2091
rect 1426 2088 1526 2091
rect 1794 2088 1862 2091
rect 1970 2088 1998 2091
rect 2246 2088 2958 2091
rect 3050 2088 3102 2091
rect 3146 2088 3150 2091
rect 3154 2088 3206 2091
rect 3258 2088 3286 2091
rect 3342 2088 3350 2091
rect 3354 2088 3366 2091
rect 3394 2088 3422 2091
rect 3682 2088 3726 2091
rect 3810 2088 3889 2091
rect 3898 2088 4214 2091
rect 4306 2088 4358 2091
rect 4370 2088 4446 2091
rect 4466 2088 4862 2091
rect 5050 2088 5081 2091
rect 5130 2088 5254 2091
rect 170 2078 294 2081
rect 298 2078 390 2081
rect 394 2078 526 2081
rect 550 2081 553 2088
rect 530 2078 553 2081
rect 558 2081 561 2088
rect 1582 2082 1585 2088
rect 558 2078 582 2081
rect 794 2078 822 2081
rect 826 2078 878 2081
rect 930 2078 934 2081
rect 938 2078 1006 2081
rect 1018 2078 1110 2081
rect 1114 2078 1198 2081
rect 1202 2078 1214 2081
rect 1238 2078 1246 2081
rect 1250 2078 1254 2081
rect 1370 2078 1494 2081
rect 1618 2078 1622 2081
rect 1650 2078 1758 2081
rect 1770 2078 1918 2081
rect 1930 2078 1934 2081
rect 1938 2078 1982 2081
rect 2238 2081 2241 2088
rect 2234 2078 2241 2081
rect 2246 2082 2249 2088
rect 2274 2078 2366 2081
rect 2426 2078 2446 2081
rect 2466 2078 2470 2081
rect 2626 2078 2694 2081
rect 2818 2078 2902 2081
rect 2966 2081 2969 2088
rect 2966 2078 3102 2081
rect 3178 2078 3190 2081
rect 3194 2078 3430 2081
rect 3434 2078 3518 2081
rect 3618 2078 3622 2081
rect 3682 2078 3686 2081
rect 3762 2078 3766 2081
rect 3778 2078 3822 2081
rect 3886 2081 3889 2088
rect 3886 2078 4030 2081
rect 4058 2078 4062 2081
rect 4106 2078 4169 2081
rect 4238 2081 4241 2088
rect 4194 2078 4334 2081
rect 4418 2078 4470 2081
rect 4482 2078 4486 2081
rect 4498 2078 4510 2081
rect 4626 2078 4734 2081
rect 5022 2078 5070 2081
rect 5078 2081 5081 2088
rect 5078 2078 5158 2081
rect 5202 2078 5230 2081
rect 1558 2072 1561 2078
rect 1566 2072 1569 2078
rect 70 2068 89 2071
rect 258 2068 270 2071
rect 274 2068 382 2071
rect 386 2068 1126 2071
rect 1130 2068 1142 2071
rect 1178 2068 1190 2071
rect 1226 2068 1238 2071
rect 1310 2068 1318 2071
rect 1338 2068 1406 2071
rect 1450 2068 1558 2071
rect 1578 2068 1774 2071
rect 1778 2068 1870 2071
rect 1890 2068 1894 2071
rect 1922 2068 1977 2071
rect 1986 2068 1998 2071
rect 2150 2071 2153 2078
rect 2750 2072 2753 2078
rect 4166 2072 4169 2078
rect 2042 2068 2153 2071
rect 2162 2068 2166 2071
rect 2298 2068 2326 2071
rect 2330 2068 2358 2071
rect 2370 2068 2502 2071
rect 2642 2068 2742 2071
rect 2826 2068 2870 2071
rect 2882 2068 2926 2071
rect 2930 2068 3374 2071
rect 3410 2068 3414 2071
rect 3466 2068 3529 2071
rect 3538 2068 3902 2071
rect 4042 2068 4046 2071
rect 4146 2068 4150 2071
rect 4178 2068 4198 2071
rect 4226 2068 4238 2071
rect 4346 2068 4350 2071
rect 4410 2068 4542 2071
rect 4738 2068 4742 2071
rect 4830 2068 4886 2071
rect 5022 2071 5025 2078
rect 5018 2068 5025 2071
rect 5042 2068 5086 2071
rect 5194 2068 5222 2071
rect 5274 2068 5278 2071
rect 70 2062 73 2068
rect 86 2062 89 2068
rect 1206 2062 1209 2068
rect 1246 2062 1249 2068
rect 1310 2062 1313 2068
rect 122 2058 190 2061
rect 310 2058 398 2061
rect 402 2058 606 2061
rect 614 2058 774 2061
rect 802 2058 806 2061
rect 810 2058 822 2061
rect 826 2058 878 2061
rect 906 2058 910 2061
rect 954 2058 958 2061
rect 1026 2058 1134 2061
rect 1218 2058 1230 2061
rect 1330 2058 1366 2061
rect 1378 2058 1382 2061
rect 1426 2058 1430 2061
rect 1498 2058 1510 2061
rect 1554 2058 1625 2061
rect 1634 2058 1662 2061
rect 1698 2058 1782 2061
rect 1850 2058 1854 2061
rect 1974 2061 1977 2068
rect 1974 2058 2062 2061
rect 2066 2058 2078 2061
rect 2106 2058 2134 2061
rect 2154 2058 2414 2061
rect 2458 2058 2574 2061
rect 2630 2058 2681 2061
rect 2698 2058 2702 2061
rect 2714 2058 2734 2061
rect 2826 2058 2918 2061
rect 2922 2058 3118 2061
rect 3122 2058 3166 2061
rect 3218 2058 3238 2061
rect 3290 2058 3297 2061
rect 3330 2058 3342 2061
rect 3410 2058 3454 2061
rect 3458 2058 3478 2061
rect 3526 2061 3529 2068
rect 3526 2058 3550 2061
rect 3602 2058 3606 2061
rect 3650 2058 3702 2061
rect 3722 2058 3726 2061
rect 3746 2058 3766 2061
rect 3842 2058 3894 2061
rect 3902 2061 3905 2068
rect 3902 2058 4006 2061
rect 4010 2058 4014 2061
rect 4026 2058 4062 2061
rect 4098 2058 4142 2061
rect 4194 2058 4398 2061
rect 4490 2058 4518 2061
rect 4522 2058 4529 2061
rect 4566 2061 4569 2068
rect 4546 2058 4569 2061
rect 4614 2062 4617 2068
rect 4654 2061 4657 2068
rect 4678 2062 4681 2068
rect 4830 2062 4833 2068
rect 4642 2058 4657 2061
rect 4666 2058 4670 2061
rect 4722 2058 4798 2061
rect 4994 2058 4998 2061
rect 5050 2058 5054 2061
rect 5082 2058 5110 2061
rect 5114 2058 5286 2061
rect 310 2052 313 2058
rect 614 2052 617 2058
rect 1182 2052 1185 2058
rect 186 2048 222 2051
rect 242 2048 246 2051
rect 498 2048 502 2051
rect 634 2048 638 2051
rect 698 2048 766 2051
rect 814 2048 822 2051
rect 906 2048 926 2051
rect 1218 2048 1574 2051
rect 1622 2051 1625 2058
rect 2630 2052 2633 2058
rect 2678 2052 2681 2058
rect 3294 2052 3297 2058
rect 1622 2048 1726 2051
rect 1730 2048 1830 2051
rect 1842 2048 1918 2051
rect 1938 2048 1942 2051
rect 1946 2048 1982 2051
rect 2018 2048 2110 2051
rect 2130 2048 2166 2051
rect 2234 2048 2294 2051
rect 2410 2048 2510 2051
rect 2514 2048 2598 2051
rect 2850 2048 2926 2051
rect 2954 2048 2958 2051
rect 3066 2048 3134 2051
rect 3210 2048 3222 2051
rect 3242 2048 3254 2051
rect 3370 2048 3382 2051
rect 3386 2048 3510 2051
rect 3514 2048 3638 2051
rect 3690 2048 3694 2051
rect 3790 2051 3793 2058
rect 3730 2048 3793 2051
rect 3810 2048 4046 2051
rect 4146 2048 4158 2051
rect 4234 2048 4238 2051
rect 4350 2048 4369 2051
rect 202 2038 350 2041
rect 354 2038 558 2041
rect 682 2038 710 2041
rect 798 2041 801 2048
rect 714 2038 801 2041
rect 814 2042 817 2048
rect 954 2038 1142 2041
rect 1146 2038 1190 2041
rect 1362 2038 1390 2041
rect 1394 2038 1446 2041
rect 1838 2038 1846 2041
rect 1850 2038 1854 2041
rect 1926 2041 1929 2048
rect 4350 2042 4353 2048
rect 4366 2042 4369 2048
rect 4490 2048 4502 2051
rect 4514 2048 4542 2051
rect 4602 2048 4630 2051
rect 4634 2048 4750 2051
rect 5018 2048 5089 2051
rect 1926 2038 1950 2041
rect 1966 2038 1974 2041
rect 1978 2038 2030 2041
rect 2146 2038 2494 2041
rect 2498 2038 2526 2041
rect 2546 2038 2926 2041
rect 2950 2038 2958 2041
rect 2962 2038 3022 2041
rect 3074 2038 3086 2041
rect 3090 2038 3174 2041
rect 3366 2038 3374 2041
rect 3378 2038 3609 2041
rect 3618 2038 3654 2041
rect 3746 2038 3846 2041
rect 3850 2038 3854 2041
rect 3882 2038 3886 2041
rect 4130 2038 4142 2041
rect 4406 2041 4409 2048
rect 4582 2042 4585 2048
rect 5086 2042 5089 2048
rect 4386 2038 4409 2041
rect 4498 2038 4518 2041
rect 4658 2038 4710 2041
rect 378 2028 662 2031
rect 666 2028 750 2031
rect 754 2028 1102 2031
rect 1174 2028 1182 2031
rect 1186 2028 1294 2031
rect 1410 2028 1422 2031
rect 1522 2028 1614 2031
rect 1686 2031 1689 2038
rect 1686 2028 1814 2031
rect 1818 2028 1934 2031
rect 1938 2028 1942 2031
rect 2034 2028 2102 2031
rect 2114 2028 2254 2031
rect 2346 2028 2390 2031
rect 2394 2028 2574 2031
rect 2602 2028 2742 2031
rect 2746 2028 2774 2031
rect 2850 2028 3502 2031
rect 3606 2031 3609 2038
rect 3606 2028 3694 2031
rect 3982 2031 3985 2038
rect 3826 2028 4030 2031
rect 4058 2028 4150 2031
rect 4226 2028 4654 2031
rect 4978 2028 5030 2031
rect 5034 2028 5102 2031
rect 266 2018 686 2021
rect 1098 2018 1230 2021
rect 1338 2018 1582 2021
rect 1586 2018 2262 2021
rect 2266 2018 2294 2021
rect 2310 2018 2318 2021
rect 2322 2018 2518 2021
rect 2578 2018 2854 2021
rect 2858 2018 2966 2021
rect 3202 2018 3334 2021
rect 3394 2018 3870 2021
rect 3874 2018 4486 2021
rect 4874 2018 4990 2021
rect 5034 2018 5246 2021
rect 230 2012 233 2018
rect 906 2008 1166 2011
rect 1426 2008 1470 2011
rect 1474 2008 1534 2011
rect 1690 2008 1694 2011
rect 1718 2008 1942 2011
rect 2010 2008 2094 2011
rect 2130 2008 2374 2011
rect 2522 2008 2566 2011
rect 2570 2008 2582 2011
rect 2586 2008 2662 2011
rect 2810 2008 2814 2011
rect 3106 2008 3150 2011
rect 3154 2008 3278 2011
rect 3474 2008 3526 2011
rect 4002 2008 4398 2011
rect 4706 2008 4862 2011
rect 328 2003 330 2007
rect 334 2003 337 2007
rect 342 2003 344 2007
rect 1352 2003 1354 2007
rect 1358 2003 1361 2007
rect 1366 2003 1368 2007
rect 194 1998 318 2001
rect 818 1998 886 2001
rect 994 1998 1254 2001
rect 1718 2001 1721 2008
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2398 2003 2400 2007
rect 3400 2003 3402 2007
rect 3406 2003 3409 2007
rect 3414 2003 3416 2007
rect 4424 2003 4426 2007
rect 4430 2003 4433 2007
rect 4438 2003 4440 2007
rect 1522 1998 1721 2001
rect 1730 1998 2134 2001
rect 2690 1998 2854 2001
rect 2858 1998 3102 2001
rect 3106 1998 3230 2001
rect 3234 1998 3254 2001
rect 3298 1998 3326 2001
rect 3786 1998 4078 2001
rect 4138 1998 4222 2001
rect 4362 1998 4366 2001
rect 4722 1998 4726 2001
rect 4730 1998 4926 2001
rect 1470 1992 1473 1998
rect 178 1988 286 1991
rect 334 1988 342 1991
rect 346 1988 486 1991
rect 762 1988 902 1991
rect 1130 1988 1158 1991
rect 1210 1988 1462 1991
rect 1586 1988 1790 1991
rect 1794 1988 1830 1991
rect 1842 1988 1846 1991
rect 1866 1988 1902 1991
rect 2098 1988 2118 1991
rect 2186 1988 2342 1991
rect 2434 1988 2502 1991
rect 2506 1988 2630 1991
rect 2634 1988 2686 1991
rect 2690 1988 2710 1991
rect 3242 1988 3526 1991
rect 4082 1988 4094 1991
rect 4114 1988 4785 1991
rect 62 1981 65 1988
rect 62 1978 470 1981
rect 834 1978 1190 1981
rect 1218 1978 1342 1981
rect 1530 1978 1566 1981
rect 1762 1978 1998 1981
rect 2002 1978 2550 1981
rect 2554 1978 2822 1981
rect 3126 1981 3129 1988
rect 4782 1982 4785 1988
rect 3126 1978 3318 1981
rect 3378 1978 3438 1981
rect 3482 1978 3542 1981
rect 3626 1978 3630 1981
rect 3690 1978 3950 1981
rect 3954 1978 3982 1981
rect 4042 1978 4086 1981
rect 4202 1978 4478 1981
rect 4834 1978 4854 1981
rect 4986 1978 5286 1981
rect 4870 1972 4873 1978
rect 230 1968 286 1971
rect 426 1968 430 1971
rect 634 1968 694 1971
rect 762 1968 782 1971
rect 794 1968 862 1971
rect 866 1968 1126 1971
rect 1162 1968 1398 1971
rect 1426 1968 1430 1971
rect 1458 1968 1558 1971
rect 1586 1968 1606 1971
rect 1618 1968 1742 1971
rect 1754 1968 1774 1971
rect 1786 1968 1798 1971
rect 1818 1968 1830 1971
rect 1834 1968 1870 1971
rect 2002 1968 2070 1971
rect 2106 1968 2126 1971
rect 2130 1968 2230 1971
rect 2242 1968 2246 1971
rect 2418 1968 2454 1971
rect 2474 1968 2478 1971
rect 2490 1968 2542 1971
rect 2562 1968 2574 1971
rect 2754 1968 2766 1971
rect 2794 1968 2838 1971
rect 3034 1968 3070 1971
rect 3242 1968 3262 1971
rect 3426 1968 3430 1971
rect 3458 1968 3582 1971
rect 3906 1968 4198 1971
rect 4202 1968 4302 1971
rect 4418 1968 4502 1971
rect 4570 1968 4630 1971
rect 4858 1968 4862 1971
rect 5026 1968 5265 1971
rect 230 1962 233 1968
rect 1438 1962 1441 1968
rect 2078 1962 2081 1968
rect 258 1958 270 1961
rect 278 1958 406 1961
rect 618 1958 654 1961
rect 658 1958 894 1961
rect 946 1958 982 1961
rect 986 1958 1206 1961
rect 1322 1958 1374 1961
rect 1410 1958 1414 1961
rect 1450 1958 2006 1961
rect 2058 1958 2062 1961
rect 2298 1958 2406 1961
rect 2450 1958 2590 1961
rect 2598 1961 2601 1968
rect 2918 1962 2921 1968
rect 2598 1958 2670 1961
rect 2674 1958 2678 1961
rect 2698 1958 2782 1961
rect 2802 1958 2806 1961
rect 2934 1961 2937 1968
rect 5262 1962 5265 1968
rect 2934 1958 3054 1961
rect 3062 1958 3078 1961
rect 3086 1958 3094 1961
rect 3098 1958 3158 1961
rect 3186 1958 3190 1961
rect 3226 1958 3278 1961
rect 3426 1958 3670 1961
rect 3674 1958 3998 1961
rect 4018 1958 4110 1961
rect 4314 1958 4318 1961
rect 4322 1958 4342 1961
rect 4370 1958 4606 1961
rect 4714 1958 4790 1961
rect 4826 1958 5062 1961
rect 278 1952 281 1958
rect 3062 1952 3065 1958
rect 130 1948 182 1951
rect 226 1948 254 1951
rect 322 1948 326 1951
rect 402 1948 646 1951
rect 658 1948 766 1951
rect 810 1948 998 1951
rect 1002 1948 1054 1951
rect 1074 1948 1118 1951
rect 1130 1948 1190 1951
rect 1194 1948 1262 1951
rect 1266 1948 1582 1951
rect 1610 1948 1614 1951
rect 1626 1948 1630 1951
rect 1698 1948 1702 1951
rect 1754 1948 1854 1951
rect 1874 1948 2006 1951
rect 2026 1948 2078 1951
rect 2114 1948 2126 1951
rect 2130 1948 2262 1951
rect 2370 1948 2414 1951
rect 2418 1948 2438 1951
rect 2442 1948 2486 1951
rect 2506 1948 2518 1951
rect 2586 1948 2614 1951
rect 2618 1948 2662 1951
rect 2666 1948 2753 1951
rect 2778 1948 2782 1951
rect 2938 1948 2969 1951
rect 3034 1948 3062 1951
rect 3082 1948 3118 1951
rect 3122 1948 3406 1951
rect 3418 1948 3438 1951
rect 3642 1948 3718 1951
rect 18 1938 334 1941
rect 578 1938 582 1941
rect 594 1938 865 1941
rect 874 1938 966 1941
rect 1122 1938 1198 1941
rect 1218 1938 1246 1941
rect 1322 1938 1342 1941
rect 1346 1938 1350 1941
rect 1354 1938 1438 1941
rect 1506 1938 1622 1941
rect 1626 1938 1654 1941
rect 1706 1938 1710 1941
rect 1722 1938 1726 1941
rect 1778 1938 1854 1941
rect 1882 1938 1886 1941
rect 1898 1938 1910 1941
rect 1970 1938 1974 1941
rect 2010 1938 2014 1941
rect 2114 1938 2118 1941
rect 2234 1938 2574 1941
rect 2674 1938 2678 1941
rect 2682 1938 2702 1941
rect 2738 1938 2742 1941
rect 2750 1941 2753 1948
rect 2814 1941 2817 1948
rect 2966 1942 2969 1948
rect 3606 1942 3609 1948
rect 3730 1948 3774 1951
rect 4046 1948 4054 1951
rect 4058 1948 4158 1951
rect 4270 1948 4318 1951
rect 4370 1948 4550 1951
rect 4642 1948 5014 1951
rect 5018 1948 5046 1951
rect 5234 1948 5278 1951
rect 2750 1938 2894 1941
rect 2898 1938 2910 1941
rect 3074 1938 3198 1941
rect 3266 1938 3270 1941
rect 3426 1938 3446 1941
rect 3546 1938 3550 1941
rect 3610 1938 4054 1941
rect 4066 1938 4070 1941
rect 4082 1938 4086 1941
rect 4114 1938 4126 1941
rect 4190 1941 4193 1948
rect 4262 1941 4265 1948
rect 4190 1938 4265 1941
rect 4270 1942 4273 1948
rect 4598 1941 4601 1948
rect 4514 1938 4601 1941
rect 4770 1938 4838 1941
rect 4858 1938 4918 1941
rect 5042 1938 5126 1941
rect 5150 1938 5214 1941
rect 670 1932 673 1938
rect 862 1932 865 1938
rect 1926 1932 1929 1938
rect 2062 1932 2065 1938
rect 2086 1932 2089 1938
rect 226 1928 398 1931
rect 638 1928 646 1931
rect 650 1928 662 1931
rect 698 1928 806 1931
rect 866 1928 934 1931
rect 938 1928 1006 1931
rect 1034 1928 1086 1931
rect 1090 1928 1134 1931
rect 1146 1928 1182 1931
rect 1186 1928 1406 1931
rect 1546 1928 1582 1931
rect 1594 1928 1598 1931
rect 1698 1928 1702 1931
rect 1706 1928 1718 1931
rect 1746 1928 1870 1931
rect 1898 1928 1918 1931
rect 1946 1928 1950 1931
rect 1954 1928 2006 1931
rect 2130 1928 2142 1931
rect 2258 1928 2334 1931
rect 2362 1928 2502 1931
rect 2514 1928 2526 1931
rect 2554 1928 2614 1931
rect 2634 1928 2646 1931
rect 2650 1928 2790 1931
rect 2794 1928 2798 1931
rect 2818 1928 2902 1931
rect 3114 1928 3150 1931
rect 3290 1928 3318 1931
rect 3366 1931 3369 1938
rect 3366 1928 3462 1931
rect 3582 1931 3585 1938
rect 4094 1932 4097 1938
rect 4566 1932 4569 1938
rect 5150 1932 5153 1938
rect 3582 1928 3630 1931
rect 3674 1928 3678 1931
rect 3866 1928 3870 1931
rect 3882 1928 4006 1931
rect 4378 1928 4558 1931
rect 4754 1928 4998 1931
rect 5002 1928 5006 1931
rect 5010 1928 5150 1931
rect 5262 1931 5265 1938
rect 5262 1928 5294 1931
rect 222 1922 225 1928
rect 278 1918 286 1921
rect 290 1918 318 1921
rect 506 1918 766 1921
rect 962 1918 1126 1921
rect 1194 1918 1278 1921
rect 1314 1918 1334 1921
rect 1338 1918 1398 1921
rect 1402 1918 1422 1921
rect 1638 1921 1641 1928
rect 1474 1918 1641 1921
rect 1710 1918 1718 1921
rect 1722 1918 2033 1921
rect 2162 1918 2262 1921
rect 2334 1921 2337 1928
rect 2334 1918 2438 1921
rect 2562 1918 2606 1921
rect 2658 1918 2766 1921
rect 2786 1918 2862 1921
rect 3098 1918 3142 1921
rect 3314 1918 3398 1921
rect 3474 1918 3494 1921
rect 3498 1918 3550 1921
rect 3554 1918 3678 1921
rect 3682 1918 3798 1921
rect 3866 1918 3886 1921
rect 3898 1918 4102 1921
rect 4394 1918 4598 1921
rect 4898 1918 4926 1921
rect 4930 1918 5046 1921
rect 5098 1918 5126 1921
rect 5138 1918 5142 1921
rect 5154 1918 5182 1921
rect 122 1908 142 1911
rect 146 1908 382 1911
rect 402 1908 422 1911
rect 458 1908 782 1911
rect 1138 1908 1862 1911
rect 2030 1911 2033 1918
rect 2870 1912 2873 1918
rect 2030 1908 2086 1911
rect 2158 1908 2326 1911
rect 2426 1908 2718 1911
rect 2738 1908 2862 1911
rect 3066 1908 3230 1911
rect 3282 1908 3454 1911
rect 3650 1908 3702 1911
rect 3810 1908 3862 1911
rect 3970 1908 4070 1911
rect 4074 1908 4142 1911
rect 4154 1908 4614 1911
rect 4618 1908 4638 1911
rect 4794 1908 4918 1911
rect 4986 1908 5062 1911
rect 5074 1908 5190 1911
rect 5226 1908 5238 1911
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 862 1903 864 1907
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1886 1903 1888 1907
rect 102 1898 838 1901
rect 1026 1898 1030 1901
rect 1082 1898 1110 1901
rect 1114 1898 1118 1901
rect 1154 1898 1358 1901
rect 1370 1898 1374 1901
rect 1378 1898 1422 1901
rect 1530 1898 1670 1901
rect 1778 1898 1830 1901
rect 1930 1898 1934 1901
rect 2158 1901 2161 1908
rect 2888 1903 2890 1907
rect 2894 1903 2897 1907
rect 2902 1903 2904 1907
rect 3920 1903 3922 1907
rect 3926 1903 3929 1907
rect 3934 1903 3936 1907
rect 3942 1902 3945 1908
rect 4936 1903 4938 1907
rect 4942 1903 4945 1907
rect 4950 1903 4952 1907
rect 2042 1898 2161 1901
rect 2218 1898 2222 1901
rect 2226 1898 2278 1901
rect 2418 1898 2446 1901
rect 2474 1898 2486 1901
rect 2578 1898 2702 1901
rect 2706 1898 2710 1901
rect 2922 1898 2974 1901
rect 3186 1898 3190 1901
rect 3282 1898 3294 1901
rect 3386 1898 3526 1901
rect 3562 1898 3598 1901
rect 3602 1898 3662 1901
rect 3674 1898 3686 1901
rect 3954 1898 3974 1901
rect 3994 1898 4174 1901
rect 4186 1898 4190 1901
rect 4290 1898 4342 1901
rect 4346 1898 4414 1901
rect 4418 1898 4446 1901
rect 4474 1898 4630 1901
rect 4854 1898 4878 1901
rect 4958 1898 5166 1901
rect 5170 1898 5278 1901
rect 6 1891 9 1898
rect 102 1892 105 1898
rect 2166 1892 2169 1898
rect 4846 1892 4849 1898
rect 4854 1892 4857 1898
rect 6 1888 102 1891
rect 258 1888 318 1891
rect 598 1888 606 1891
rect 610 1888 710 1891
rect 1014 1888 1022 1891
rect 1026 1888 1070 1891
rect 1090 1888 1446 1891
rect 1450 1888 1718 1891
rect 1866 1888 2046 1891
rect 2058 1888 2062 1891
rect 2074 1888 2166 1891
rect 2274 1888 2286 1891
rect 2330 1888 2334 1891
rect 2346 1888 2406 1891
rect 2410 1888 2430 1891
rect 2442 1888 2462 1891
rect 2466 1888 2470 1891
rect 2482 1888 2486 1891
rect 2578 1888 2582 1891
rect 2610 1888 2630 1891
rect 2634 1888 2678 1891
rect 2846 1888 3102 1891
rect 3162 1888 3262 1891
rect 3266 1888 3294 1891
rect 3618 1888 4214 1891
rect 4218 1888 4270 1891
rect 4314 1888 4529 1891
rect 182 1881 185 1888
rect 74 1878 185 1881
rect 266 1878 270 1881
rect 290 1878 310 1881
rect 314 1878 366 1881
rect 386 1878 614 1881
rect 642 1878 702 1881
rect 754 1878 790 1881
rect 842 1878 1102 1881
rect 1146 1878 1198 1881
rect 1210 1878 1270 1881
rect 1274 1878 1310 1881
rect 1354 1878 1454 1881
rect 1554 1878 1566 1881
rect 1570 1878 1614 1881
rect 1626 1878 1726 1881
rect 1730 1878 1790 1881
rect 1866 1878 1990 1881
rect 2234 1878 2270 1881
rect 2274 1878 2550 1881
rect 2562 1878 2766 1881
rect 2790 1881 2793 1888
rect 2846 1882 2849 1888
rect 3614 1882 3617 1888
rect 2790 1878 2846 1881
rect 2874 1878 3038 1881
rect 3138 1878 3294 1881
rect 3578 1878 3598 1881
rect 3642 1878 3678 1881
rect 3690 1878 3750 1881
rect 3786 1878 3966 1881
rect 3970 1878 3998 1881
rect 4018 1878 4102 1881
rect 4114 1878 4193 1881
rect 4294 1881 4297 1888
rect 4210 1878 4297 1881
rect 4526 1882 4529 1888
rect 4762 1888 4806 1891
rect 4958 1891 4961 1898
rect 4930 1888 4961 1891
rect 4982 1888 5014 1891
rect 5122 1888 5161 1891
rect 4534 1882 4537 1888
rect 4590 1882 4593 1888
rect 4982 1882 4985 1888
rect 5158 1882 5161 1888
rect 5166 1882 5169 1888
rect 4818 1878 4822 1881
rect 4826 1878 4958 1881
rect 5010 1878 5142 1881
rect 1318 1872 1321 1878
rect 194 1868 225 1871
rect 290 1868 374 1871
rect 466 1868 510 1871
rect 690 1868 694 1871
rect 818 1868 838 1871
rect 946 1868 1030 1871
rect 1066 1868 1086 1871
rect 1098 1868 1126 1871
rect 1378 1868 1510 1871
rect 1562 1868 1606 1871
rect 1858 1868 1862 1871
rect 2014 1871 2017 1878
rect 1970 1868 2017 1871
rect 2034 1868 2054 1871
rect 2074 1868 2118 1871
rect 2174 1871 2177 1878
rect 3046 1872 3049 1878
rect 2122 1868 2177 1871
rect 2234 1868 2238 1871
rect 2242 1868 2806 1871
rect 2826 1868 2982 1871
rect 3034 1868 3046 1871
rect 3154 1868 3190 1871
rect 3266 1868 3326 1871
rect 3366 1871 3369 1878
rect 4190 1872 4193 1878
rect 3366 1868 3518 1871
rect 3530 1868 3550 1871
rect 3586 1868 3622 1871
rect 3642 1868 3649 1871
rect 3658 1868 3694 1871
rect 3738 1868 3814 1871
rect 3930 1868 3958 1871
rect 3978 1868 4014 1871
rect 4058 1868 4150 1871
rect 4154 1868 4158 1871
rect 4214 1868 4222 1871
rect 4282 1868 4366 1871
rect 4394 1868 4414 1871
rect 4530 1868 4537 1871
rect 4578 1868 4638 1871
rect 4690 1868 4750 1871
rect 4754 1868 5022 1871
rect 5026 1868 5094 1871
rect 5098 1868 5182 1871
rect 5186 1868 5230 1871
rect 5258 1868 5278 1871
rect 70 1858 126 1861
rect 150 1861 153 1868
rect 150 1858 214 1861
rect 222 1861 225 1868
rect 718 1862 721 1868
rect 222 1858 334 1861
rect 354 1858 374 1861
rect 434 1858 510 1861
rect 514 1858 542 1861
rect 610 1858 614 1861
rect 682 1858 686 1861
rect 698 1858 702 1861
rect 770 1858 774 1861
rect 818 1858 878 1861
rect 930 1858 1046 1861
rect 1050 1858 1118 1861
rect 1130 1858 1158 1861
rect 1278 1861 1281 1868
rect 1210 1858 1281 1861
rect 1334 1861 1337 1868
rect 1298 1858 1374 1861
rect 1410 1858 1526 1861
rect 1546 1858 1574 1861
rect 1586 1858 1662 1861
rect 1742 1861 1745 1868
rect 2190 1862 2193 1868
rect 3646 1862 3649 1868
rect 1742 1858 1758 1861
rect 1778 1858 1846 1861
rect 1962 1858 2070 1861
rect 2330 1858 2334 1861
rect 2370 1858 2422 1861
rect 2426 1858 2486 1861
rect 2490 1858 2566 1861
rect 2586 1858 2590 1861
rect 2594 1858 2638 1861
rect 2682 1858 2710 1861
rect 2714 1858 2750 1861
rect 2794 1858 2814 1861
rect 2986 1858 3022 1861
rect 3026 1858 3078 1861
rect 3170 1858 3222 1861
rect 3242 1858 3270 1861
rect 3486 1858 3494 1861
rect 3538 1858 3598 1861
rect 3658 1858 3681 1861
rect 3726 1861 3729 1868
rect 4214 1862 4217 1868
rect 4246 1862 4249 1868
rect 3714 1858 3729 1861
rect 3810 1858 3870 1861
rect 3922 1858 3950 1861
rect 3978 1858 3982 1861
rect 4098 1858 4158 1861
rect 4250 1858 4409 1861
rect 4418 1858 4646 1861
rect 4762 1858 4790 1861
rect 4794 1858 4846 1861
rect 4858 1858 4878 1861
rect 5018 1858 5030 1861
rect 5042 1858 5046 1861
rect 5106 1858 5110 1861
rect 70 1852 73 1858
rect 710 1852 713 1858
rect 210 1848 254 1851
rect 258 1848 358 1851
rect 386 1848 574 1851
rect 578 1848 646 1851
rect 770 1848 846 1851
rect 1002 1848 1094 1851
rect 1298 1848 1326 1851
rect 1570 1848 1606 1851
rect 1610 1848 1622 1851
rect 1634 1848 1694 1851
rect 1698 1848 1718 1851
rect 1722 1848 1894 1851
rect 1946 1848 1990 1851
rect 2026 1848 2030 1851
rect 2210 1848 2470 1851
rect 2506 1848 2510 1851
rect 2546 1848 2550 1851
rect 2570 1848 2614 1851
rect 2666 1848 2670 1851
rect 2778 1848 2870 1851
rect 2882 1848 2886 1851
rect 2890 1848 3038 1851
rect 3094 1851 3097 1858
rect 3486 1852 3489 1858
rect 3678 1852 3681 1858
rect 4022 1852 4025 1858
rect 4406 1852 4409 1858
rect 3094 1848 3142 1851
rect 3154 1848 3182 1851
rect 3218 1848 3222 1851
rect 3506 1848 3510 1851
rect 3514 1848 3670 1851
rect 3710 1848 3774 1851
rect 3778 1848 3790 1851
rect 3834 1848 3878 1851
rect 3982 1848 3990 1851
rect 3994 1848 4014 1851
rect 4066 1848 4254 1851
rect 4562 1848 4582 1851
rect 4654 1848 4670 1851
rect 4714 1848 4790 1851
rect 4794 1848 4870 1851
rect 5042 1848 5222 1851
rect 1126 1842 1129 1848
rect 234 1838 494 1841
rect 562 1838 598 1841
rect 770 1838 822 1841
rect 1294 1841 1297 1848
rect 1266 1838 1297 1841
rect 1346 1838 1590 1841
rect 1594 1838 1686 1841
rect 1754 1838 2190 1841
rect 2194 1838 2358 1841
rect 2434 1838 2454 1841
rect 2458 1838 2518 1841
rect 2550 1841 2553 1848
rect 3710 1842 3713 1848
rect 2550 1838 2582 1841
rect 2586 1838 2630 1841
rect 2634 1838 2654 1841
rect 2658 1838 2686 1841
rect 2770 1838 2830 1841
rect 2858 1838 2910 1841
rect 2946 1838 3006 1841
rect 3026 1838 3038 1841
rect 3442 1838 3502 1841
rect 3850 1838 3870 1841
rect 4178 1838 4342 1841
rect 4614 1841 4617 1848
rect 4538 1838 4617 1841
rect 4654 1842 4657 1848
rect 4982 1842 4985 1848
rect 4698 1838 4769 1841
rect 3870 1832 3873 1838
rect 4766 1832 4769 1838
rect 522 1828 550 1831
rect 554 1828 590 1831
rect 858 1828 1350 1831
rect 1426 1828 1646 1831
rect 1794 1828 2150 1831
rect 2178 1828 2270 1831
rect 2330 1828 2686 1831
rect 2850 1828 2942 1831
rect 3050 1828 3142 1831
rect 3146 1828 3390 1831
rect 3410 1828 3526 1831
rect 3530 1828 3590 1831
rect 3674 1828 3862 1831
rect 4218 1828 4230 1831
rect 4242 1828 4294 1831
rect 4322 1828 4574 1831
rect 4578 1828 4742 1831
rect 4746 1828 4758 1831
rect 4858 1828 5206 1831
rect 66 1818 830 1821
rect 1042 1818 1190 1821
rect 1242 1818 1462 1821
rect 1618 1818 1678 1821
rect 1682 1818 1814 1821
rect 2010 1818 2070 1821
rect 2074 1818 2230 1821
rect 2258 1818 2286 1821
rect 2290 1818 2310 1821
rect 2322 1818 2574 1821
rect 2702 1821 2705 1828
rect 2702 1818 3022 1821
rect 3034 1818 3070 1821
rect 3074 1818 3078 1821
rect 3130 1818 3142 1821
rect 3186 1818 3358 1821
rect 3458 1818 3734 1821
rect 3770 1818 3910 1821
rect 3994 1818 4166 1821
rect 4218 1818 4406 1821
rect 4458 1818 4574 1821
rect 4634 1818 4678 1821
rect 290 1808 318 1811
rect 674 1808 710 1811
rect 714 1808 726 1811
rect 754 1808 774 1811
rect 906 1808 1006 1811
rect 1010 1808 1142 1811
rect 1146 1808 1342 1811
rect 1674 1808 1766 1811
rect 2034 1808 2038 1811
rect 2122 1808 2286 1811
rect 2322 1808 2366 1811
rect 2546 1808 2662 1811
rect 2674 1808 2710 1811
rect 2722 1808 2814 1811
rect 3130 1808 3382 1811
rect 3698 1808 3830 1811
rect 4170 1808 4262 1811
rect 4626 1808 5014 1811
rect 328 1803 330 1807
rect 334 1803 337 1807
rect 342 1803 344 1807
rect 1352 1803 1354 1807
rect 1358 1803 1361 1807
rect 1366 1803 1368 1807
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2398 1803 2400 1807
rect 3400 1803 3402 1807
rect 3406 1803 3409 1807
rect 3414 1803 3416 1807
rect 4424 1803 4426 1807
rect 4430 1803 4433 1807
rect 4438 1803 4440 1807
rect 210 1798 238 1801
rect 522 1798 526 1801
rect 530 1798 958 1801
rect 1098 1798 1134 1801
rect 1162 1798 1174 1801
rect 1178 1798 1310 1801
rect 1562 1798 1838 1801
rect 1938 1798 2046 1801
rect 2098 1798 2150 1801
rect 2154 1798 2222 1801
rect 2450 1798 2494 1801
rect 2626 1798 2950 1801
rect 3034 1798 3054 1801
rect 3082 1798 3238 1801
rect 3586 1798 3878 1801
rect 3882 1798 4182 1801
rect 4546 1798 4710 1801
rect 3070 1792 3073 1798
rect 170 1788 262 1791
rect 430 1788 766 1791
rect 786 1788 2542 1791
rect 2550 1788 2630 1791
rect 2714 1788 2742 1791
rect 2746 1788 2902 1791
rect 3202 1788 3726 1791
rect 4010 1788 4198 1791
rect 4202 1788 4294 1791
rect 4370 1788 4662 1791
rect 430 1782 433 1788
rect 2550 1782 2553 1788
rect 530 1778 582 1781
rect 730 1778 838 1781
rect 1290 1778 1494 1781
rect 2050 1778 2102 1781
rect 2162 1778 2502 1781
rect 2602 1778 2750 1781
rect 2966 1781 2969 1788
rect 2966 1778 3006 1781
rect 3010 1778 3102 1781
rect 3114 1778 3518 1781
rect 3522 1778 3966 1781
rect 3978 1778 4281 1781
rect 4354 1778 4382 1781
rect 4506 1778 4726 1781
rect 4882 1778 5046 1781
rect 5050 1778 5118 1781
rect 402 1768 566 1771
rect 730 1768 798 1771
rect 1082 1768 1102 1771
rect 1106 1768 1113 1771
rect 1186 1768 1198 1771
rect 1202 1768 1206 1771
rect 1210 1768 1558 1771
rect 1570 1768 1726 1771
rect 1738 1768 1798 1771
rect 1818 1768 1974 1771
rect 2170 1768 2174 1771
rect 2202 1768 2206 1771
rect 2210 1768 2534 1771
rect 2538 1768 2606 1771
rect 2766 1771 2769 1778
rect 4278 1772 4281 1778
rect 2650 1768 2769 1771
rect 2834 1768 2846 1771
rect 2866 1768 2974 1771
rect 3186 1768 3990 1771
rect 4006 1768 4062 1771
rect 4090 1768 4110 1771
rect 4354 1768 4510 1771
rect 4578 1768 4726 1771
rect 4986 1768 4998 1771
rect 5074 1768 5166 1771
rect 378 1758 382 1761
rect 418 1758 422 1761
rect 546 1758 590 1761
rect 762 1758 910 1761
rect 1090 1758 1329 1761
rect 1434 1758 1510 1761
rect 1562 1758 1654 1761
rect 1714 1758 1718 1761
rect 1746 1758 1758 1761
rect 1762 1758 1990 1761
rect 2054 1761 2057 1768
rect 3038 1762 3041 1768
rect 4006 1762 4009 1768
rect 2018 1758 2057 1761
rect 2066 1758 2246 1761
rect 2410 1758 2422 1761
rect 2490 1758 2510 1761
rect 2514 1758 2606 1761
rect 2642 1758 2678 1761
rect 2730 1758 2782 1761
rect 2786 1758 2838 1761
rect 2866 1758 2934 1761
rect 3146 1758 3182 1761
rect 3322 1758 3374 1761
rect 3498 1758 3630 1761
rect 3698 1758 3838 1761
rect 3842 1758 4006 1761
rect 4050 1758 4142 1761
rect 4178 1758 4182 1761
rect 4226 1758 4246 1761
rect 4274 1758 4334 1761
rect 4410 1758 4454 1761
rect 4458 1758 4510 1761
rect 4546 1758 4614 1761
rect 4706 1758 4710 1761
rect 4866 1758 4966 1761
rect 5098 1758 5294 1761
rect 1326 1752 1329 1758
rect 290 1748 358 1751
rect 442 1748 518 1751
rect 586 1748 590 1751
rect 602 1748 734 1751
rect 738 1748 742 1751
rect 782 1748 790 1751
rect 794 1748 854 1751
rect 18 1738 70 1741
rect 142 1741 145 1748
rect 254 1741 257 1748
rect 978 1748 982 1751
rect 1026 1748 1097 1751
rect 1138 1748 1158 1751
rect 1274 1748 1318 1751
rect 1330 1748 1382 1751
rect 1426 1748 1430 1751
rect 1554 1748 1566 1751
rect 1658 1748 1710 1751
rect 1802 1748 1902 1751
rect 1922 1748 1966 1751
rect 1986 1748 2030 1751
rect 2138 1748 2534 1751
rect 2726 1751 2729 1758
rect 2602 1748 2729 1751
rect 2766 1748 2886 1751
rect 2990 1751 2993 1758
rect 2922 1748 2993 1751
rect 3010 1748 3046 1751
rect 3122 1748 3126 1751
rect 3130 1748 3262 1751
rect 3298 1748 3302 1751
rect 3306 1748 3326 1751
rect 3346 1748 3382 1751
rect 3386 1748 3438 1751
rect 3514 1748 3521 1751
rect 3546 1748 3550 1751
rect 3570 1748 3654 1751
rect 3830 1748 3838 1751
rect 3842 1748 3870 1751
rect 3906 1748 3942 1751
rect 4194 1748 4270 1751
rect 4290 1748 4550 1751
rect 4610 1748 4614 1751
rect 4690 1748 4702 1751
rect 4718 1751 4721 1758
rect 4734 1751 4737 1758
rect 4718 1748 4830 1751
rect 4850 1748 4862 1751
rect 5026 1748 5038 1751
rect 5078 1751 5081 1758
rect 5066 1748 5081 1751
rect 1094 1742 1097 1748
rect 1406 1742 1409 1748
rect 2766 1742 2769 1748
rect 142 1738 257 1741
rect 378 1738 414 1741
rect 442 1738 510 1741
rect 586 1738 726 1741
rect 754 1738 806 1741
rect 906 1738 934 1741
rect 1058 1738 1070 1741
rect 1146 1738 1150 1741
rect 1178 1738 1326 1741
rect 1330 1738 1334 1741
rect 1426 1738 1542 1741
rect 1578 1738 1582 1741
rect 1722 1738 1766 1741
rect 1794 1738 1830 1741
rect 1946 1738 1974 1741
rect 1978 1738 2142 1741
rect 2178 1738 2550 1741
rect 2586 1738 2630 1741
rect 2930 1738 2958 1741
rect 3062 1741 3065 1748
rect 3982 1742 3985 1748
rect 3062 1738 3086 1741
rect 3138 1738 3142 1741
rect 3178 1738 3238 1741
rect 3258 1738 3361 1741
rect 3394 1738 3534 1741
rect 3586 1738 3670 1741
rect 3754 1738 3838 1741
rect 3922 1738 3942 1741
rect 4066 1738 4134 1741
rect 4202 1738 4270 1741
rect 4282 1738 4502 1741
rect 4506 1738 4606 1741
rect 4670 1741 4673 1748
rect 4642 1738 4673 1741
rect 4802 1738 4846 1741
rect 4898 1738 4942 1741
rect 4946 1738 5094 1741
rect 5114 1738 5174 1741
rect 5214 1741 5217 1748
rect 5230 1741 5233 1748
rect 5214 1738 5233 1741
rect 66 1728 158 1731
rect 162 1728 238 1731
rect 562 1728 614 1731
rect 834 1728 990 1731
rect 1226 1728 1254 1731
rect 1322 1728 1374 1731
rect 1406 1728 1670 1731
rect 1678 1731 1681 1738
rect 1678 1728 1782 1731
rect 1786 1728 1934 1731
rect 1958 1728 2014 1731
rect 2042 1728 2062 1731
rect 2106 1728 2158 1731
rect 2218 1728 2358 1731
rect 2574 1731 2577 1738
rect 2450 1728 2577 1731
rect 2742 1731 2745 1738
rect 2742 1728 2806 1731
rect 2830 1731 2833 1738
rect 3358 1732 3361 1738
rect 2830 1728 3041 1731
rect 3050 1728 3110 1731
rect 3250 1728 3294 1731
rect 3298 1728 3342 1731
rect 3506 1728 3518 1731
rect 3546 1728 3606 1731
rect 3642 1728 3854 1731
rect 3858 1728 3894 1731
rect 4122 1728 4238 1731
rect 4306 1728 4462 1731
rect 4466 1728 4473 1731
rect 4658 1728 4710 1731
rect 4714 1728 4734 1731
rect 4738 1728 4814 1731
rect 4818 1728 4886 1731
rect 5058 1728 5086 1731
rect 162 1718 198 1721
rect 202 1718 398 1721
rect 770 1718 918 1721
rect 1406 1721 1409 1728
rect 1958 1722 1961 1728
rect 930 1718 1409 1721
rect 1418 1718 1430 1721
rect 1434 1718 1734 1721
rect 1826 1718 1830 1721
rect 1862 1718 1950 1721
rect 1970 1718 2174 1721
rect 2514 1718 2518 1721
rect 2546 1718 2590 1721
rect 2594 1718 2614 1721
rect 2794 1718 2982 1721
rect 2986 1718 2998 1721
rect 3038 1721 3041 1728
rect 3038 1718 3206 1721
rect 4170 1718 4198 1721
rect 4242 1718 4270 1721
rect 4314 1718 4318 1721
rect 4346 1718 4358 1721
rect 4378 1718 4390 1721
rect 4906 1718 5126 1721
rect 98 1708 134 1711
rect 138 1708 294 1711
rect 338 1708 390 1711
rect 394 1708 718 1711
rect 918 1711 921 1718
rect 918 1708 1406 1711
rect 1626 1708 1630 1711
rect 1862 1711 1865 1718
rect 3022 1712 3025 1718
rect 1690 1708 1865 1711
rect 2042 1708 2262 1711
rect 2522 1708 2526 1711
rect 2538 1708 2598 1711
rect 2618 1708 2670 1711
rect 3386 1708 3414 1711
rect 3418 1708 3902 1711
rect 4138 1708 4206 1711
rect 4978 1708 5030 1711
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 862 1703 864 1707
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1886 1703 1888 1707
rect 1958 1702 1961 1708
rect 2888 1703 2890 1707
rect 2894 1703 2897 1707
rect 2902 1703 2904 1707
rect 3920 1703 3922 1707
rect 3926 1703 3929 1707
rect 3934 1703 3936 1707
rect 4936 1703 4938 1707
rect 4942 1703 4945 1707
rect 4950 1703 4952 1707
rect 258 1698 438 1701
rect 482 1698 590 1701
rect 978 1698 1014 1701
rect 1122 1698 1414 1701
rect 1522 1698 1622 1701
rect 2042 1698 2046 1701
rect 2106 1698 2566 1701
rect 2818 1698 2870 1701
rect 3018 1698 3030 1701
rect 3042 1698 3102 1701
rect 3162 1698 3638 1701
rect 3658 1698 3870 1701
rect 3874 1698 3902 1701
rect 4042 1698 4166 1701
rect 4170 1698 4334 1701
rect 4338 1698 4358 1701
rect 4362 1698 4462 1701
rect 4466 1698 4518 1701
rect 4602 1698 4750 1701
rect 3150 1692 3153 1698
rect 122 1688 382 1691
rect 402 1688 558 1691
rect 754 1688 782 1691
rect 786 1688 894 1691
rect 1326 1688 1334 1691
rect 1338 1688 1710 1691
rect 1722 1688 1769 1691
rect 1810 1688 1926 1691
rect 1938 1688 1974 1691
rect 1994 1688 2049 1691
rect 2058 1688 2086 1691
rect 2098 1688 2182 1691
rect 2498 1688 2606 1691
rect 2610 1688 2654 1691
rect 2762 1688 2814 1691
rect 2830 1688 2910 1691
rect 2938 1688 3070 1691
rect 3074 1688 3118 1691
rect 3122 1688 3145 1691
rect 3170 1688 3222 1691
rect 3226 1688 3238 1691
rect 3306 1688 3358 1691
rect 3466 1688 3489 1691
rect 3554 1688 3614 1691
rect 3618 1688 3718 1691
rect 4026 1688 4070 1691
rect 4074 1688 4214 1691
rect 4234 1688 4254 1691
rect 4330 1688 4438 1691
rect 4666 1688 4718 1691
rect 4898 1688 5126 1691
rect 5202 1688 5206 1691
rect 5242 1688 5254 1691
rect 1766 1682 1769 1688
rect 2046 1682 2049 1688
rect 130 1678 166 1681
rect 170 1678 406 1681
rect 426 1678 518 1681
rect 522 1678 542 1681
rect 570 1678 646 1681
rect 650 1678 750 1681
rect 874 1678 950 1681
rect 1114 1678 1134 1681
rect 1202 1678 1302 1681
rect 1306 1678 1310 1681
rect 1370 1678 1406 1681
rect 1570 1678 1670 1681
rect 1730 1678 1750 1681
rect 1786 1678 1942 1681
rect 1946 1678 2038 1681
rect 2050 1678 2486 1681
rect 2694 1681 2697 1688
rect 2830 1682 2833 1688
rect 3142 1682 3145 1688
rect 3486 1682 3489 1688
rect 2694 1678 2750 1681
rect 2754 1678 2761 1681
rect 2850 1678 2854 1681
rect 2878 1678 2886 1681
rect 2890 1678 2998 1681
rect 3098 1678 3126 1681
rect 3146 1678 3470 1681
rect 3634 1678 3662 1681
rect 3802 1678 3854 1681
rect 3906 1678 4174 1681
rect 4226 1678 4774 1681
rect 4778 1678 4926 1681
rect 4970 1678 4974 1681
rect 5010 1678 5078 1681
rect 218 1668 454 1671
rect 570 1668 606 1671
rect 610 1668 638 1671
rect 642 1668 902 1671
rect 914 1668 918 1671
rect 922 1668 926 1671
rect 946 1668 1046 1671
rect 1082 1668 1110 1671
rect 1130 1668 1206 1671
rect 1282 1668 1326 1671
rect 1362 1668 1422 1671
rect 1466 1668 1494 1671
rect 1498 1668 1502 1671
rect 1578 1668 1582 1671
rect 1650 1668 1654 1671
rect 1690 1668 2118 1671
rect 2130 1668 2230 1671
rect 2370 1668 2390 1671
rect 2510 1671 2513 1678
rect 5238 1672 5241 1678
rect 2394 1668 2513 1671
rect 2538 1668 2598 1671
rect 2674 1668 2726 1671
rect 2810 1668 2878 1671
rect 2978 1668 3070 1671
rect 3082 1668 3086 1671
rect 3090 1668 3174 1671
rect 3218 1668 3222 1671
rect 3242 1668 3270 1671
rect 3274 1668 3334 1671
rect 3346 1668 3446 1671
rect 3450 1668 3558 1671
rect 3650 1668 3654 1671
rect 3714 1668 3742 1671
rect 3954 1668 4030 1671
rect 4098 1668 4158 1671
rect 4202 1668 4214 1671
rect 4290 1668 4318 1671
rect 4446 1668 4470 1671
rect 4490 1668 4678 1671
rect 4722 1668 4790 1671
rect 4862 1668 4918 1671
rect 5050 1668 5070 1671
rect 5074 1668 5166 1671
rect 5170 1668 5190 1671
rect 58 1658 102 1661
rect 162 1658 190 1661
rect 194 1658 217 1661
rect 226 1658 257 1661
rect 290 1658 350 1661
rect 354 1658 566 1661
rect 618 1658 646 1661
rect 754 1658 1126 1661
rect 1146 1658 1262 1661
rect 1266 1658 1390 1661
rect 1426 1658 1430 1661
rect 1514 1658 1569 1661
rect 1578 1659 1638 1661
rect 1574 1658 1638 1659
rect 1746 1658 1782 1661
rect 1786 1658 1902 1661
rect 1946 1658 2110 1661
rect 2118 1661 2121 1668
rect 2622 1662 2625 1668
rect 2118 1658 2182 1661
rect 2258 1658 2278 1661
rect 2282 1658 2294 1661
rect 2298 1658 2326 1661
rect 2330 1658 2342 1661
rect 2482 1658 2486 1661
rect 2642 1658 2646 1661
rect 2658 1658 2678 1661
rect 2682 1658 2686 1661
rect 2722 1658 2838 1661
rect 2858 1658 2902 1661
rect 3010 1658 3046 1661
rect 3050 1658 3078 1661
rect 3146 1658 3150 1661
rect 3218 1658 3334 1661
rect 3402 1658 3406 1661
rect 3426 1658 3446 1661
rect 3482 1658 3550 1661
rect 3650 1658 3654 1661
rect 3674 1658 3702 1661
rect 3750 1661 3753 1668
rect 3750 1658 3830 1661
rect 3946 1658 4014 1661
rect 4034 1658 4150 1661
rect 4154 1658 4158 1661
rect 4162 1658 4174 1661
rect 4202 1658 4206 1661
rect 4446 1661 4449 1668
rect 4862 1662 4865 1668
rect 5262 1662 5265 1668
rect 4258 1658 4449 1661
rect 4458 1658 4478 1661
rect 4498 1658 4502 1661
rect 4522 1658 4582 1661
rect 4690 1658 4694 1661
rect 4714 1658 4718 1661
rect 4746 1658 4774 1661
rect 4882 1658 4886 1661
rect 5050 1658 5086 1661
rect 5170 1658 5174 1661
rect 5178 1658 5185 1661
rect 5226 1658 5238 1661
rect 214 1652 217 1658
rect 254 1652 257 1658
rect 114 1648 142 1651
rect 314 1648 334 1651
rect 338 1648 374 1651
rect 442 1648 462 1651
rect 482 1648 582 1651
rect 586 1648 806 1651
rect 850 1648 1006 1651
rect 1010 1648 1310 1651
rect 1330 1648 1494 1651
rect 1498 1648 1534 1651
rect 1566 1651 1569 1658
rect 1566 1648 1622 1651
rect 1674 1648 1678 1651
rect 1710 1648 1718 1651
rect 1722 1648 1750 1651
rect 1762 1648 1814 1651
rect 1898 1648 1934 1651
rect 2010 1648 2014 1651
rect 2090 1648 2126 1651
rect 2470 1651 2473 1658
rect 3390 1652 3393 1658
rect 5182 1652 5185 1658
rect 2470 1648 2526 1651
rect 2650 1648 2758 1651
rect 2762 1648 3038 1651
rect 3106 1648 3110 1651
rect 3194 1648 3254 1651
rect 3258 1648 3270 1651
rect 3330 1648 3350 1651
rect 3354 1648 3374 1651
rect 3650 1648 3670 1651
rect 3770 1648 3830 1651
rect 3834 1648 3998 1651
rect 4002 1648 4030 1651
rect 4098 1648 4190 1651
rect 4274 1648 4334 1651
rect 4594 1648 4646 1651
rect 4762 1648 4822 1651
rect 4866 1648 5030 1651
rect 5066 1648 5126 1651
rect 2070 1642 2073 1648
rect 4238 1642 4241 1648
rect 130 1638 174 1641
rect 178 1638 182 1641
rect 210 1638 446 1641
rect 458 1638 550 1641
rect 554 1638 566 1641
rect 586 1638 590 1641
rect 594 1638 758 1641
rect 762 1638 878 1641
rect 882 1638 1702 1641
rect 1706 1638 1990 1641
rect 2090 1638 2118 1641
rect 2266 1638 2774 1641
rect 2818 1638 2958 1641
rect 3010 1638 3054 1641
rect 3154 1638 3198 1641
rect 3218 1638 3230 1641
rect 3682 1638 4086 1641
rect 4330 1638 4862 1641
rect 4866 1638 5038 1641
rect 578 1628 614 1631
rect 690 1628 766 1631
rect 818 1628 838 1631
rect 1058 1628 1630 1631
rect 1858 1628 1958 1631
rect 1962 1628 2214 1631
rect 2466 1628 2614 1631
rect 2622 1628 2630 1631
rect 2634 1628 2862 1631
rect 3098 1628 3230 1631
rect 3762 1628 3854 1631
rect 4206 1628 4630 1631
rect 4634 1628 4646 1631
rect 4658 1628 5062 1631
rect 194 1618 390 1621
rect 394 1618 398 1621
rect 410 1618 654 1621
rect 690 1618 1302 1621
rect 1306 1618 2142 1621
rect 2442 1618 2873 1621
rect 2882 1618 3310 1621
rect 3314 1618 3574 1621
rect 3578 1618 4062 1621
rect 4206 1621 4209 1628
rect 4066 1618 4209 1621
rect 4410 1618 4502 1621
rect 4962 1618 5030 1621
rect 5098 1618 5110 1621
rect 386 1608 430 1611
rect 650 1608 686 1611
rect 690 1608 798 1611
rect 962 1608 1278 1611
rect 1394 1608 1398 1611
rect 1490 1608 1526 1611
rect 1542 1608 1686 1611
rect 1698 1608 1734 1611
rect 1738 1608 1758 1611
rect 1818 1608 1950 1611
rect 2010 1608 2374 1611
rect 2426 1608 2654 1611
rect 2850 1608 2854 1611
rect 2870 1611 2873 1618
rect 2870 1608 2990 1611
rect 3146 1608 3366 1611
rect 3986 1608 4134 1611
rect 4146 1608 4286 1611
rect 4570 1608 5094 1611
rect 328 1603 330 1607
rect 334 1603 337 1607
rect 342 1603 344 1607
rect 1352 1603 1354 1607
rect 1358 1603 1361 1607
rect 1366 1603 1368 1607
rect 626 1598 694 1601
rect 702 1598 1054 1601
rect 1130 1598 1134 1601
rect 1542 1601 1545 1608
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2398 1603 2400 1607
rect 3400 1603 3402 1607
rect 3406 1603 3409 1607
rect 3414 1603 3416 1607
rect 4424 1603 4426 1607
rect 4430 1603 4433 1607
rect 4438 1603 4440 1607
rect 1410 1598 1545 1601
rect 1554 1598 1678 1601
rect 1682 1598 1726 1601
rect 1754 1598 1790 1601
rect 1802 1598 1894 1601
rect 1954 1598 2246 1601
rect 2274 1598 2278 1601
rect 2778 1598 2910 1601
rect 2930 1598 3014 1601
rect 3506 1598 4022 1601
rect 4042 1598 4230 1601
rect 4706 1598 4902 1601
rect 702 1592 705 1598
rect 314 1588 702 1591
rect 1026 1588 1182 1591
rect 1186 1588 1854 1591
rect 1906 1588 2022 1591
rect 2114 1588 2166 1591
rect 2234 1588 2454 1591
rect 2458 1588 2470 1591
rect 2610 1588 2750 1591
rect 2754 1588 2790 1591
rect 2906 1588 3030 1591
rect 3034 1588 3118 1591
rect 3122 1588 3622 1591
rect 3778 1588 3846 1591
rect 3850 1588 4166 1591
rect 4226 1588 4278 1591
rect 4466 1588 4582 1591
rect 274 1578 318 1581
rect 410 1578 422 1581
rect 522 1578 598 1581
rect 610 1578 638 1581
rect 1018 1578 1086 1581
rect 1402 1578 1566 1581
rect 1714 1578 1718 1581
rect 1818 1578 1942 1581
rect 1986 1578 2350 1581
rect 2402 1578 2462 1581
rect 2586 1578 2630 1581
rect 2878 1581 2881 1588
rect 2878 1578 2942 1581
rect 3026 1578 3078 1581
rect 3386 1578 3782 1581
rect 3786 1578 3846 1581
rect 3850 1578 4030 1581
rect 4194 1578 4262 1581
rect 4266 1578 4454 1581
rect 4458 1578 4494 1581
rect 4498 1578 4614 1581
rect 4674 1578 4702 1581
rect 4994 1578 5022 1581
rect 106 1568 134 1571
rect 402 1568 670 1571
rect 674 1568 710 1571
rect 1050 1568 1054 1571
rect 1134 1571 1137 1578
rect 1166 1571 1169 1578
rect 1134 1568 1169 1571
rect 1346 1568 1454 1571
rect 1498 1568 1558 1571
rect 1666 1568 1718 1571
rect 1834 1568 1918 1571
rect 2502 1571 2505 1578
rect 1922 1568 2505 1571
rect 2570 1568 2678 1571
rect 2826 1568 2846 1571
rect 2850 1568 2934 1571
rect 2958 1571 2961 1578
rect 2958 1568 3022 1571
rect 3026 1568 3046 1571
rect 3110 1571 3113 1578
rect 3074 1568 3113 1571
rect 3226 1568 3366 1571
rect 3378 1568 3422 1571
rect 3834 1568 3838 1571
rect 3858 1568 3886 1571
rect 3906 1568 3910 1571
rect 4234 1568 4238 1571
rect 4258 1568 4294 1571
rect 4314 1568 4334 1571
rect 4402 1568 4438 1571
rect 4658 1568 4662 1571
rect 4690 1568 4702 1571
rect 4706 1568 4766 1571
rect 4770 1568 4878 1571
rect 4882 1568 4886 1571
rect 4930 1568 5054 1571
rect 5146 1568 5262 1571
rect 146 1558 166 1561
rect 254 1561 257 1568
rect 1118 1562 1121 1568
rect 1462 1562 1465 1568
rect 250 1558 257 1561
rect 386 1558 678 1561
rect 1322 1558 1358 1561
rect 1362 1558 1406 1561
rect 1418 1558 1422 1561
rect 1482 1558 1486 1561
rect 1506 1558 1510 1561
rect 1574 1561 1577 1568
rect 1574 1558 1622 1561
rect 1650 1558 1718 1561
rect 1734 1561 1737 1568
rect 1734 1558 1742 1561
rect 1782 1561 1785 1568
rect 4102 1562 4105 1568
rect 1778 1558 1785 1561
rect 1866 1558 1966 1561
rect 1994 1558 1998 1561
rect 2034 1558 2054 1561
rect 2114 1558 2230 1561
rect 2290 1558 2358 1561
rect 2422 1558 2446 1561
rect 2594 1558 3254 1561
rect 3282 1558 3478 1561
rect 3570 1558 3646 1561
rect 3698 1558 3734 1561
rect 3866 1558 4070 1561
rect 4174 1561 4177 1568
rect 4566 1562 4569 1568
rect 4598 1562 4601 1568
rect 4162 1558 4177 1561
rect 4250 1558 4470 1561
rect 4474 1558 4534 1561
rect 4586 1558 4590 1561
rect 4622 1558 4630 1561
rect 4686 1561 4689 1568
rect 4650 1558 4689 1561
rect 4698 1558 4702 1561
rect 4706 1558 4830 1561
rect 106 1548 126 1551
rect 154 1548 214 1551
rect 250 1548 278 1551
rect 374 1551 377 1558
rect 338 1548 406 1551
rect 418 1548 470 1551
rect 562 1548 590 1551
rect 626 1548 630 1551
rect 646 1542 649 1548
rect 654 1542 657 1548
rect 662 1542 665 1551
rect 674 1548 734 1551
rect 738 1548 758 1551
rect 810 1548 814 1551
rect 914 1548 990 1551
rect 1018 1548 1022 1551
rect 1082 1548 1094 1551
rect 1170 1548 1174 1551
rect 1290 1548 1342 1551
rect 1346 1548 1582 1551
rect 1586 1548 1638 1551
rect 1730 1548 1974 1551
rect 2002 1548 2038 1551
rect 2138 1548 2174 1551
rect 2422 1551 2425 1558
rect 3542 1552 3545 1558
rect 2346 1548 2425 1551
rect 2434 1548 2646 1551
rect 2786 1548 2854 1551
rect 2922 1548 2926 1551
rect 2938 1548 2950 1551
rect 2986 1548 3086 1551
rect 3090 1548 3126 1551
rect 3242 1548 3270 1551
rect 3346 1548 3350 1551
rect 3682 1548 3790 1551
rect 3838 1551 3841 1558
rect 3818 1548 3841 1551
rect 3882 1548 3886 1551
rect 3906 1548 4158 1551
rect 4162 1548 4302 1551
rect 4542 1551 4545 1558
rect 4622 1552 4625 1558
rect 4338 1548 4545 1551
rect 4570 1548 4598 1551
rect 1742 1542 1745 1548
rect 3846 1542 3849 1548
rect 4318 1542 4321 1548
rect 4762 1548 4817 1551
rect 4838 1551 4841 1558
rect 4826 1548 4841 1551
rect 4858 1548 4862 1551
rect 4882 1548 4894 1551
rect 5034 1548 5038 1551
rect 5066 1548 5070 1551
rect 5090 1548 5134 1551
rect 5154 1548 5241 1551
rect 4814 1542 4817 1548
rect 42 1538 110 1541
rect 122 1538 142 1541
rect 146 1538 454 1541
rect 458 1538 526 1541
rect 586 1538 590 1541
rect 754 1538 982 1541
rect 986 1538 1014 1541
rect 1122 1538 1126 1541
rect 1162 1538 1166 1541
rect 1250 1538 1326 1541
rect 1466 1538 1470 1541
rect 1530 1538 1534 1541
rect 1546 1538 1558 1541
rect 1562 1538 1662 1541
rect 1770 1538 1838 1541
rect 1930 1538 1934 1541
rect 1978 1538 1990 1541
rect 2010 1538 2030 1541
rect 2050 1538 2254 1541
rect 2322 1538 2486 1541
rect 2498 1538 2545 1541
rect 2578 1538 2713 1541
rect 2794 1538 2798 1541
rect 2818 1538 2974 1541
rect 2994 1538 3078 1541
rect 3098 1538 3102 1541
rect 3122 1538 3150 1541
rect 3258 1538 3262 1541
rect 3266 1538 3286 1541
rect 3306 1538 3350 1541
rect 3490 1538 3494 1541
rect 3530 1538 3590 1541
rect 3626 1538 3630 1541
rect 3634 1538 3670 1541
rect 3698 1538 3702 1541
rect 3706 1538 3718 1541
rect 3986 1538 4046 1541
rect 4106 1538 4110 1541
rect 4146 1538 4150 1541
rect 4170 1538 4190 1541
rect 4210 1538 4238 1541
rect 4250 1538 4286 1541
rect 4378 1538 4382 1541
rect 4402 1538 4406 1541
rect 4442 1538 4494 1541
rect 4498 1538 4806 1541
rect 4850 1538 4886 1541
rect 5014 1541 5017 1548
rect 5238 1542 5241 1548
rect 5014 1538 5150 1541
rect 218 1528 222 1531
rect 346 1528 366 1531
rect 370 1528 438 1531
rect 482 1528 558 1531
rect 658 1528 878 1531
rect 922 1528 1150 1531
rect 1298 1528 1430 1531
rect 1494 1531 1497 1538
rect 2542 1532 2545 1538
rect 2614 1532 2617 1538
rect 2710 1532 2713 1538
rect 3086 1532 3089 1538
rect 1458 1528 1497 1531
rect 1522 1528 1718 1531
rect 1770 1528 1774 1531
rect 1850 1528 1862 1531
rect 1898 1528 1966 1531
rect 2002 1528 2006 1531
rect 2042 1528 2118 1531
rect 2146 1528 2406 1531
rect 2466 1528 2518 1531
rect 2790 1528 2822 1531
rect 2874 1528 2902 1531
rect 2934 1528 2990 1531
rect 3034 1528 3070 1531
rect 3302 1531 3305 1538
rect 3266 1528 3305 1531
rect 3346 1528 3430 1531
rect 3578 1528 3606 1531
rect 3754 1528 3822 1531
rect 3826 1528 3966 1531
rect 4226 1528 4638 1531
rect 4642 1528 4798 1531
rect 4802 1528 5006 1531
rect 5050 1528 5078 1531
rect 174 1521 177 1528
rect 174 1518 390 1521
rect 586 1518 590 1521
rect 602 1518 1142 1521
rect 1146 1518 1582 1521
rect 1586 1518 1726 1521
rect 1734 1521 1737 1528
rect 2790 1522 2793 1528
rect 2934 1522 2937 1528
rect 1734 1518 1993 1521
rect 2050 1518 2078 1521
rect 2090 1518 2134 1521
rect 2186 1518 2286 1521
rect 2434 1518 2518 1521
rect 2522 1518 2574 1521
rect 2578 1518 2598 1521
rect 2714 1518 2726 1521
rect 2746 1518 2790 1521
rect 3018 1518 3046 1521
rect 3234 1518 3273 1521
rect 3534 1521 3537 1528
rect 5238 1522 5241 1528
rect 3394 1518 3537 1521
rect 3650 1518 3694 1521
rect 3698 1518 3902 1521
rect 4066 1518 4102 1521
rect 4114 1518 4206 1521
rect 4234 1518 4462 1521
rect 4466 1518 4718 1521
rect 4866 1518 4974 1521
rect 122 1508 342 1511
rect 370 1508 582 1511
rect 1106 1508 1542 1511
rect 1546 1508 1766 1511
rect 1770 1508 1782 1511
rect 1906 1508 1942 1511
rect 1990 1511 1993 1518
rect 3270 1512 3273 1518
rect 1990 1508 2150 1511
rect 2266 1508 2318 1511
rect 2322 1508 2486 1511
rect 2490 1508 2550 1511
rect 2554 1508 2574 1511
rect 2658 1508 2814 1511
rect 2914 1508 2934 1511
rect 2938 1508 3006 1511
rect 3018 1508 3062 1511
rect 3082 1508 3190 1511
rect 3330 1508 3486 1511
rect 3490 1508 3558 1511
rect 4090 1508 4102 1511
rect 4106 1508 4222 1511
rect 4266 1508 4270 1511
rect 4362 1508 4366 1511
rect 4410 1508 4470 1511
rect 4498 1508 4502 1511
rect 4562 1508 4606 1511
rect 4634 1508 4694 1511
rect 5154 1508 5206 1511
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 862 1503 864 1507
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1886 1503 1888 1507
rect 1958 1502 1961 1508
rect 2888 1503 2890 1507
rect 2894 1503 2897 1507
rect 2902 1503 2904 1507
rect 3920 1503 3922 1507
rect 3926 1503 3929 1507
rect 3934 1503 3936 1507
rect 4622 1502 4625 1508
rect 4936 1503 4938 1507
rect 4942 1503 4945 1507
rect 4950 1503 4952 1507
rect 130 1498 214 1501
rect 242 1498 326 1501
rect 354 1498 710 1501
rect 754 1498 814 1501
rect 1218 1498 1494 1501
rect 1498 1498 1638 1501
rect 1706 1498 1750 1501
rect 1762 1498 1862 1501
rect 1922 1498 1926 1501
rect 2050 1498 2054 1501
rect 2058 1498 2062 1501
rect 2202 1498 2238 1501
rect 2250 1498 2806 1501
rect 2994 1498 3022 1501
rect 3034 1498 3038 1501
rect 3114 1498 3150 1501
rect 3154 1498 3206 1501
rect 3258 1498 3286 1501
rect 3298 1498 3382 1501
rect 3474 1498 3526 1501
rect 3530 1498 3638 1501
rect 4034 1498 4174 1501
rect 4242 1498 4270 1501
rect 4274 1498 4318 1501
rect 4386 1498 4566 1501
rect 4578 1498 4614 1501
rect 306 1488 310 1491
rect 322 1488 382 1491
rect 386 1488 462 1491
rect 566 1488 654 1491
rect 682 1488 830 1491
rect 850 1488 990 1491
rect 1314 1488 1334 1491
rect 1482 1488 1566 1491
rect 1590 1488 1598 1491
rect 1602 1488 1678 1491
rect 1698 1488 1702 1491
rect 1710 1488 1737 1491
rect 1762 1488 1966 1491
rect 1970 1488 2102 1491
rect 2130 1488 2233 1491
rect 2242 1488 2278 1491
rect 2282 1488 2430 1491
rect 2434 1488 2446 1491
rect 2698 1488 3310 1491
rect 3434 1488 3486 1491
rect 3658 1488 3974 1491
rect 4050 1488 4350 1491
rect 4386 1488 4590 1491
rect 4594 1488 4734 1491
rect 4762 1488 4790 1491
rect 4842 1488 4902 1491
rect 4906 1488 4950 1491
rect 5058 1488 5062 1491
rect 566 1482 569 1488
rect 98 1478 134 1481
rect 138 1478 166 1481
rect 378 1478 414 1481
rect 450 1478 454 1481
rect 778 1478 894 1481
rect 1710 1481 1713 1488
rect 1098 1478 1713 1481
rect 1734 1481 1737 1488
rect 1734 1478 1790 1481
rect 1794 1478 1822 1481
rect 1858 1478 2134 1481
rect 2178 1478 2222 1481
rect 2230 1481 2233 1488
rect 2590 1482 2593 1488
rect 2230 1478 2246 1481
rect 2458 1478 2462 1481
rect 2706 1478 2726 1481
rect 2730 1478 2998 1481
rect 3002 1478 3262 1481
rect 3282 1478 3286 1481
rect 3306 1478 3638 1481
rect 3642 1478 3662 1481
rect 3666 1478 3790 1481
rect 3794 1478 3854 1481
rect 3858 1478 3870 1481
rect 3874 1478 3894 1481
rect 3914 1478 3982 1481
rect 3986 1478 4054 1481
rect 4146 1478 4217 1481
rect 4250 1478 4278 1481
rect 4354 1478 4390 1481
rect 4410 1478 4481 1481
rect 4530 1478 4766 1481
rect 4818 1478 4894 1481
rect 5058 1478 5182 1481
rect 302 1472 305 1478
rect 614 1472 617 1478
rect 1726 1472 1729 1478
rect 106 1468 145 1471
rect 202 1468 230 1471
rect 738 1468 790 1471
rect 794 1468 798 1471
rect 922 1468 926 1471
rect 1050 1468 1105 1471
rect 142 1462 145 1468
rect 390 1462 393 1468
rect 870 1462 873 1468
rect 1102 1462 1105 1468
rect 1338 1468 1374 1471
rect 1570 1468 1574 1471
rect 1634 1468 1638 1471
rect 1682 1468 1694 1471
rect 1738 1468 1742 1471
rect 1754 1468 1758 1471
rect 1778 1468 1782 1471
rect 1802 1468 1926 1471
rect 1930 1468 1934 1471
rect 1954 1468 1974 1471
rect 2018 1468 2062 1471
rect 2066 1468 2078 1471
rect 2122 1468 2214 1471
rect 2270 1471 2273 1478
rect 2310 1471 2313 1478
rect 2218 1468 2494 1471
rect 2530 1468 2542 1471
rect 2562 1468 2654 1471
rect 2998 1468 3390 1471
rect 3482 1468 3510 1471
rect 3514 1468 3646 1471
rect 3650 1468 3654 1471
rect 3874 1468 3982 1471
rect 3986 1468 4078 1471
rect 4098 1468 4166 1471
rect 4170 1468 4177 1471
rect 4186 1468 4190 1471
rect 4214 1471 4217 1478
rect 4478 1472 4481 1478
rect 5190 1472 5193 1478
rect 4214 1468 4270 1471
rect 4314 1468 4318 1471
rect 4402 1468 4462 1471
rect 4490 1468 4494 1471
rect 4562 1468 4654 1471
rect 4810 1468 4822 1471
rect 4930 1468 4934 1471
rect 5198 1471 5201 1478
rect 5198 1468 5246 1471
rect 58 1458 113 1461
rect 162 1458 190 1461
rect 194 1458 230 1461
rect 234 1458 246 1461
rect 354 1458 358 1461
rect 394 1458 446 1461
rect 506 1458 510 1461
rect 618 1458 622 1461
rect 794 1458 846 1461
rect 986 1458 1070 1461
rect 1114 1458 1118 1461
rect 1170 1458 1174 1461
rect 1246 1461 1249 1468
rect 1246 1458 1254 1461
rect 1270 1461 1273 1468
rect 1502 1462 1505 1468
rect 1266 1458 1273 1461
rect 1282 1458 1334 1461
rect 1354 1458 1390 1461
rect 1454 1458 1486 1461
rect 1550 1461 1553 1468
rect 2542 1462 2545 1468
rect 1550 1458 1822 1461
rect 1826 1458 1846 1461
rect 1890 1458 1894 1461
rect 1906 1458 1910 1461
rect 1922 1458 1942 1461
rect 1946 1458 1990 1461
rect 1994 1458 2054 1461
rect 2154 1458 2230 1461
rect 2306 1458 2390 1461
rect 2434 1458 2454 1461
rect 2554 1459 2598 1461
rect 2694 1461 2697 1468
rect 2554 1458 2601 1459
rect 2694 1458 2750 1461
rect 2754 1458 2758 1461
rect 2778 1458 2886 1461
rect 2950 1461 2953 1468
rect 2950 1458 2966 1461
rect 2998 1461 3001 1468
rect 2970 1458 3001 1461
rect 3074 1458 3110 1461
rect 3122 1458 3350 1461
rect 3354 1458 3470 1461
rect 3474 1458 3630 1461
rect 3650 1458 3654 1461
rect 3970 1458 4030 1461
rect 4122 1458 4158 1461
rect 4174 1461 4177 1468
rect 4174 1458 4190 1461
rect 4206 1461 4209 1468
rect 4782 1462 4785 1468
rect 4206 1458 4270 1461
rect 4282 1458 4342 1461
rect 4474 1458 4486 1461
rect 4626 1458 4694 1461
rect 4810 1458 4814 1461
rect 4846 1458 4918 1461
rect 4922 1458 4929 1461
rect 4938 1458 5006 1461
rect 5102 1461 5105 1468
rect 5066 1458 5105 1461
rect 5122 1458 5150 1461
rect 5170 1458 5174 1461
rect 5186 1458 5198 1461
rect 5202 1458 5222 1461
rect 110 1452 113 1458
rect 1446 1452 1449 1458
rect 1454 1452 1457 1458
rect 178 1448 406 1451
rect 418 1448 430 1451
rect 442 1448 582 1451
rect 1010 1448 1142 1451
rect 1146 1448 1222 1451
rect 1242 1448 1254 1451
rect 1258 1448 1262 1451
rect 1282 1448 1294 1451
rect 1370 1448 1446 1451
rect 1562 1448 1654 1451
rect 1698 1448 1702 1451
rect 1722 1448 1734 1451
rect 1918 1451 1921 1458
rect 1738 1448 1921 1451
rect 1946 1448 2022 1451
rect 2078 1448 2105 1451
rect 2130 1448 2222 1451
rect 2298 1448 2326 1451
rect 2430 1451 2433 1458
rect 2346 1448 2433 1451
rect 2462 1452 2465 1458
rect 2514 1448 2598 1451
rect 2602 1448 2862 1451
rect 2898 1448 2942 1451
rect 2946 1448 3014 1451
rect 3018 1448 3102 1451
rect 3106 1448 3166 1451
rect 3170 1448 3390 1451
rect 3442 1448 3542 1451
rect 3586 1448 3614 1451
rect 3622 1448 3678 1451
rect 3794 1448 3806 1451
rect 3850 1448 3854 1451
rect 3858 1448 4398 1451
rect 4454 1451 4457 1458
rect 4846 1452 4849 1458
rect 4454 1448 4550 1451
rect 4890 1448 4990 1451
rect 4994 1448 5134 1451
rect 2078 1442 2081 1448
rect 2102 1442 2105 1448
rect 3622 1442 3625 1448
rect 178 1438 246 1441
rect 250 1438 334 1441
rect 354 1438 366 1441
rect 698 1438 838 1441
rect 1018 1438 1054 1441
rect 1058 1438 1078 1441
rect 1082 1438 1214 1441
rect 1258 1438 1734 1441
rect 1738 1438 1782 1441
rect 1794 1438 1854 1441
rect 1906 1438 1966 1441
rect 2010 1438 2014 1441
rect 2138 1438 2438 1441
rect 2770 1438 2806 1441
rect 2866 1438 2878 1441
rect 2994 1438 2998 1441
rect 3002 1438 3102 1441
rect 3114 1438 3134 1441
rect 3314 1438 3366 1441
rect 3678 1441 3681 1448
rect 3678 1438 3790 1441
rect 3890 1438 3958 1441
rect 4162 1438 4182 1441
rect 4218 1438 4878 1441
rect 4882 1438 5110 1441
rect 5114 1438 5126 1441
rect 5202 1438 5206 1441
rect 586 1428 774 1431
rect 886 1431 889 1438
rect 4054 1432 4057 1438
rect 778 1428 889 1431
rect 1130 1428 1302 1431
rect 1334 1428 1342 1431
rect 1346 1428 1374 1431
rect 1394 1428 1430 1431
rect 1442 1428 1558 1431
rect 1570 1428 1574 1431
rect 1594 1428 1830 1431
rect 1834 1428 2070 1431
rect 2218 1428 2238 1431
rect 2250 1428 2286 1431
rect 2290 1428 2446 1431
rect 2450 1428 2582 1431
rect 2882 1428 3078 1431
rect 3362 1428 3438 1431
rect 3442 1428 3566 1431
rect 3594 1428 3686 1431
rect 3842 1428 3958 1431
rect 4202 1428 4798 1431
rect 4906 1428 4966 1431
rect 5034 1428 5078 1431
rect 430 1421 433 1428
rect 430 1418 590 1421
rect 786 1418 806 1421
rect 842 1418 1022 1421
rect 1138 1418 1182 1421
rect 1186 1418 1982 1421
rect 2130 1418 2158 1421
rect 2162 1418 2246 1421
rect 2258 1418 2302 1421
rect 2434 1418 2686 1421
rect 2690 1418 2766 1421
rect 2930 1418 3854 1421
rect 4066 1418 4430 1421
rect 4434 1418 4558 1421
rect 4578 1418 4670 1421
rect 4746 1418 4750 1421
rect 4778 1418 4790 1421
rect 4818 1418 5158 1421
rect 1030 1412 1033 1418
rect 434 1408 478 1411
rect 1082 1408 1222 1411
rect 1234 1408 1318 1411
rect 1466 1408 1526 1411
rect 1530 1408 1838 1411
rect 1962 1408 1974 1411
rect 2274 1408 2350 1411
rect 2506 1408 2878 1411
rect 2978 1408 3222 1411
rect 3522 1408 3798 1411
rect 3826 1408 4014 1411
rect 4050 1408 4326 1411
rect 4458 1408 4702 1411
rect 4914 1408 4998 1411
rect 5042 1408 5070 1411
rect 328 1403 330 1407
rect 334 1403 337 1407
rect 342 1403 344 1407
rect 1352 1403 1354 1407
rect 1358 1403 1361 1407
rect 1366 1403 1368 1407
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2398 1403 2400 1407
rect 3400 1403 3402 1407
rect 3406 1403 3409 1407
rect 3414 1403 3416 1407
rect 4382 1402 4385 1408
rect 4424 1403 4426 1407
rect 4430 1403 4433 1407
rect 4438 1403 4440 1407
rect 410 1398 654 1401
rect 658 1398 1102 1401
rect 1538 1398 1894 1401
rect 2226 1398 2286 1401
rect 2298 1398 2310 1401
rect 2466 1398 2470 1401
rect 2546 1398 2550 1401
rect 2674 1398 2761 1401
rect 2770 1398 2958 1401
rect 3130 1398 3214 1401
rect 3218 1398 3366 1401
rect 3530 1398 3766 1401
rect 3946 1398 4150 1401
rect 4282 1398 4374 1401
rect 4546 1398 4638 1401
rect 4918 1398 5046 1401
rect 5050 1398 5206 1401
rect 474 1388 486 1391
rect 658 1388 1030 1391
rect 1110 1388 1118 1391
rect 1122 1388 1150 1391
rect 1162 1388 1166 1391
rect 1322 1388 1342 1391
rect 1402 1388 1422 1391
rect 1434 1388 1486 1391
rect 1514 1388 1630 1391
rect 1634 1388 1774 1391
rect 1826 1388 2454 1391
rect 2542 1388 2742 1391
rect 2758 1391 2761 1398
rect 4918 1392 4921 1398
rect 2758 1388 3086 1391
rect 3090 1388 3118 1391
rect 3178 1388 3390 1391
rect 3746 1388 3822 1391
rect 4258 1388 4494 1391
rect 4722 1388 4750 1391
rect 4754 1388 4918 1391
rect 2542 1382 2545 1388
rect 458 1378 502 1381
rect 762 1378 790 1381
rect 970 1378 990 1381
rect 994 1378 1174 1381
rect 1346 1378 1374 1381
rect 1378 1378 2198 1381
rect 2522 1378 2542 1381
rect 2578 1378 2590 1381
rect 2874 1378 3070 1381
rect 3082 1378 3326 1381
rect 3330 1378 3502 1381
rect 3546 1378 3598 1381
rect 3754 1378 3966 1381
rect 3970 1378 4078 1381
rect 4306 1378 4438 1381
rect 4506 1378 4510 1381
rect 4518 1378 4686 1381
rect 4778 1378 4830 1381
rect 4834 1378 4950 1381
rect 5062 1381 5065 1388
rect 4970 1378 5065 1381
rect 2214 1372 2217 1378
rect 178 1368 1014 1371
rect 1038 1368 1086 1371
rect 1122 1368 2014 1371
rect 2098 1368 2166 1371
rect 2178 1368 2198 1371
rect 2242 1368 2342 1371
rect 2498 1368 2558 1371
rect 2566 1371 2569 1378
rect 2566 1368 2614 1371
rect 2726 1368 2950 1371
rect 2954 1368 2958 1371
rect 2978 1368 3054 1371
rect 3394 1368 3398 1371
rect 3754 1368 3790 1371
rect 4010 1368 4118 1371
rect 4246 1371 4249 1378
rect 4518 1372 4521 1378
rect 4246 1368 4502 1371
rect 4890 1368 4934 1371
rect 5058 1368 5102 1371
rect 206 1362 209 1368
rect 1038 1362 1041 1368
rect 226 1358 278 1361
rect 314 1358 526 1361
rect 562 1358 766 1361
rect 818 1358 1014 1361
rect 1050 1358 1134 1361
rect 1146 1358 1198 1361
rect 1210 1358 1462 1361
rect 1466 1358 1582 1361
rect 1610 1358 1622 1361
rect 1866 1358 1958 1361
rect 2014 1361 2017 1368
rect 1986 1358 2017 1361
rect 2146 1358 2198 1361
rect 2202 1358 2238 1361
rect 2254 1358 2262 1361
rect 2266 1358 2318 1361
rect 2330 1358 2433 1361
rect 2482 1358 2518 1361
rect 2526 1358 2534 1361
rect 2726 1361 2729 1368
rect 2538 1358 2729 1361
rect 3158 1361 3161 1368
rect 3154 1358 3161 1361
rect 3174 1361 3177 1368
rect 3294 1362 3297 1368
rect 3174 1358 3270 1361
rect 3354 1358 3358 1361
rect 3378 1358 3406 1361
rect 3426 1358 3454 1361
rect 3602 1358 3638 1361
rect 3682 1358 3774 1361
rect 4226 1358 4278 1361
rect 4314 1358 4390 1361
rect 4418 1358 4422 1361
rect 4474 1358 4478 1361
rect 4514 1358 4518 1361
rect 4578 1358 4582 1361
rect 4598 1361 4601 1368
rect 4598 1358 4606 1361
rect 4618 1358 4622 1361
rect 4810 1358 4814 1361
rect 4858 1358 5046 1361
rect 5130 1358 5182 1361
rect 5302 1361 5305 1368
rect 5186 1358 5305 1361
rect 110 1351 113 1358
rect 110 1348 198 1351
rect 266 1348 270 1351
rect 378 1348 390 1351
rect 418 1348 494 1351
rect 522 1348 526 1351
rect 622 1348 670 1351
rect 706 1348 758 1351
rect 786 1348 942 1351
rect 946 1348 974 1351
rect 1170 1348 1214 1351
rect 1226 1348 1470 1351
rect 1474 1348 1582 1351
rect 1686 1351 1689 1358
rect 1586 1348 1681 1351
rect 1686 1348 1694 1351
rect 1798 1351 1801 1358
rect 2046 1352 2049 1358
rect 1794 1348 1801 1351
rect 1962 1348 2014 1351
rect 2034 1348 2038 1351
rect 2098 1348 2422 1351
rect 2430 1351 2433 1358
rect 2526 1352 2529 1358
rect 2798 1352 2801 1358
rect 3054 1352 3057 1358
rect 2430 1348 2510 1351
rect 2514 1348 2521 1351
rect 2554 1348 2558 1351
rect 2578 1348 2582 1351
rect 2618 1348 2673 1351
rect 2706 1348 2734 1351
rect 3002 1348 3006 1351
rect 3138 1348 3158 1351
rect 3162 1348 3606 1351
rect 3654 1351 3657 1358
rect 3634 1348 3657 1351
rect 3666 1348 3734 1351
rect 3770 1348 4014 1351
rect 4214 1351 4217 1358
rect 4718 1352 4721 1358
rect 4766 1352 4769 1358
rect 4106 1348 4217 1351
rect 4226 1348 4230 1351
rect 4274 1348 4374 1351
rect 4386 1348 4590 1351
rect 4618 1348 4630 1351
rect 4634 1348 4678 1351
rect 4762 1348 4766 1351
rect 4770 1348 5022 1351
rect 5030 1348 5038 1351
rect 5062 1351 5065 1358
rect 5094 1352 5097 1358
rect 5042 1348 5065 1351
rect 5074 1348 5086 1351
rect 5146 1348 5166 1351
rect 5186 1348 5246 1351
rect 130 1338 166 1341
rect 242 1338 246 1341
rect 266 1338 278 1341
rect 282 1338 318 1341
rect 398 1341 401 1348
rect 414 1341 417 1348
rect 622 1342 625 1348
rect 1054 1342 1057 1348
rect 398 1338 417 1341
rect 426 1338 534 1341
rect 722 1338 849 1341
rect 874 1338 950 1341
rect 1018 1338 1038 1341
rect 1066 1338 1238 1341
rect 1306 1338 1422 1341
rect 1522 1338 1566 1341
rect 1602 1338 1606 1341
rect 1618 1338 1638 1341
rect 1642 1338 1654 1341
rect 1678 1341 1681 1348
rect 1702 1341 1705 1348
rect 1678 1338 1705 1341
rect 1718 1342 1721 1348
rect 1782 1342 1785 1348
rect 1878 1341 1881 1348
rect 2670 1342 2673 1348
rect 2966 1342 2969 1348
rect 1858 1338 1881 1341
rect 1986 1338 1998 1341
rect 2026 1338 2190 1341
rect 2226 1338 2230 1341
rect 2290 1338 2334 1341
rect 2410 1338 2414 1341
rect 2506 1338 2577 1341
rect 3042 1338 3062 1341
rect 3146 1338 3206 1341
rect 3274 1338 3334 1341
rect 3362 1338 3366 1341
rect 3378 1338 3502 1341
rect 3802 1338 3902 1341
rect 4058 1338 4062 1341
rect 4098 1338 4134 1341
rect 4314 1338 4406 1341
rect 4410 1338 4454 1341
rect 4498 1338 4542 1341
rect 4610 1338 4622 1341
rect 4650 1338 4654 1341
rect 4706 1338 4734 1341
rect 4762 1338 4774 1341
rect 4922 1338 4926 1341
rect 4930 1338 4942 1341
rect 5010 1338 5030 1341
rect 5050 1338 5094 1341
rect 5106 1338 5142 1341
rect 5186 1338 5198 1341
rect 846 1332 849 1338
rect 1246 1332 1249 1338
rect 74 1328 478 1331
rect 482 1328 510 1331
rect 530 1328 558 1331
rect 562 1328 774 1331
rect 1042 1328 1118 1331
rect 1290 1328 1302 1331
rect 1518 1331 1521 1338
rect 1966 1332 1969 1338
rect 2262 1332 2265 1338
rect 1306 1328 1521 1331
rect 1530 1328 1582 1331
rect 1650 1328 1654 1331
rect 1706 1328 1942 1331
rect 1946 1328 1958 1331
rect 2026 1328 2030 1331
rect 2266 1328 2310 1331
rect 2338 1328 2342 1331
rect 2410 1328 2462 1331
rect 2546 1328 2558 1331
rect 2574 1331 2577 1338
rect 2726 1331 2729 1338
rect 3558 1332 3561 1338
rect 3582 1332 3585 1338
rect 2574 1328 2729 1331
rect 2738 1328 2894 1331
rect 2898 1328 2905 1331
rect 2994 1328 3302 1331
rect 3322 1328 3438 1331
rect 3678 1331 3681 1338
rect 3678 1328 3718 1331
rect 3746 1328 3910 1331
rect 4098 1328 4206 1331
rect 4282 1328 4286 1331
rect 4670 1331 4673 1338
rect 4290 1328 4673 1331
rect 4986 1328 5222 1331
rect 2326 1322 2329 1328
rect 4742 1322 4745 1328
rect 18 1318 86 1321
rect 218 1318 238 1321
rect 778 1318 790 1321
rect 978 1318 1062 1321
rect 1338 1318 1350 1321
rect 1354 1318 1614 1321
rect 1746 1318 1822 1321
rect 1842 1318 1998 1321
rect 2450 1318 2462 1321
rect 2498 1318 2582 1321
rect 2586 1318 2614 1321
rect 2642 1318 2782 1321
rect 2922 1318 3150 1321
rect 3234 1318 3238 1321
rect 3298 1318 3302 1321
rect 3594 1318 3814 1321
rect 3858 1318 4254 1321
rect 4274 1318 4326 1321
rect 4482 1318 4574 1321
rect 4930 1318 5030 1321
rect 5038 1318 5046 1321
rect 5050 1318 5086 1321
rect 5122 1318 5206 1321
rect 130 1308 526 1311
rect 930 1308 974 1311
rect 986 1308 1070 1311
rect 1074 1308 1270 1311
rect 1314 1308 1406 1311
rect 1418 1308 1558 1311
rect 1590 1308 1606 1311
rect 1762 1308 1838 1311
rect 2018 1308 2110 1311
rect 2114 1308 2182 1311
rect 2186 1308 2286 1311
rect 2290 1308 2486 1311
rect 2506 1308 2870 1311
rect 3074 1308 3158 1311
rect 3162 1308 3694 1311
rect 3698 1308 3766 1311
rect 3810 1308 3814 1311
rect 3826 1308 3854 1311
rect 3978 1308 4246 1311
rect 4250 1308 4326 1311
rect 4394 1308 4774 1311
rect 5018 1308 5094 1311
rect 5114 1308 5126 1311
rect 5202 1308 5214 1311
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 862 1303 864 1307
rect 186 1298 238 1301
rect 242 1298 246 1301
rect 250 1298 750 1301
rect 798 1298 841 1301
rect 986 1298 1062 1301
rect 1074 1298 1198 1301
rect 1590 1301 1593 1308
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1886 1303 1888 1307
rect 2888 1303 2890 1307
rect 2894 1303 2897 1307
rect 2902 1303 2904 1307
rect 3920 1303 3922 1307
rect 3926 1303 3929 1307
rect 3934 1303 3936 1307
rect 4936 1303 4938 1307
rect 4942 1303 4945 1307
rect 4950 1303 4952 1307
rect 1394 1298 1593 1301
rect 1602 1298 1614 1301
rect 1682 1298 1718 1301
rect 1722 1298 1838 1301
rect 1986 1298 2070 1301
rect 2074 1298 2150 1301
rect 2314 1298 2398 1301
rect 2410 1298 2734 1301
rect 3082 1298 3102 1301
rect 3106 1298 3126 1301
rect 3138 1298 3286 1301
rect 3290 1298 3430 1301
rect 3594 1298 3606 1301
rect 3842 1298 3910 1301
rect 3994 1298 4398 1301
rect 4450 1298 4542 1301
rect 5082 1298 5150 1301
rect 798 1292 801 1298
rect 154 1288 182 1291
rect 458 1288 486 1291
rect 738 1288 798 1291
rect 838 1291 841 1298
rect 1382 1292 1385 1298
rect 1862 1292 1865 1298
rect 3830 1292 3833 1298
rect 838 1288 870 1291
rect 882 1288 1166 1291
rect 1430 1288 1814 1291
rect 1874 1288 1974 1291
rect 1978 1288 2014 1291
rect 2050 1288 2334 1291
rect 2450 1288 2502 1291
rect 2530 1288 2774 1291
rect 2794 1288 2862 1291
rect 2866 1288 2966 1291
rect 2970 1288 3118 1291
rect 3186 1288 3238 1291
rect 3322 1288 3342 1291
rect 3462 1288 3758 1291
rect 3906 1288 4070 1291
rect 4074 1288 4190 1291
rect 4194 1288 4310 1291
rect 4330 1288 4470 1291
rect 4626 1288 4766 1291
rect 4770 1288 4854 1291
rect 4962 1288 5006 1291
rect 5074 1288 5113 1291
rect 182 1281 185 1288
rect 182 1278 222 1281
rect 234 1278 462 1281
rect 466 1278 614 1281
rect 706 1278 774 1281
rect 806 1281 809 1288
rect 1430 1282 1433 1288
rect 1526 1282 1529 1288
rect 3462 1282 3465 1288
rect 3782 1282 3785 1288
rect 794 1278 809 1281
rect 834 1278 870 1281
rect 954 1278 990 1281
rect 1050 1278 1358 1281
rect 1362 1278 1390 1281
rect 1642 1278 1710 1281
rect 1714 1278 1734 1281
rect 1838 1278 1926 1281
rect 1946 1278 1982 1281
rect 2066 1278 2190 1281
rect 2194 1278 2238 1281
rect 2242 1278 2406 1281
rect 2426 1278 2446 1281
rect 2450 1278 2702 1281
rect 2778 1278 2798 1281
rect 2962 1278 3358 1281
rect 3482 1278 3502 1281
rect 3806 1281 3809 1288
rect 5110 1282 5113 1288
rect 3806 1278 3870 1281
rect 3890 1278 3990 1281
rect 4266 1278 4270 1281
rect 4290 1278 4350 1281
rect 4378 1278 4510 1281
rect 4570 1278 4574 1281
rect 4818 1278 4990 1281
rect 4994 1278 5102 1281
rect 42 1268 110 1271
rect 130 1268 134 1271
rect 290 1268 422 1271
rect 442 1268 446 1271
rect 602 1268 665 1271
rect 754 1268 822 1271
rect 866 1268 886 1271
rect 906 1268 942 1271
rect 954 1268 958 1271
rect 970 1268 974 1271
rect 1010 1268 1014 1271
rect 1098 1268 1302 1271
rect 1406 1271 1409 1278
rect 1838 1272 1841 1278
rect 3510 1272 3513 1278
rect 1386 1268 1409 1271
rect 1650 1268 1825 1271
rect 1914 1268 2486 1271
rect 2490 1268 2694 1271
rect 2802 1268 2814 1271
rect 2834 1268 2854 1271
rect 2858 1268 3150 1271
rect 3154 1268 3214 1271
rect 3386 1268 3470 1271
rect 3622 1271 3625 1278
rect 3546 1268 3625 1271
rect 3762 1268 3822 1271
rect 3850 1268 3974 1271
rect 4034 1268 4046 1271
rect 4178 1268 4246 1271
rect 4250 1268 4257 1271
rect 4266 1268 4294 1271
rect 4330 1268 4334 1271
rect 4346 1268 4390 1271
rect 4410 1268 4510 1271
rect 4514 1268 4694 1271
rect 4826 1268 4870 1271
rect 4906 1268 4982 1271
rect 5058 1268 5126 1271
rect 5190 1268 5246 1271
rect 106 1258 126 1261
rect 210 1258 230 1261
rect 270 1261 273 1268
rect 662 1262 665 1268
rect 838 1262 841 1268
rect 270 1258 286 1261
rect 290 1258 406 1261
rect 426 1258 430 1261
rect 762 1258 774 1261
rect 810 1258 814 1261
rect 842 1258 1006 1261
rect 1086 1261 1089 1268
rect 1086 1259 1142 1261
rect 1086 1258 1145 1259
rect 1170 1258 1214 1261
rect 1318 1261 1321 1268
rect 1250 1258 1321 1261
rect 1414 1261 1417 1268
rect 1402 1258 1417 1261
rect 1478 1261 1481 1268
rect 1822 1262 1825 1268
rect 2982 1262 2985 1268
rect 3222 1262 3225 1268
rect 3246 1262 3249 1268
rect 3278 1262 3281 1268
rect 5190 1262 5193 1268
rect 1458 1258 1481 1261
rect 1530 1258 1558 1261
rect 1562 1258 1654 1261
rect 1674 1258 1678 1261
rect 1690 1258 1766 1261
rect 2018 1258 2033 1261
rect 2042 1258 2134 1261
rect 2138 1258 2302 1261
rect 2386 1258 2406 1261
rect 2482 1258 2486 1261
rect 2522 1258 2526 1261
rect 2546 1258 2550 1261
rect 2554 1258 2561 1261
rect 2570 1258 2646 1261
rect 2722 1258 2734 1261
rect 2762 1258 2766 1261
rect 2786 1258 2854 1261
rect 2874 1258 2910 1261
rect 2946 1258 2950 1261
rect 3002 1258 3006 1261
rect 3082 1258 3086 1261
rect 3098 1258 3158 1261
rect 3334 1258 3342 1261
rect 3562 1258 3598 1261
rect 3730 1258 3742 1261
rect 3746 1258 3758 1261
rect 3762 1258 3846 1261
rect 3850 1258 3862 1261
rect 3918 1258 4078 1261
rect 4082 1258 4102 1261
rect 4114 1258 4126 1261
rect 4130 1258 4326 1261
rect 4338 1258 4366 1261
rect 4538 1258 4606 1261
rect 4690 1258 4718 1261
rect 4722 1258 4862 1261
rect 4866 1258 4894 1261
rect 5002 1258 5182 1261
rect 98 1248 142 1251
rect 146 1248 190 1251
rect 254 1251 257 1258
rect 1838 1252 1841 1258
rect 254 1248 374 1251
rect 642 1248 662 1251
rect 906 1248 1190 1251
rect 1298 1248 1342 1251
rect 1346 1248 1358 1251
rect 1378 1248 1430 1251
rect 1474 1248 1478 1251
rect 1570 1248 1574 1251
rect 1618 1248 1726 1251
rect 1922 1248 1934 1251
rect 1962 1248 2022 1251
rect 2030 1251 2033 1258
rect 2454 1252 2457 1258
rect 3294 1252 3297 1258
rect 3334 1252 3337 1258
rect 3918 1252 3921 1258
rect 4398 1252 4401 1258
rect 4446 1252 4449 1258
rect 5094 1252 5097 1258
rect 2030 1248 2070 1251
rect 2106 1248 2150 1251
rect 2178 1248 2254 1251
rect 2482 1248 2598 1251
rect 2690 1248 2710 1251
rect 2722 1248 2926 1251
rect 2946 1248 3054 1251
rect 3058 1248 3270 1251
rect 3714 1248 3918 1251
rect 3946 1248 4174 1251
rect 4178 1248 4294 1251
rect 4338 1248 4342 1251
rect 4386 1248 4390 1251
rect 4546 1248 4590 1251
rect 4914 1248 4918 1251
rect 4938 1248 5054 1251
rect 170 1238 278 1241
rect 282 1238 310 1241
rect 314 1238 550 1241
rect 554 1238 1446 1241
rect 1450 1238 1606 1241
rect 1730 1238 1958 1241
rect 2010 1238 2025 1241
rect 2270 1241 2273 1248
rect 2242 1238 2273 1241
rect 2302 1242 2305 1248
rect 2326 1241 2329 1248
rect 2326 1238 2342 1241
rect 2346 1238 2774 1241
rect 2954 1238 3262 1241
rect 3274 1238 3561 1241
rect 3730 1238 3734 1241
rect 3746 1238 3766 1241
rect 3882 1238 4022 1241
rect 4426 1238 4654 1241
rect 2022 1232 2025 1238
rect 578 1228 638 1231
rect 650 1228 1118 1231
rect 1354 1228 1414 1231
rect 1490 1228 2017 1231
rect 2330 1228 3078 1231
rect 3098 1228 3550 1231
rect 3558 1231 3561 1238
rect 3558 1228 3766 1231
rect 3794 1228 3846 1231
rect 3850 1228 3894 1231
rect 3978 1228 4750 1231
rect 5090 1228 5174 1231
rect 158 1222 161 1228
rect 746 1218 886 1221
rect 890 1218 902 1221
rect 954 1218 958 1221
rect 994 1218 1054 1221
rect 1066 1218 1990 1221
rect 2014 1221 2017 1228
rect 2014 1218 2102 1221
rect 2202 1218 2342 1221
rect 2554 1218 2566 1221
rect 2626 1218 2878 1221
rect 3034 1218 3150 1221
rect 3298 1218 3390 1221
rect 3394 1218 3494 1221
rect 3514 1218 3926 1221
rect 3930 1218 3990 1221
rect 4662 1218 4686 1221
rect 4898 1218 5102 1221
rect 5106 1218 5158 1221
rect 2958 1212 2961 1218
rect 4662 1212 4665 1218
rect 842 1208 926 1211
rect 962 1208 982 1211
rect 1018 1208 1174 1211
rect 1410 1208 1486 1211
rect 1490 1208 1894 1211
rect 1986 1208 2262 1211
rect 2450 1208 2462 1211
rect 2786 1208 2838 1211
rect 2842 1208 2878 1211
rect 3018 1208 3030 1211
rect 3074 1208 3150 1211
rect 3218 1208 3310 1211
rect 3330 1208 3366 1211
rect 4290 1208 4414 1211
rect 5106 1208 5118 1211
rect 328 1203 330 1207
rect 334 1203 337 1207
rect 342 1203 344 1207
rect 1352 1203 1354 1207
rect 1358 1203 1361 1207
rect 1366 1203 1368 1207
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2398 1203 2400 1207
rect 3400 1203 3402 1207
rect 3406 1203 3409 1207
rect 3414 1203 3416 1207
rect 4424 1203 4426 1207
rect 4430 1203 4433 1207
rect 4438 1203 4440 1207
rect 834 1198 1094 1201
rect 1378 1198 1398 1201
rect 1402 1198 1550 1201
rect 1866 1198 1894 1201
rect 1898 1198 1950 1201
rect 2426 1198 2478 1201
rect 2674 1198 2921 1201
rect 2930 1198 3182 1201
rect 3234 1198 3238 1201
rect 3242 1198 3374 1201
rect 3530 1198 3566 1201
rect 3818 1198 4302 1201
rect 4458 1198 4646 1201
rect 4650 1198 4734 1201
rect 4738 1198 4902 1201
rect 4906 1198 5086 1201
rect 5090 1198 5150 1201
rect 1310 1192 1313 1198
rect 882 1188 886 1191
rect 890 1188 1102 1191
rect 1330 1188 1414 1191
rect 1466 1188 1558 1191
rect 1562 1188 1606 1191
rect 1610 1188 2046 1191
rect 2050 1188 2070 1191
rect 2082 1188 2326 1191
rect 2378 1188 2494 1191
rect 2498 1188 2542 1191
rect 2546 1188 2670 1191
rect 2674 1188 2870 1191
rect 2918 1191 2921 1198
rect 2918 1188 3070 1191
rect 3374 1191 3377 1198
rect 3374 1188 3430 1191
rect 3434 1188 3542 1191
rect 3658 1188 3686 1191
rect 3690 1188 3726 1191
rect 3786 1188 4214 1191
rect 4330 1188 4630 1191
rect 4674 1188 4998 1191
rect 5234 1188 5286 1191
rect 162 1178 214 1181
rect 218 1178 222 1181
rect 330 1178 606 1181
rect 1162 1178 1598 1181
rect 1698 1178 1854 1181
rect 2034 1178 2582 1181
rect 2594 1178 2598 1181
rect 2602 1178 2838 1181
rect 3126 1181 3129 1188
rect 2850 1178 3129 1181
rect 3234 1178 3246 1181
rect 3554 1178 3558 1181
rect 3634 1178 4326 1181
rect 4466 1178 4550 1181
rect 4638 1181 4641 1188
rect 4638 1178 4662 1181
rect 5218 1178 5262 1181
rect 150 1171 153 1178
rect 106 1168 153 1171
rect 230 1171 233 1178
rect 194 1168 233 1171
rect 818 1168 830 1171
rect 918 1171 921 1178
rect 906 1168 921 1171
rect 962 1168 1022 1171
rect 1122 1168 1222 1171
rect 1226 1168 1350 1171
rect 2090 1168 2182 1171
rect 2274 1168 2278 1171
rect 2554 1168 2574 1171
rect 2730 1168 2766 1171
rect 2770 1168 2830 1171
rect 3034 1168 3046 1171
rect 3050 1168 3606 1171
rect 3754 1168 3814 1171
rect 3962 1168 4070 1171
rect 4074 1168 4166 1171
rect 4250 1168 4382 1171
rect 4410 1168 4670 1171
rect 4886 1171 4889 1178
rect 4786 1168 4873 1171
rect 4886 1168 4902 1171
rect 5170 1168 5198 1171
rect 94 1161 97 1168
rect 94 1158 126 1161
rect 130 1158 166 1161
rect 182 1161 185 1168
rect 182 1158 270 1161
rect 410 1158 414 1161
rect 438 1161 441 1168
rect 434 1158 441 1161
rect 454 1161 457 1168
rect 454 1158 494 1161
rect 570 1158 606 1161
rect 610 1158 670 1161
rect 722 1158 726 1161
rect 898 1158 910 1161
rect 914 1158 1046 1161
rect 1094 1161 1097 1168
rect 1094 1158 1150 1161
rect 1218 1158 1222 1161
rect 1290 1158 1318 1161
rect 1338 1158 1406 1161
rect 1410 1158 1438 1161
rect 1454 1161 1457 1168
rect 1454 1158 1494 1161
rect 1822 1161 1825 1168
rect 1822 1158 2094 1161
rect 2114 1158 2302 1161
rect 2306 1158 2318 1161
rect 2454 1161 2457 1168
rect 4870 1162 4873 1168
rect 2370 1158 2457 1161
rect 2482 1158 2486 1161
rect 2570 1158 2862 1161
rect 2946 1158 2985 1161
rect 2994 1158 3022 1161
rect 3082 1158 3102 1161
rect 3114 1158 3278 1161
rect 3314 1158 3318 1161
rect 3378 1158 3414 1161
rect 3482 1158 3518 1161
rect 3546 1158 3550 1161
rect 3570 1158 3574 1161
rect 3634 1158 3638 1161
rect 3810 1158 3838 1161
rect 4042 1158 4182 1161
rect 4362 1158 4678 1161
rect 4986 1158 5046 1161
rect 5118 1161 5121 1168
rect 5134 1161 5137 1168
rect 5118 1158 5137 1161
rect 822 1152 825 1158
rect 58 1148 94 1151
rect 130 1148 198 1151
rect 202 1148 278 1151
rect 282 1148 390 1151
rect 410 1148 574 1151
rect 642 1148 646 1151
rect 722 1148 726 1151
rect 810 1148 814 1151
rect 842 1148 846 1151
rect 930 1148 934 1151
rect 938 1148 990 1151
rect 1070 1151 1073 1158
rect 1026 1148 1302 1151
rect 1306 1148 1334 1151
rect 1378 1148 1390 1151
rect 1394 1148 1406 1151
rect 1434 1148 1470 1151
rect 1530 1148 1534 1151
rect 1594 1148 1606 1151
rect 1610 1148 1614 1151
rect 1654 1151 1657 1158
rect 2566 1152 2569 1158
rect 2982 1152 2985 1158
rect 3350 1152 3353 1158
rect 3358 1152 3361 1158
rect 4006 1152 4009 1158
rect 4022 1152 4025 1158
rect 1634 1148 1657 1151
rect 1682 1148 1766 1151
rect 1770 1148 1846 1151
rect 1850 1148 1878 1151
rect 1882 1148 2046 1151
rect 2066 1148 2198 1151
rect 2226 1148 2238 1151
rect 2242 1148 2254 1151
rect 2274 1148 2366 1151
rect 2418 1148 2470 1151
rect 2474 1148 2518 1151
rect 2586 1148 2598 1151
rect 2730 1148 2734 1151
rect 2810 1148 2846 1151
rect 2850 1148 2958 1151
rect 2998 1148 3006 1151
rect 3010 1148 3022 1151
rect 3170 1148 3254 1151
rect 3266 1148 3270 1151
rect 3290 1148 3334 1151
rect 3410 1148 3574 1151
rect 3602 1148 3710 1151
rect 3770 1148 3774 1151
rect 3786 1148 3966 1151
rect 4138 1148 4142 1151
rect 4162 1148 4166 1151
rect 4370 1148 4390 1151
rect 4546 1148 4550 1151
rect 4594 1148 4622 1151
rect 4674 1148 4678 1151
rect 4742 1151 4745 1158
rect 4738 1148 4745 1151
rect 4830 1151 4833 1158
rect 4894 1151 4897 1158
rect 4830 1148 4897 1151
rect 4918 1151 4921 1158
rect 5166 1152 5169 1158
rect 5190 1152 5193 1158
rect 4914 1148 4921 1151
rect 4970 1148 5041 1151
rect 5058 1148 5110 1151
rect 5114 1148 5118 1151
rect 5274 1148 5286 1151
rect 130 1138 134 1141
rect 138 1138 150 1141
rect 158 1138 230 1141
rect 234 1138 262 1141
rect 306 1138 422 1141
rect 498 1138 694 1141
rect 722 1138 758 1141
rect 762 1138 1070 1141
rect 1074 1138 1102 1141
rect 1226 1138 2014 1141
rect 2018 1138 2142 1141
rect 2450 1138 2454 1141
rect 2458 1138 2606 1141
rect 2658 1138 2742 1141
rect 2826 1138 2894 1141
rect 2914 1138 2918 1141
rect 2958 1141 2961 1148
rect 3134 1142 3137 1148
rect 2958 1138 3014 1141
rect 3026 1138 3046 1141
rect 3162 1138 3182 1141
rect 3186 1138 3310 1141
rect 3362 1138 3374 1141
rect 3506 1138 3510 1141
rect 3578 1138 3598 1141
rect 4134 1141 4137 1148
rect 3610 1138 4137 1141
rect 4294 1142 4297 1148
rect 5038 1142 5041 1148
rect 4330 1138 4398 1141
rect 4474 1138 4558 1141
rect 4570 1138 4582 1141
rect 4602 1138 4638 1141
rect 4650 1138 4654 1141
rect 4898 1138 4918 1141
rect 4938 1138 4982 1141
rect 4986 1138 4990 1141
rect 5058 1138 5110 1141
rect 5122 1138 5134 1141
rect 5210 1138 5254 1141
rect 158 1132 161 1138
rect 2174 1132 2177 1138
rect 5150 1132 5153 1138
rect 402 1128 406 1131
rect 514 1128 582 1131
rect 694 1128 782 1131
rect 794 1128 814 1131
rect 818 1128 886 1131
rect 954 1128 998 1131
rect 1010 1128 1166 1131
rect 1274 1128 1654 1131
rect 1658 1128 1662 1131
rect 1666 1128 1814 1131
rect 2154 1128 2166 1131
rect 2290 1128 2718 1131
rect 2794 1128 2806 1131
rect 2818 1128 2846 1131
rect 2850 1128 3174 1131
rect 3178 1128 3238 1131
rect 3266 1128 3270 1131
rect 3362 1128 3502 1131
rect 3506 1128 3958 1131
rect 4090 1128 4254 1131
rect 4354 1128 4358 1131
rect 4586 1128 4590 1131
rect 4746 1128 4750 1131
rect 4898 1128 5126 1131
rect 694 1122 697 1128
rect 82 1118 214 1121
rect 266 1118 430 1121
rect 458 1118 574 1121
rect 706 1118 1062 1121
rect 1298 1118 1438 1121
rect 1554 1118 1630 1121
rect 1786 1118 1822 1121
rect 1826 1118 1934 1121
rect 1938 1118 2038 1121
rect 2042 1118 2078 1121
rect 2246 1121 2249 1128
rect 3326 1122 3329 1128
rect 3334 1122 3337 1128
rect 4654 1122 4657 1128
rect 2122 1118 2249 1121
rect 2618 1118 2862 1121
rect 2986 1118 3022 1121
rect 3034 1118 3086 1121
rect 3138 1118 3150 1121
rect 3290 1118 3310 1121
rect 3562 1118 3606 1121
rect 3626 1118 3654 1121
rect 3730 1118 3806 1121
rect 3826 1118 3934 1121
rect 4018 1118 4022 1121
rect 4026 1118 4030 1121
rect 4122 1118 4190 1121
rect 4282 1118 4350 1121
rect 4362 1118 4366 1121
rect 4418 1118 4454 1121
rect 4530 1118 4614 1121
rect 4698 1118 4886 1121
rect 4890 1118 4934 1121
rect 4954 1118 4966 1121
rect 4970 1118 5009 1121
rect 1294 1112 1297 1118
rect 2870 1112 2873 1118
rect 2950 1112 2953 1118
rect 5006 1112 5009 1118
rect 306 1108 702 1111
rect 706 1108 830 1111
rect 1258 1108 1278 1111
rect 1762 1108 1766 1111
rect 1898 1108 2134 1111
rect 2162 1108 2334 1111
rect 3098 1108 3158 1111
rect 3210 1108 3230 1111
rect 3306 1108 3454 1111
rect 3746 1108 3854 1111
rect 4042 1108 4078 1111
rect 4114 1108 4174 1111
rect 4754 1108 4766 1111
rect 5090 1108 5094 1111
rect 182 1102 185 1108
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 862 1103 864 1107
rect 1838 1102 1841 1108
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1886 1103 1888 1107
rect 2888 1103 2890 1107
rect 2894 1103 2897 1107
rect 2902 1103 2904 1107
rect 3920 1103 3922 1107
rect 3926 1103 3929 1107
rect 3934 1103 3936 1107
rect 4936 1103 4938 1107
rect 4942 1103 4945 1107
rect 4950 1103 4952 1107
rect 274 1098 302 1101
rect 562 1098 766 1101
rect 778 1098 798 1101
rect 1090 1098 1182 1101
rect 1218 1098 1518 1101
rect 1746 1098 1758 1101
rect 2050 1098 2166 1101
rect 2170 1098 2198 1101
rect 2202 1098 2214 1101
rect 2274 1098 2342 1101
rect 2386 1098 2502 1101
rect 2778 1098 2870 1101
rect 2922 1098 3334 1101
rect 3370 1098 3374 1101
rect 3442 1098 3494 1101
rect 3962 1098 4086 1101
rect 4402 1098 4606 1101
rect 4610 1098 4638 1101
rect 4666 1098 4758 1101
rect 5018 1098 5102 1101
rect 154 1088 334 1091
rect 374 1091 377 1098
rect 346 1088 377 1091
rect 602 1088 646 1091
rect 650 1088 686 1091
rect 802 1088 1454 1091
rect 1474 1088 1478 1091
rect 1642 1088 1798 1091
rect 2010 1088 2094 1091
rect 2330 1088 2446 1091
rect 2666 1088 2686 1091
rect 2690 1088 2798 1091
rect 2890 1088 2966 1091
rect 3154 1088 3270 1091
rect 3274 1088 3366 1091
rect 3490 1088 3566 1091
rect 3634 1088 3662 1091
rect 3722 1088 3806 1091
rect 3962 1088 4126 1091
rect 4210 1088 4238 1091
rect 4258 1088 4286 1091
rect 4290 1088 4326 1091
rect 4354 1088 4462 1091
rect 4490 1088 4590 1091
rect 4626 1088 4670 1091
rect 4714 1088 4758 1091
rect 4778 1088 4846 1091
rect 4850 1088 4910 1091
rect 5162 1088 5166 1091
rect 42 1078 118 1081
rect 130 1078 142 1081
rect 162 1078 174 1081
rect 442 1078 486 1081
rect 526 1081 529 1088
rect 3070 1082 3073 1088
rect 490 1078 529 1081
rect 678 1078 750 1081
rect 970 1078 990 1081
rect 994 1078 998 1081
rect 1010 1078 1038 1081
rect 1066 1078 1070 1081
rect 1306 1078 1366 1081
rect 1690 1078 1798 1081
rect 2146 1078 2422 1081
rect 2430 1078 2518 1081
rect 2530 1078 2558 1081
rect 2578 1078 2646 1081
rect 2714 1078 2774 1081
rect 2786 1078 2814 1081
rect 3138 1078 3262 1081
rect 3334 1078 3534 1081
rect 3594 1078 3630 1081
rect 3650 1078 3758 1081
rect 3762 1078 3774 1081
rect 3810 1078 3902 1081
rect 4058 1078 4574 1081
rect 4578 1078 4678 1081
rect 4682 1078 4894 1081
rect 4898 1078 4926 1081
rect 4930 1078 5094 1081
rect 66 1068 177 1071
rect 294 1071 297 1078
rect 678 1072 681 1078
rect 266 1068 297 1071
rect 418 1068 430 1071
rect 618 1068 630 1071
rect 690 1068 814 1071
rect 1102 1071 1105 1078
rect 2430 1072 2433 1078
rect 882 1068 1105 1071
rect 1226 1068 1318 1071
rect 1386 1068 1422 1071
rect 1458 1068 1505 1071
rect 1530 1068 1606 1071
rect 1722 1068 1734 1071
rect 1962 1068 1990 1071
rect 2002 1068 2334 1071
rect 2574 1071 2577 1078
rect 2498 1068 2577 1071
rect 2658 1068 2662 1071
rect 2730 1068 2734 1071
rect 2754 1068 2878 1071
rect 3134 1071 3137 1078
rect 3302 1072 3305 1078
rect 3334 1072 3337 1078
rect 5158 1072 5161 1078
rect 3042 1068 3137 1071
rect 3218 1068 3246 1071
rect 3626 1068 3670 1071
rect 3690 1068 3710 1071
rect 3714 1068 3721 1071
rect 3754 1068 3758 1071
rect 3986 1068 3990 1071
rect 4178 1068 4182 1071
rect 4242 1068 4262 1071
rect 4306 1068 4369 1071
rect 174 1062 177 1068
rect 114 1058 142 1061
rect 226 1058 262 1061
rect 546 1058 622 1061
rect 830 1061 833 1068
rect 1502 1062 1505 1068
rect 1854 1062 1857 1068
rect 2686 1062 2689 1068
rect 2718 1062 2721 1068
rect 830 1058 910 1061
rect 1018 1058 1022 1061
rect 1050 1058 1070 1061
rect 1258 1058 1294 1061
rect 1618 1058 1630 1061
rect 1650 1058 1734 1061
rect 1754 1058 1806 1061
rect 1914 1058 1942 1061
rect 1946 1058 1966 1061
rect 1970 1058 1990 1061
rect 2274 1058 2350 1061
rect 2418 1058 2534 1061
rect 2538 1058 2574 1061
rect 2610 1058 2678 1061
rect 2730 1058 2782 1061
rect 2786 1058 2910 1061
rect 2914 1058 2934 1061
rect 3026 1058 3086 1061
rect 3206 1061 3209 1068
rect 3254 1061 3257 1068
rect 3350 1062 3353 1068
rect 3206 1058 3257 1061
rect 3266 1058 3294 1061
rect 3330 1058 3342 1061
rect 3430 1061 3433 1068
rect 3394 1058 3433 1061
rect 3534 1062 3537 1068
rect 3546 1058 3638 1061
rect 3682 1058 3710 1061
rect 3770 1058 3774 1061
rect 3810 1058 3822 1061
rect 3870 1061 3873 1068
rect 3998 1062 4001 1068
rect 4046 1062 4049 1068
rect 3870 1058 3918 1061
rect 4018 1058 4046 1061
rect 4094 1061 4097 1068
rect 4366 1062 4369 1068
rect 4538 1068 4542 1071
rect 4638 1068 4710 1071
rect 4738 1068 4910 1071
rect 5082 1068 5134 1071
rect 5202 1068 5246 1071
rect 4094 1058 4110 1061
rect 4170 1058 4198 1061
rect 4234 1058 4238 1061
rect 4374 1061 4377 1068
rect 4630 1062 4633 1068
rect 4638 1062 4641 1068
rect 4374 1058 4382 1061
rect 4386 1058 4414 1061
rect 4418 1058 4566 1061
rect 4726 1061 4729 1068
rect 4726 1058 4798 1061
rect 4874 1058 4886 1061
rect 5166 1061 5169 1068
rect 5066 1058 5169 1061
rect 374 1051 377 1058
rect 298 1048 377 1051
rect 578 1048 598 1051
rect 602 1048 654 1051
rect 666 1048 838 1051
rect 1034 1048 1190 1051
rect 1254 1051 1257 1058
rect 1194 1048 1257 1051
rect 1298 1048 1310 1051
rect 1390 1051 1393 1058
rect 1390 1048 1430 1051
rect 1890 1048 1926 1051
rect 1982 1048 2038 1051
rect 2122 1048 2150 1051
rect 2218 1048 2382 1051
rect 2426 1048 2462 1051
rect 2562 1048 3526 1051
rect 3546 1048 3550 1051
rect 3642 1048 3646 1051
rect 3930 1048 3958 1051
rect 4154 1048 4166 1051
rect 4178 1048 4182 1051
rect 4338 1048 4390 1051
rect 4402 1048 4406 1051
rect 4530 1048 4534 1051
rect 4566 1051 4569 1058
rect 4566 1048 4582 1051
rect 4630 1051 4633 1058
rect 4630 1048 4830 1051
rect 4882 1048 4974 1051
rect 5122 1048 5134 1051
rect 1982 1042 1985 1048
rect 322 1038 358 1041
rect 802 1038 966 1041
rect 1002 1038 1238 1041
rect 1262 1038 1270 1041
rect 1274 1038 1406 1041
rect 1434 1038 1710 1041
rect 2130 1038 2142 1041
rect 2330 1038 2358 1041
rect 2674 1038 2734 1041
rect 2778 1038 3214 1041
rect 3498 1038 3822 1041
rect 4134 1041 4137 1048
rect 3826 1038 4137 1041
rect 4146 1038 4150 1041
rect 4182 1041 4185 1048
rect 4182 1038 4614 1041
rect 4634 1038 4646 1041
rect 4786 1038 4862 1041
rect 5114 1038 5198 1041
rect 226 1028 550 1031
rect 818 1028 950 1031
rect 1050 1028 1118 1031
rect 1194 1028 1206 1031
rect 1282 1028 2550 1031
rect 2610 1028 2734 1031
rect 2842 1028 2942 1031
rect 2970 1028 3006 1031
rect 3010 1028 3022 1031
rect 3242 1028 3462 1031
rect 3514 1028 4246 1031
rect 4250 1028 4310 1031
rect 4394 1028 4486 1031
rect 4682 1028 4838 1031
rect 210 1018 326 1021
rect 842 1018 846 1021
rect 922 1018 1054 1021
rect 1058 1018 2126 1021
rect 2810 1018 2966 1021
rect 2994 1018 3198 1021
rect 3238 1021 3241 1028
rect 3202 1018 3241 1021
rect 3322 1018 3590 1021
rect 3746 1018 3886 1021
rect 3906 1018 4054 1021
rect 4114 1018 4246 1021
rect 4266 1018 5190 1021
rect 5274 1018 5278 1021
rect 378 1008 894 1011
rect 1290 1008 1294 1011
rect 1410 1008 1534 1011
rect 1658 1008 1902 1011
rect 2034 1008 2070 1011
rect 2762 1008 3174 1011
rect 3442 1008 3830 1011
rect 3834 1008 4102 1011
rect 4498 1008 4526 1011
rect 4642 1008 4758 1011
rect 4794 1008 5110 1011
rect 328 1003 330 1007
rect 334 1003 337 1007
rect 342 1003 344 1007
rect 1352 1003 1354 1007
rect 1358 1003 1361 1007
rect 1366 1003 1368 1007
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2398 1003 2400 1007
rect 3400 1003 3402 1007
rect 3406 1003 3409 1007
rect 3414 1003 3416 1007
rect 4424 1003 4426 1007
rect 4430 1003 4433 1007
rect 4438 1003 4440 1007
rect 162 998 222 1001
rect 474 998 950 1001
rect 1050 998 1238 1001
rect 1442 998 1446 1001
rect 1618 998 1654 1001
rect 2770 998 3142 1001
rect 3466 998 3582 1001
rect 3586 998 3622 1001
rect 3770 998 3782 1001
rect 4194 998 4414 1001
rect 4562 998 4590 1001
rect 5270 992 5273 998
rect 634 988 670 991
rect 674 988 718 991
rect 754 988 942 991
rect 1034 988 1094 991
rect 1098 988 1222 991
rect 1242 988 1278 991
rect 1322 988 1422 991
rect 1426 988 1462 991
rect 2002 988 2054 991
rect 2074 988 2126 991
rect 2586 988 3510 991
rect 3690 988 3774 991
rect 3786 988 3958 991
rect 3978 988 4142 991
rect 4202 988 4238 991
rect 4434 988 4446 991
rect 4490 988 5150 991
rect 5226 988 5262 991
rect 198 978 438 981
rect 566 978 646 981
rect 834 978 1774 981
rect 1906 978 1918 981
rect 2106 978 2198 981
rect 2562 978 2670 981
rect 2674 978 2710 981
rect 2834 978 3046 981
rect 3146 978 3542 981
rect 3754 978 4126 981
rect 4130 978 4134 981
rect 4258 978 4649 981
rect 4658 978 5014 981
rect 198 972 201 978
rect 566 972 569 978
rect 106 968 137 971
rect 134 962 137 968
rect 258 968 310 971
rect 318 968 326 971
rect 330 968 398 971
rect 686 971 689 978
rect 686 968 942 971
rect 958 968 982 971
rect 1002 968 1158 971
rect 1162 968 1494 971
rect 1498 968 1518 971
rect 1970 968 1998 971
rect 2010 968 2030 971
rect 2038 968 2046 971
rect 2050 968 2054 971
rect 2098 968 2134 971
rect 2594 968 2630 971
rect 2634 968 2694 971
rect 2718 971 2721 978
rect 4646 972 4649 978
rect 2718 968 2918 971
rect 2962 968 3094 971
rect 3106 968 3494 971
rect 3738 968 3782 971
rect 3794 968 4198 971
rect 4290 968 4454 971
rect 4714 968 4806 971
rect 4858 968 5054 971
rect 5194 968 5278 971
rect 182 962 185 968
rect 958 962 961 968
rect 4206 962 4209 968
rect 42 958 118 961
rect 138 958 166 961
rect 274 958 286 961
rect 322 958 334 961
rect 354 958 414 961
rect 658 958 702 961
rect 834 958 846 961
rect 978 958 982 961
rect 1026 958 1030 961
rect 1266 958 1286 961
rect 1446 958 1454 961
rect 1458 958 1558 961
rect 1690 958 1966 961
rect 1970 958 2070 961
rect 2122 958 2134 961
rect 2338 958 2430 961
rect 2434 958 2558 961
rect 2562 958 2606 961
rect 2642 958 2646 961
rect 2666 958 2702 961
rect 2746 958 2758 961
rect 2786 958 2790 961
rect 2858 958 2910 961
rect 3058 958 3166 961
rect 3178 958 3310 961
rect 3738 958 3758 961
rect 4274 958 4446 961
rect 4450 958 4638 961
rect 4754 958 4758 961
rect 4922 958 4926 961
rect 4938 958 4998 961
rect 5002 958 5150 961
rect 5218 958 5286 961
rect 234 948 254 951
rect 262 951 265 958
rect 262 948 270 951
rect 274 948 342 951
rect 394 948 422 951
rect 470 951 473 958
rect 470 948 478 951
rect 554 948 582 951
rect 586 948 598 951
rect 674 948 678 951
rect 734 951 737 958
rect 698 948 737 951
rect 814 952 817 958
rect 1118 952 1121 958
rect 1166 952 1169 958
rect 1174 952 1177 958
rect 1414 952 1417 958
rect 1670 952 1673 958
rect 2806 952 2809 958
rect 906 948 910 951
rect 970 948 998 951
rect 1050 948 1062 951
rect 1126 948 1134 951
rect 1274 948 1302 951
rect 1306 948 1334 951
rect 1434 948 1446 951
rect 1658 948 1662 951
rect 1714 948 1742 951
rect 1746 948 1974 951
rect 1978 948 1990 951
rect 1994 948 2022 951
rect 2026 948 2134 951
rect 2138 948 2246 951
rect 2266 948 2270 951
rect 2298 948 2302 951
rect 2326 948 2374 951
rect 2482 948 2510 951
rect 2514 948 2654 951
rect 2682 948 2710 951
rect 2914 948 2958 951
rect 3010 948 3078 951
rect 3122 948 3278 951
rect 3318 951 3321 958
rect 3446 952 3449 958
rect 3470 952 3473 958
rect 3798 952 3801 958
rect 3318 948 3438 951
rect 3474 948 3486 951
rect 3674 948 3750 951
rect 3802 948 3974 951
rect 4074 948 4078 951
rect 4210 948 4222 951
rect 4474 948 4478 951
rect 4618 948 4622 951
rect 4674 948 4694 951
rect 4786 948 4878 951
rect 4882 948 4926 951
rect 4938 948 4998 951
rect 5066 948 5102 951
rect 5210 948 5214 951
rect 5334 951 5338 952
rect 5290 948 5338 951
rect 114 938 118 941
rect 226 938 238 941
rect 290 938 686 941
rect 938 938 958 941
rect 1038 941 1041 948
rect 1038 938 1078 941
rect 1102 941 1105 948
rect 1678 942 1681 948
rect 2326 942 2329 948
rect 4510 942 4513 948
rect 1102 938 1214 941
rect 1218 938 1222 941
rect 1246 938 1318 941
rect 1482 938 1502 941
rect 1730 938 1806 941
rect 1914 938 1985 941
rect 2026 938 2038 941
rect 2074 938 2081 941
rect 2090 938 2110 941
rect 2114 938 2262 941
rect 2338 938 2422 941
rect 2450 938 2462 941
rect 2522 938 2598 941
rect 2658 938 2702 941
rect 2714 938 2750 941
rect 2778 938 2782 941
rect 2874 938 2902 941
rect 2906 938 2974 941
rect 2978 938 3086 941
rect 3250 938 3286 941
rect 3362 938 3478 941
rect 3522 938 3550 941
rect 3554 938 3574 941
rect 3594 938 3606 941
rect 3626 938 3710 941
rect 3714 938 3726 941
rect 3730 938 3734 941
rect 3918 938 3993 941
rect 4074 938 4134 941
rect 4138 938 4174 941
rect 4194 938 4262 941
rect 4374 938 4398 941
rect 4474 938 4478 941
rect 4490 938 4494 941
rect 4618 938 4838 941
rect 4842 938 4862 941
rect 4866 938 4894 941
rect 4922 938 4966 941
rect 5038 941 5041 948
rect 5134 941 5137 948
rect 5038 938 5206 941
rect 1246 932 1249 938
rect 1982 932 1985 938
rect 2078 932 2081 938
rect 3142 932 3145 938
rect 3918 932 3921 938
rect 3990 932 3993 938
rect 4374 932 4377 938
rect 466 928 478 931
rect 514 928 598 931
rect 634 928 646 931
rect 898 928 1086 931
rect 1114 928 1118 931
rect 1490 928 1966 931
rect 2050 928 2070 931
rect 2258 928 2270 931
rect 2410 928 2846 931
rect 2898 928 2966 931
rect 2986 928 2998 931
rect 3002 928 3102 931
rect 3442 928 3518 931
rect 3826 928 3870 931
rect 4018 928 4097 931
rect 4226 928 4302 931
rect 4410 928 4502 931
rect 4618 928 4742 931
rect 4914 928 4942 931
rect 4986 928 5038 931
rect 154 918 166 921
rect 186 918 206 921
rect 398 921 401 928
rect 4094 922 4097 928
rect 398 918 886 921
rect 978 918 1198 921
rect 1338 918 1638 921
rect 1722 918 1766 921
rect 1810 918 1950 921
rect 1954 918 2022 921
rect 2058 918 2182 921
rect 2186 918 2318 921
rect 2362 918 2606 921
rect 2642 918 2710 921
rect 2762 918 2854 921
rect 2986 918 3134 921
rect 3194 918 3670 921
rect 3730 918 3750 921
rect 3754 918 3774 921
rect 3914 918 3950 921
rect 4322 918 4374 921
rect 4514 918 4542 921
rect 4562 918 4590 921
rect 4738 918 4742 921
rect 4882 918 4958 921
rect 5018 918 5182 921
rect 5242 918 5254 921
rect 894 912 897 918
rect 122 908 406 911
rect 450 908 486 911
rect 578 908 654 911
rect 1122 908 1478 911
rect 1506 908 1542 911
rect 1546 908 1702 911
rect 1730 908 1830 911
rect 2122 908 2126 911
rect 2178 908 2182 911
rect 2234 908 2302 911
rect 2306 908 2350 911
rect 3506 908 3902 911
rect 3962 908 4198 911
rect 4202 908 4222 911
rect 4282 908 4342 911
rect 4450 908 4686 911
rect 4690 908 4814 911
rect 5058 908 5078 911
rect 5250 908 5254 911
rect 848 903 850 907
rect 854 903 857 907
rect 862 903 864 907
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1886 903 1888 907
rect 162 898 294 901
rect 298 898 606 901
rect 634 898 662 901
rect 826 898 830 901
rect 890 898 918 901
rect 922 898 934 901
rect 1018 898 1046 901
rect 1226 898 1390 901
rect 1458 898 1534 901
rect 1538 898 1686 901
rect 1994 898 2006 901
rect 2230 901 2233 908
rect 2888 903 2890 907
rect 2894 903 2897 907
rect 2902 903 2904 907
rect 3920 903 3922 907
rect 3926 903 3929 907
rect 3934 903 3936 907
rect 4936 903 4938 907
rect 4942 903 4945 907
rect 4950 903 4952 907
rect 2058 898 2233 901
rect 2330 898 2358 901
rect 2730 898 2838 901
rect 3658 898 3718 901
rect 3770 898 3814 901
rect 4090 898 4094 901
rect 4098 898 4110 901
rect 4154 898 4182 901
rect 4218 898 4534 901
rect 4538 898 4598 901
rect 5242 898 5262 901
rect 106 888 150 891
rect 242 888 334 891
rect 338 888 494 891
rect 650 888 718 891
rect 986 888 1070 891
rect 1198 888 1230 891
rect 1234 888 1270 891
rect 1338 888 1542 891
rect 1762 888 1862 891
rect 1866 888 1910 891
rect 2082 888 2174 891
rect 2258 888 2926 891
rect 2938 888 3049 891
rect 150 881 153 888
rect 1198 882 1201 888
rect 3046 882 3049 888
rect 3146 888 3257 891
rect 3314 888 3366 891
rect 3498 888 3526 891
rect 3906 888 3950 891
rect 3962 888 4006 891
rect 4010 888 4094 891
rect 4506 888 4526 891
rect 4530 888 4550 891
rect 4582 888 4614 891
rect 4802 888 4822 891
rect 4962 888 5150 891
rect 3070 882 3073 888
rect 3094 882 3097 888
rect 3254 882 3257 888
rect 3822 882 3825 888
rect 4102 882 4105 888
rect 4582 882 4585 888
rect 150 878 166 881
rect 178 878 246 881
rect 426 878 486 881
rect 714 878 766 881
rect 786 878 878 881
rect 882 878 958 881
rect 1050 878 1054 881
rect 1330 878 1422 881
rect 1706 878 2086 881
rect 2090 878 2150 881
rect 2218 878 2222 881
rect 2226 878 2270 881
rect 2474 878 2494 881
rect 2514 878 2518 881
rect 2694 878 2702 881
rect 2706 878 2774 881
rect 2858 878 3038 881
rect 3098 878 3182 881
rect 3258 878 3358 881
rect 3386 878 3438 881
rect 3442 878 3462 881
rect 3466 878 3542 881
rect 3546 878 3766 881
rect 3970 878 4014 881
rect 4258 878 4286 881
rect 4458 878 4542 881
rect 4594 878 4598 881
rect 4698 878 4766 881
rect 4934 881 4937 888
rect 4842 878 4937 881
rect 5002 878 5166 881
rect 170 868 182 871
rect 546 868 590 871
rect 618 868 638 871
rect 662 871 665 878
rect 662 868 830 871
rect 834 868 886 871
rect 938 868 942 871
rect 1118 871 1121 878
rect 1686 872 1689 878
rect 1694 872 1697 878
rect 982 868 1121 871
rect 1146 868 1246 871
rect 1262 868 1454 871
rect 1466 868 1470 871
rect 1570 868 1654 871
rect 1714 868 1718 871
rect 1826 868 1918 871
rect 1954 868 1982 871
rect 1986 868 2110 871
rect 2218 868 2246 871
rect 2430 871 2433 878
rect 3806 872 3809 878
rect 4678 872 4681 878
rect 2354 868 2433 871
rect 2450 868 2526 871
rect 2650 868 2798 871
rect 2802 868 2814 871
rect 2866 868 3078 871
rect 3090 868 3358 871
rect 3362 868 3366 871
rect 3370 868 3390 871
rect 3426 868 3430 871
rect 3458 868 3486 871
rect 3674 868 3678 871
rect 3818 868 3974 871
rect 3978 868 4054 871
rect 4066 868 4118 871
rect 4210 868 4358 871
rect 4370 868 4473 871
rect 4498 868 4606 871
rect 4706 868 4718 871
rect 4906 868 4966 871
rect 4986 868 5006 871
rect 5010 868 5158 871
rect 5210 868 5238 871
rect 462 862 465 868
rect 50 858 126 861
rect 330 858 401 861
rect 466 858 486 861
rect 506 858 574 861
rect 578 858 582 861
rect 618 858 622 861
rect 682 858 710 861
rect 714 858 798 861
rect 818 858 862 861
rect 866 858 926 861
rect 982 861 985 868
rect 1262 862 1265 868
rect 946 858 985 861
rect 1066 858 1254 861
rect 1418 858 1462 861
rect 1626 858 1646 861
rect 1650 858 1694 861
rect 1706 858 1734 861
rect 1738 858 1758 861
rect 1786 858 1830 861
rect 1882 859 1958 861
rect 1878 858 1958 859
rect 1978 858 2158 861
rect 2270 861 2273 868
rect 2218 858 2273 861
rect 2378 858 2382 861
rect 2402 858 2414 861
rect 2590 861 2593 868
rect 3494 862 3497 868
rect 3798 862 3801 868
rect 2590 858 2606 861
rect 2722 858 2814 861
rect 2930 858 2974 861
rect 2986 858 2990 861
rect 3066 858 3081 861
rect 3090 858 3118 861
rect 3138 858 3182 861
rect 3206 858 3270 861
rect 3350 858 3406 861
rect 3410 858 3462 861
rect 3634 858 3646 861
rect 3658 858 3662 861
rect 3722 858 3726 861
rect 3738 858 3742 861
rect 3874 858 3918 861
rect 3970 858 3974 861
rect 4150 861 4153 868
rect 4470 862 4473 868
rect 5182 862 5185 868
rect 3994 858 4153 861
rect 4218 858 4238 861
rect 4242 858 4310 861
rect 4314 858 4342 861
rect 4394 858 4406 861
rect 4422 858 4454 861
rect 4530 858 4990 861
rect 4994 858 5054 861
rect 5058 858 5086 861
rect 5090 858 5126 861
rect 5246 861 5249 868
rect 5202 858 5249 861
rect 106 848 174 851
rect 214 851 217 858
rect 398 852 401 858
rect 214 848 382 851
rect 434 848 470 851
rect 506 848 550 851
rect 674 848 686 851
rect 722 848 806 851
rect 906 848 918 851
rect 1098 848 1214 851
rect 1234 848 1238 851
rect 1250 848 1630 851
rect 1634 848 1670 851
rect 1714 848 1718 851
rect 1746 848 1806 851
rect 1850 848 2190 851
rect 2218 848 2225 851
rect 114 838 134 841
rect 138 838 422 841
rect 830 841 833 848
rect 2222 842 2225 848
rect 2458 848 2462 851
rect 2610 848 2614 851
rect 2634 848 2638 851
rect 2826 848 2958 851
rect 3014 851 3017 858
rect 2978 848 3017 851
rect 3046 851 3049 858
rect 3026 848 3049 851
rect 3078 852 3081 858
rect 3206 852 3209 858
rect 3350 852 3353 858
rect 3186 848 3206 851
rect 3490 848 3510 851
rect 3794 848 3838 851
rect 3854 851 3857 858
rect 3842 848 3857 851
rect 3870 848 3889 851
rect 3946 848 3950 851
rect 3954 848 4094 851
rect 4202 848 4238 851
rect 4266 848 4270 851
rect 4422 851 4425 858
rect 4286 848 4425 851
rect 4434 848 4502 851
rect 4594 848 4614 851
rect 4618 848 4998 851
rect 5098 848 5102 851
rect 762 838 833 841
rect 850 838 1102 841
rect 1122 838 1302 841
rect 1466 838 1742 841
rect 1754 838 1982 841
rect 2238 841 2241 848
rect 3870 842 3873 848
rect 3886 842 3889 848
rect 4286 842 4289 848
rect 5030 842 5033 848
rect 2238 838 2286 841
rect 2290 838 2326 841
rect 2394 838 2462 841
rect 2490 838 2550 841
rect 2554 838 2926 841
rect 2986 838 2990 841
rect 3042 838 3046 841
rect 3122 838 3358 841
rect 3790 838 3798 841
rect 3802 838 3806 841
rect 4082 838 4230 841
rect 4394 838 4454 841
rect 4514 838 4638 841
rect 4642 838 4662 841
rect 4898 838 4918 841
rect 4922 838 5022 841
rect 82 828 494 831
rect 498 828 718 831
rect 802 828 918 831
rect 1082 828 1134 831
rect 1170 828 1310 831
rect 1314 828 1374 831
rect 1594 828 1718 831
rect 2178 828 2342 831
rect 2346 828 2598 831
rect 2602 828 2654 831
rect 2658 828 2710 831
rect 2818 828 2830 831
rect 2834 828 2910 831
rect 2914 828 3206 831
rect 3674 828 4174 831
rect 4186 828 4198 831
rect 4258 828 4446 831
rect 4474 828 4742 831
rect 5018 828 5046 831
rect 250 818 710 821
rect 714 818 1238 821
rect 1246 818 1518 821
rect 1610 818 1854 821
rect 1930 818 2142 821
rect 2426 818 2742 821
rect 2762 818 2934 821
rect 3082 818 4462 821
rect 4642 818 4718 821
rect 4898 818 5038 821
rect 5042 818 5158 821
rect 5266 818 5278 821
rect 1246 812 1249 818
rect 354 808 358 811
rect 490 808 902 811
rect 914 808 1182 811
rect 1618 808 1622 811
rect 1770 808 1782 811
rect 2418 808 2422 811
rect 2586 808 2598 811
rect 2602 808 2646 811
rect 3034 808 3078 811
rect 3554 808 3558 811
rect 3698 808 3878 811
rect 3890 808 4158 811
rect 4178 808 4390 811
rect 4730 808 4966 811
rect 5090 808 5158 811
rect 328 803 330 807
rect 334 803 337 807
rect 342 803 344 807
rect 1352 803 1354 807
rect 1358 803 1361 807
rect 1366 803 1368 807
rect 2062 802 2065 808
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2398 803 2400 807
rect 3400 803 3402 807
rect 3406 803 3409 807
rect 3414 803 3416 807
rect 4166 802 4169 808
rect 4424 803 4426 807
rect 4430 803 4433 807
rect 4438 803 4440 807
rect 4494 802 4497 808
rect 618 798 630 801
rect 778 798 822 801
rect 986 798 1062 801
rect 1410 798 1590 801
rect 1618 798 2030 801
rect 2138 798 2294 801
rect 2826 798 2926 801
rect 2930 798 2998 801
rect 3242 798 3318 801
rect 3538 798 3702 801
rect 4018 798 4150 801
rect 4506 798 4614 801
rect 4658 798 5102 801
rect 130 788 246 791
rect 250 788 518 791
rect 522 788 1206 791
rect 1298 788 1374 791
rect 1386 788 1646 791
rect 1682 788 1742 791
rect 1746 788 1766 791
rect 1770 788 1990 791
rect 2090 788 2630 791
rect 3066 788 3086 791
rect 3210 788 3302 791
rect 3306 788 3566 791
rect 3570 788 3814 791
rect 3850 788 3886 791
rect 3890 788 4038 791
rect 4354 788 4497 791
rect 4654 791 4657 798
rect 4506 788 4657 791
rect 5126 792 5129 798
rect 4494 782 4497 788
rect 178 778 318 781
rect 418 778 662 781
rect 666 778 822 781
rect 826 778 1014 781
rect 1018 778 1046 781
rect 1194 778 1262 781
rect 1290 778 1790 781
rect 1986 778 2398 781
rect 2402 778 2454 781
rect 2906 778 3310 781
rect 3314 778 3462 781
rect 3522 778 3542 781
rect 3546 778 3566 781
rect 4058 778 4086 781
rect 4170 778 4382 781
rect 4418 778 4430 781
rect 4834 778 4958 781
rect 5166 781 5169 788
rect 5130 778 5169 781
rect 122 768 262 771
rect 410 768 622 771
rect 626 768 1326 771
rect 1698 768 1822 771
rect 2042 768 2118 771
rect 2130 768 2158 771
rect 2162 768 2214 771
rect 2434 768 2590 771
rect 2878 771 2881 778
rect 2878 768 2910 771
rect 3034 768 3334 771
rect 3530 768 3862 771
rect 3866 768 3950 771
rect 3954 768 4062 771
rect 4074 768 4134 771
rect 4154 768 4446 771
rect 4458 768 4814 771
rect 4898 768 5086 771
rect 5258 768 5262 771
rect 170 758 198 761
rect 314 758 358 761
rect 434 758 502 761
rect 722 758 854 761
rect 874 758 934 761
rect 1042 758 1118 761
rect 1154 758 1190 761
rect 1326 761 1329 768
rect 1326 758 1422 761
rect 1426 758 1750 761
rect 1890 758 2022 761
rect 2302 761 2305 768
rect 2282 758 2305 761
rect 2322 758 2326 761
rect 2354 758 2446 761
rect 2638 761 2641 768
rect 2618 758 2641 761
rect 2862 761 2865 768
rect 3022 762 3025 768
rect 2842 758 2865 761
rect 2890 758 2918 761
rect 3098 758 3134 761
rect 3138 758 3230 761
rect 3386 758 3446 761
rect 3498 758 3502 761
rect 3514 758 3678 761
rect 3698 758 3801 761
rect 3922 758 3966 761
rect 3970 758 3998 761
rect 4050 758 4078 761
rect 4114 758 4142 761
rect 4146 758 4150 761
rect 4162 758 4294 761
rect 4306 758 4422 761
rect 4426 758 4438 761
rect 4578 758 4606 761
rect 4818 758 5006 761
rect 5010 758 5094 761
rect 5150 761 5153 768
rect 5150 758 5222 761
rect 34 748 38 751
rect 66 748 102 751
rect 162 748 209 751
rect 234 748 254 751
rect 258 748 278 751
rect 362 748 377 751
rect 426 748 454 751
rect 458 748 462 751
rect 646 751 649 758
rect 998 752 1001 758
rect 578 748 649 751
rect 762 748 766 751
rect 778 748 798 751
rect 818 748 830 751
rect 1058 748 1078 751
rect 18 738 30 741
rect 102 741 105 748
rect 118 741 121 748
rect 102 738 121 741
rect 206 742 209 748
rect 374 742 377 748
rect 1198 751 1201 758
rect 1194 748 1201 751
rect 1226 748 1230 751
rect 1282 748 1334 751
rect 1458 748 1526 751
rect 1666 748 1750 751
rect 1850 748 1854 751
rect 2002 748 2030 751
rect 2158 751 2161 758
rect 2090 748 2161 751
rect 2238 752 2241 758
rect 2310 752 2313 758
rect 3798 752 3801 758
rect 4030 752 4033 758
rect 2250 748 2254 751
rect 2338 748 2414 751
rect 2650 748 2918 751
rect 2962 748 2990 751
rect 3042 748 3046 751
rect 3166 748 3222 751
rect 3274 748 3302 751
rect 3306 748 3358 751
rect 3450 748 3502 751
rect 3562 748 3566 751
rect 3714 748 3718 751
rect 3958 748 3974 751
rect 3986 748 3993 751
rect 4010 748 4014 751
rect 4146 748 4342 751
rect 4554 748 4574 751
rect 4610 748 4622 751
rect 4774 751 4777 758
rect 5118 752 5121 758
rect 4770 748 4777 751
rect 4794 748 4798 751
rect 4874 748 4878 751
rect 4990 748 5030 751
rect 5050 748 5054 751
rect 5082 748 5102 751
rect 5162 748 5174 751
rect 378 738 414 741
rect 466 738 470 741
rect 578 738 750 741
rect 770 738 774 741
rect 986 738 993 741
rect 1010 738 1342 741
rect 1630 741 1633 748
rect 3054 742 3057 748
rect 3166 742 3169 748
rect 1546 738 1633 741
rect 1714 738 1742 741
rect 1746 738 1758 741
rect 1866 738 2046 741
rect 2074 738 2078 741
rect 2098 738 2110 741
rect 2114 738 2150 741
rect 2266 738 2270 741
rect 2282 738 2286 741
rect 2298 738 2358 741
rect 2626 738 2630 741
rect 2738 738 2782 741
rect 2834 738 3038 741
rect 3246 741 3249 748
rect 3814 742 3817 748
rect 3958 742 3961 748
rect 3990 742 3993 748
rect 3242 738 3249 741
rect 3338 738 3478 741
rect 3482 738 3510 741
rect 3538 738 3550 741
rect 3770 738 3806 741
rect 3882 738 3910 741
rect 3914 738 3934 741
rect 4014 741 4017 748
rect 4966 742 4969 748
rect 4974 742 4977 748
rect 4990 742 4993 748
rect 4014 738 4390 741
rect 4482 738 4646 741
rect 4650 738 4734 741
rect 5002 738 5014 741
rect 5074 738 5198 741
rect 990 732 993 738
rect 1782 732 1785 738
rect 2486 732 2489 738
rect 122 728 230 731
rect 306 728 473 731
rect 482 728 710 731
rect 762 728 782 731
rect 826 728 838 731
rect 842 728 926 731
rect 946 728 982 731
rect 1186 728 1206 731
rect 1218 728 1230 731
rect 1258 728 1302 731
rect 1338 728 1606 731
rect 1866 728 1894 731
rect 1962 728 2009 731
rect 2702 731 2705 738
rect 2830 732 2833 738
rect 2702 728 2774 731
rect 2866 728 2926 731
rect 3078 731 3081 738
rect 3078 728 3313 731
rect 3322 728 3430 731
rect 3550 728 3558 731
rect 3562 728 3614 731
rect 3810 728 3814 731
rect 3974 731 3977 738
rect 3866 728 3977 731
rect 3986 728 4062 731
rect 4090 728 4094 731
rect 4122 728 4182 731
rect 4194 728 4222 731
rect 4282 728 4334 731
rect 4450 728 4694 731
rect 4778 728 4793 731
rect 4930 728 5006 731
rect 5010 728 5038 731
rect 5050 728 5158 731
rect 5186 728 5262 731
rect 5274 728 5278 731
rect 470 722 473 728
rect 2006 722 2009 728
rect 2974 722 2977 728
rect 2990 722 2993 728
rect 3014 722 3017 728
rect 186 718 190 721
rect 274 718 390 721
rect 498 718 718 721
rect 730 718 878 721
rect 946 718 1054 721
rect 1234 718 1350 721
rect 1354 718 1470 721
rect 1522 718 1534 721
rect 1674 718 1718 721
rect 1722 718 1905 721
rect 2362 718 2398 721
rect 2490 718 2606 721
rect 2722 718 2910 721
rect 3042 718 3150 721
rect 3154 718 3206 721
rect 3310 721 3313 728
rect 4414 722 4417 728
rect 4790 722 4793 728
rect 3310 718 3406 721
rect 3426 718 3606 721
rect 3610 718 3734 721
rect 3818 718 4086 721
rect 4106 718 4326 721
rect 4458 718 4654 721
rect 4954 718 4982 721
rect 5026 718 5062 721
rect 5066 718 5094 721
rect 1902 712 1905 718
rect 178 708 318 711
rect 354 708 366 711
rect 370 708 478 711
rect 514 708 702 711
rect 810 708 830 711
rect 1290 708 1398 711
rect 1434 708 1502 711
rect 1506 708 1526 711
rect 1642 708 1782 711
rect 1802 708 1854 711
rect 1858 708 1862 711
rect 1906 708 2246 711
rect 2250 708 2662 711
rect 2938 708 2982 711
rect 2986 708 3774 711
rect 4106 708 4150 711
rect 4154 708 4222 711
rect 4226 708 4454 711
rect 4514 708 4542 711
rect 4562 708 4758 711
rect 848 703 850 707
rect 854 703 857 707
rect 862 703 864 707
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1886 703 1888 707
rect 2888 703 2890 707
rect 2894 703 2897 707
rect 2902 703 2904 707
rect 3920 703 3922 707
rect 3926 703 3929 707
rect 3934 703 3936 707
rect 234 698 366 701
rect 450 698 486 701
rect 562 698 638 701
rect 1274 698 1798 701
rect 1962 698 1966 701
rect 1994 698 2174 701
rect 2186 698 2262 701
rect 2442 698 2590 701
rect 2690 698 2862 701
rect 3066 698 3078 701
rect 3106 698 3302 701
rect 3306 698 3318 701
rect 3330 698 3494 701
rect 3498 698 3614 701
rect 3618 698 3638 701
rect 3650 698 3782 701
rect 3786 698 3870 701
rect 4066 698 4142 701
rect 4146 698 4174 701
rect 4402 698 4510 701
rect 4558 701 4561 708
rect 4936 703 4938 707
rect 4942 703 4945 707
rect 4950 703 4952 707
rect 4514 698 4561 701
rect 4794 698 4878 701
rect 5002 698 5126 701
rect 226 688 438 691
rect 474 688 478 691
rect 610 688 670 691
rect 674 688 726 691
rect 1090 688 1142 691
rect 1290 688 1542 691
rect 1618 688 1678 691
rect 1850 688 2006 691
rect 2170 688 2230 691
rect 2234 688 2241 691
rect 2838 688 2878 691
rect 2886 688 2894 691
rect 2898 688 2982 691
rect 3074 688 3142 691
rect 3146 688 3286 691
rect 3298 688 3430 691
rect 3674 688 3686 691
rect 3690 688 3710 691
rect 3714 688 3982 691
rect 4058 688 4190 691
rect 4402 688 4614 691
rect 4618 688 4726 691
rect 4890 688 4934 691
rect 5010 688 5166 691
rect 130 678 262 681
rect 362 678 374 681
rect 450 678 534 681
rect 538 678 734 681
rect 738 678 758 681
rect 878 681 881 688
rect 878 678 1094 681
rect 1210 678 1318 681
rect 1394 678 1574 681
rect 1686 681 1689 688
rect 2838 682 2841 688
rect 3454 682 3457 688
rect 1686 678 1774 681
rect 1794 678 2070 681
rect 2090 678 2094 681
rect 2194 678 2278 681
rect 2370 678 2438 681
rect 2442 678 2486 681
rect 2514 678 2606 681
rect 2714 678 2814 681
rect 2874 678 2958 681
rect 2962 678 3046 681
rect 3050 678 3110 681
rect 3170 678 3390 681
rect 3498 678 3502 681
rect 3526 681 3529 688
rect 3526 678 3550 681
rect 3874 678 3926 681
rect 3994 678 4038 681
rect 4090 678 4113 681
rect 4194 678 4198 681
rect 4530 678 4574 681
rect 4578 678 4590 681
rect 4610 678 4654 681
rect 4674 678 4678 681
rect 4854 681 4857 688
rect 4854 678 4910 681
rect 4990 681 4993 688
rect 4938 678 4993 681
rect 5006 682 5009 688
rect 5050 678 5062 681
rect 66 668 94 671
rect 106 668 134 671
rect 162 668 206 671
rect 210 668 214 671
rect 274 668 294 671
rect 390 671 393 678
rect 1198 672 1201 678
rect 1374 672 1377 678
rect 390 668 670 671
rect 970 668 998 671
rect 1050 668 1054 671
rect 1058 668 1110 671
rect 1146 668 1174 671
rect 1618 668 1654 671
rect 1722 668 1798 671
rect 1850 668 1926 671
rect 1930 668 1966 671
rect 2046 668 2142 671
rect 2226 668 2246 671
rect 2258 668 2334 671
rect 2338 668 2406 671
rect 2418 668 2454 671
rect 2578 668 2622 671
rect 2658 668 2694 671
rect 2714 668 2742 671
rect 2754 668 2846 671
rect 2866 668 2966 671
rect 2970 668 3094 671
rect 3122 668 3126 671
rect 3426 668 3430 671
rect 3718 671 3721 678
rect 3838 672 3841 678
rect 4062 672 4065 678
rect 4110 672 4113 678
rect 3718 668 3766 671
rect 3770 668 3814 671
rect 3842 668 3862 671
rect 3914 668 3982 671
rect 3986 668 3993 671
rect 4018 668 4030 671
rect 4306 668 4310 671
rect 4390 671 4393 678
rect 4314 668 4478 671
rect 4570 668 4686 671
rect 4914 668 5014 671
rect 5150 671 5153 678
rect 5150 668 5246 671
rect 38 661 41 668
rect 302 662 305 668
rect 870 662 873 668
rect 38 658 54 661
rect 74 658 118 661
rect 130 658 278 661
rect 282 658 302 661
rect 370 658 406 661
rect 410 658 422 661
rect 634 658 646 661
rect 706 658 710 661
rect 1002 658 1006 661
rect 1066 658 1190 661
rect 1214 658 1222 661
rect 1270 661 1273 668
rect 1226 658 1273 661
rect 1450 658 1454 661
rect 1490 658 1494 661
rect 1570 658 1625 661
rect 1650 658 1678 661
rect 1822 661 1825 668
rect 1818 658 1825 661
rect 2046 662 2049 668
rect 2074 658 2214 661
rect 2250 658 2270 661
rect 2274 658 2342 661
rect 2482 658 2494 661
rect 2634 658 2646 661
rect 2706 658 2726 661
rect 2818 658 2894 661
rect 2898 658 2942 661
rect 3034 658 3126 661
rect 3146 658 3198 661
rect 3438 661 3441 668
rect 3438 658 3454 661
rect 3502 661 3505 668
rect 3502 658 3526 661
rect 3538 658 3542 661
rect 3622 661 3625 668
rect 3990 662 3993 668
rect 4126 662 4129 668
rect 3622 658 3686 661
rect 3714 658 3870 661
rect 4002 658 4006 661
rect 4026 658 4038 661
rect 4202 658 4206 661
rect 4298 658 4302 661
rect 4410 658 4502 661
rect 4530 658 4550 661
rect 4554 658 4582 661
rect 4610 658 4641 661
rect 4658 658 4670 661
rect 4714 658 4718 661
rect 4806 661 4809 668
rect 4806 658 4870 661
rect 4902 661 4905 668
rect 5062 662 5065 668
rect 4898 658 4905 661
rect 4922 658 4958 661
rect 5042 658 5046 661
rect 5070 661 5073 668
rect 5070 658 5110 661
rect 1382 652 1385 658
rect 1622 652 1625 658
rect 1806 652 1809 658
rect 4078 652 4081 658
rect 4638 652 4641 658
rect 50 648 350 651
rect 394 648 486 651
rect 666 648 710 651
rect 754 648 886 651
rect 1250 648 1366 651
rect 1666 648 1726 651
rect 1950 648 1958 651
rect 1962 648 2022 651
rect 2106 648 2334 651
rect 2346 648 2406 651
rect 2710 648 2750 651
rect 2826 648 2849 651
rect 2866 648 2870 651
rect 2962 648 2969 651
rect 1702 642 1705 648
rect 2710 642 2713 648
rect 2846 642 2849 648
rect 2966 642 2969 648
rect 2982 648 3078 651
rect 3102 648 3121 651
rect 2982 642 2985 648
rect 3102 642 3105 648
rect 3118 642 3121 648
rect 3170 648 3190 651
rect 3442 648 3462 651
rect 3482 648 3566 651
rect 3570 648 3670 651
rect 3678 648 3686 651
rect 3762 648 3846 651
rect 3962 648 4070 651
rect 4178 648 4302 651
rect 4306 648 4318 651
rect 4834 648 4934 651
rect 4954 648 5006 651
rect 5034 648 5038 651
rect 5050 648 5086 651
rect 5090 648 5166 651
rect 3166 642 3169 648
rect 3678 642 3681 648
rect 58 638 78 641
rect 258 638 273 641
rect 482 638 494 641
rect 650 638 678 641
rect 762 638 902 641
rect 906 638 1278 641
rect 1514 638 1598 641
rect 1602 638 1702 641
rect 1802 638 2014 641
rect 2082 638 2110 641
rect 2130 638 2206 641
rect 2222 638 2238 641
rect 2250 638 2406 641
rect 3258 638 3366 641
rect 3370 638 3422 641
rect 3426 638 3510 641
rect 3514 638 3662 641
rect 4310 638 4318 641
rect 4322 638 4606 641
rect 4634 638 5030 641
rect 5034 638 5073 641
rect 174 632 177 638
rect 270 632 273 638
rect 2222 632 2225 638
rect 5070 632 5073 638
rect 618 628 798 631
rect 842 628 990 631
rect 1018 628 1510 631
rect 1634 628 1678 631
rect 2362 628 2502 631
rect 2746 628 3174 631
rect 3186 628 3262 631
rect 3450 628 3582 631
rect 3634 628 3806 631
rect 3946 628 4446 631
rect 4450 628 4702 631
rect 4978 628 4982 631
rect 338 618 646 621
rect 674 618 1902 621
rect 1914 618 2102 621
rect 2386 618 2654 621
rect 2914 618 2966 621
rect 3050 618 3534 621
rect 3546 618 4086 621
rect 4202 618 4342 621
rect 4402 618 4494 621
rect 4498 618 4710 621
rect 4738 618 4806 621
rect 4826 618 5078 621
rect 194 608 198 611
rect 490 608 518 611
rect 522 608 542 611
rect 746 608 758 611
rect 850 608 1334 611
rect 1578 608 1942 611
rect 1946 608 2030 611
rect 2042 608 2062 611
rect 3002 608 3182 611
rect 3426 608 3518 611
rect 4490 608 4654 611
rect 4770 608 4798 611
rect 4874 608 5254 611
rect 328 603 330 607
rect 334 603 337 607
rect 342 603 344 607
rect 1352 603 1354 607
rect 1358 603 1361 607
rect 1366 603 1368 607
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2398 603 2400 607
rect 3400 603 3402 607
rect 3406 603 3409 607
rect 3414 603 3416 607
rect 4424 603 4426 607
rect 4430 603 4433 607
rect 4438 603 4440 607
rect 194 598 318 601
rect 1474 598 1766 601
rect 1770 598 1798 601
rect 1802 598 2033 601
rect 2434 598 2510 601
rect 2650 598 2806 601
rect 2810 598 2918 601
rect 2922 598 3302 601
rect 3690 598 4134 601
rect 4650 598 5294 601
rect 138 588 182 591
rect 290 588 454 591
rect 1066 588 1070 591
rect 1434 588 1486 591
rect 1770 588 1934 591
rect 2030 591 2033 598
rect 2030 588 2446 591
rect 2506 588 3230 591
rect 3562 588 3806 591
rect 3810 588 3886 591
rect 4002 588 4110 591
rect 4138 588 4598 591
rect 362 578 582 581
rect 778 578 870 581
rect 1010 578 1022 581
rect 1402 578 1430 581
rect 1678 581 1681 588
rect 1678 578 1718 581
rect 1786 578 1878 581
rect 2074 578 2198 581
rect 2202 578 3062 581
rect 3066 578 3206 581
rect 3562 578 3702 581
rect 3794 578 3862 581
rect 3882 578 3942 581
rect 3978 578 4030 581
rect 4362 578 4510 581
rect 4666 578 4718 581
rect 4770 578 5182 581
rect 1238 572 1241 578
rect 242 568 398 571
rect 770 568 854 571
rect 986 568 1014 571
rect 1370 568 1398 571
rect 1594 568 1614 571
rect 1658 568 1790 571
rect 1794 568 1910 571
rect 1950 568 1958 571
rect 1962 568 2022 571
rect 2082 568 2094 571
rect 2306 568 2441 571
rect 2490 568 2662 571
rect 2666 568 2790 571
rect 2850 568 2854 571
rect 2858 568 2894 571
rect 2938 568 3134 571
rect 3202 568 3454 571
rect 3610 568 3910 571
rect 3922 568 4006 571
rect 4154 568 4198 571
rect 4218 568 4598 571
rect 4602 568 4638 571
rect 4922 568 5110 571
rect 5138 568 5150 571
rect 210 558 534 561
rect 538 558 542 561
rect 666 558 678 561
rect 774 558 814 561
rect 898 558 918 561
rect 1018 558 1022 561
rect 1046 561 1049 568
rect 1342 562 1345 568
rect 2438 562 2441 568
rect 1046 558 1230 561
rect 1242 558 1302 561
rect 1386 558 1574 561
rect 1610 558 1614 561
rect 1618 558 1638 561
rect 1706 558 1870 561
rect 1874 558 1958 561
rect 1962 558 1982 561
rect 2042 558 2046 561
rect 2098 558 2134 561
rect 2138 558 2182 561
rect 2234 558 2238 561
rect 2282 558 2390 561
rect 2482 558 2486 561
rect 2578 558 2662 561
rect 2666 558 2822 561
rect 2898 558 3017 561
rect 3034 558 3038 561
rect 3130 558 3278 561
rect 3566 561 3569 568
rect 3490 558 3686 561
rect 3690 558 3798 561
rect 3802 558 3902 561
rect 3906 558 3950 561
rect 3978 558 4134 561
rect 4138 558 4222 561
rect 4898 558 4982 561
rect 5034 558 5206 561
rect 126 551 129 558
rect 82 548 129 551
rect 306 548 334 551
rect 338 548 342 551
rect 354 548 358 551
rect 498 548 502 551
rect 774 551 777 558
rect 666 548 777 551
rect 786 548 798 551
rect 802 548 862 551
rect 866 548 942 551
rect 946 548 974 551
rect 978 548 1030 551
rect 1042 548 1086 551
rect 1282 548 1286 551
rect 1298 548 1302 551
rect 1378 548 1422 551
rect 1562 548 1598 551
rect 1602 548 1614 551
rect 1682 548 1686 551
rect 1810 548 1830 551
rect 1978 548 1990 551
rect 1994 548 2374 551
rect 66 538 209 541
rect 234 538 302 541
rect 306 538 313 541
rect 322 538 790 541
rect 810 538 814 541
rect 890 538 950 541
rect 1034 538 1110 541
rect 1114 538 1134 541
rect 1138 538 1150 541
rect 1270 541 1273 548
rect 1266 538 1273 541
rect 1290 538 1305 541
rect 1554 538 1606 541
rect 1790 541 1793 548
rect 2570 548 2630 551
rect 2726 548 2782 551
rect 2882 548 2886 551
rect 3014 551 3017 558
rect 3014 548 3038 551
rect 3202 548 3302 551
rect 3466 548 3494 551
rect 3498 548 3502 551
rect 3586 548 3638 551
rect 3650 548 3694 551
rect 3778 548 3830 551
rect 3834 548 3894 551
rect 3962 548 3982 551
rect 4018 548 4022 551
rect 4154 548 4190 551
rect 4194 548 4214 551
rect 4522 548 4566 551
rect 4570 548 4574 551
rect 4586 548 4590 551
rect 4634 548 4670 551
rect 4738 548 4926 551
rect 4986 548 5086 551
rect 5090 548 5166 551
rect 5170 548 5190 551
rect 2726 542 2729 548
rect 1682 538 1793 541
rect 1802 538 1838 541
rect 1842 538 2054 541
rect 2154 538 2158 541
rect 2170 538 2174 541
rect 2178 538 2286 541
rect 2306 538 2334 541
rect 2370 538 2558 541
rect 2778 538 2806 541
rect 2842 538 2982 541
rect 3006 541 3009 548
rect 3006 538 3294 541
rect 3434 538 3486 541
rect 3530 538 3590 541
rect 3658 538 3670 541
rect 3746 538 3886 541
rect 3990 541 3993 548
rect 3962 538 3993 541
rect 4002 538 4030 541
rect 4170 538 4182 541
rect 4286 541 4289 548
rect 4286 538 4334 541
rect 4346 538 4446 541
rect 4474 538 4534 541
rect 4702 538 4798 541
rect 5002 538 5078 541
rect 5170 538 5174 541
rect 5186 538 5270 541
rect 110 532 113 538
rect 206 532 209 538
rect 1302 532 1305 538
rect 210 528 382 531
rect 506 528 646 531
rect 650 528 958 531
rect 1058 528 1158 531
rect 1506 528 1566 531
rect 1678 531 1681 538
rect 1570 528 1681 531
rect 1706 528 1894 531
rect 1930 528 2014 531
rect 2106 528 2358 531
rect 2362 528 2430 531
rect 2434 528 2446 531
rect 2514 528 2606 531
rect 2626 528 2646 531
rect 2674 528 2854 531
rect 2874 528 3086 531
rect 3098 528 3126 531
rect 3218 528 3222 531
rect 3314 528 3598 531
rect 3730 528 3822 531
rect 3898 528 3942 531
rect 3954 528 4022 531
rect 4150 531 4153 538
rect 4034 528 4153 531
rect 4182 528 4190 531
rect 4194 528 4246 531
rect 4446 531 4449 538
rect 4702 532 4705 538
rect 4446 528 4534 531
rect 4754 528 4934 531
rect 5010 528 5030 531
rect 5034 528 5118 531
rect 5186 528 5214 531
rect 5274 528 5294 531
rect 382 521 385 528
rect 2646 522 2649 528
rect 382 518 566 521
rect 706 518 790 521
rect 802 518 1022 521
rect 1122 518 1230 521
rect 1266 518 1294 521
rect 1666 518 1790 521
rect 1866 518 1998 521
rect 2018 518 2046 521
rect 2050 518 2086 521
rect 2114 518 2118 521
rect 2266 518 2318 521
rect 2658 518 2718 521
rect 3378 518 3478 521
rect 3490 518 3502 521
rect 3794 518 3830 521
rect 3882 518 3982 521
rect 3986 518 4142 521
rect 4514 518 4550 521
rect 4934 521 4937 528
rect 5174 522 5177 528
rect 4934 518 5022 521
rect 5026 518 5054 521
rect 5058 518 5102 521
rect 5106 518 5142 521
rect 2166 512 2169 518
rect 130 508 246 511
rect 250 508 302 511
rect 698 508 710 511
rect 1298 508 1326 511
rect 1346 508 1622 511
rect 1626 508 1742 511
rect 1914 508 1966 511
rect 2026 508 2102 511
rect 2298 508 2318 511
rect 2506 508 2574 511
rect 2634 508 2670 511
rect 2674 508 2686 511
rect 2922 508 3054 511
rect 3074 508 3078 511
rect 3282 508 3606 511
rect 3786 508 3854 511
rect 4098 508 4230 511
rect 4410 508 4438 511
rect 4482 508 4590 511
rect 4650 508 4758 511
rect 4762 508 4894 511
rect 4962 508 5030 511
rect 5042 508 5062 511
rect 5114 508 5158 511
rect 848 503 850 507
rect 854 503 857 507
rect 862 503 864 507
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1886 503 1888 507
rect 2888 503 2890 507
rect 2894 503 2897 507
rect 2902 503 2904 507
rect 3920 503 3922 507
rect 3926 503 3929 507
rect 3934 503 3936 507
rect 4936 503 4938 507
rect 4942 503 4945 507
rect 4950 503 4952 507
rect 5094 502 5097 508
rect 250 498 326 501
rect 546 498 630 501
rect 634 498 686 501
rect 690 498 782 501
rect 946 498 1302 501
rect 1330 498 1334 501
rect 1730 498 1822 501
rect 2026 498 2145 501
rect 2154 498 2182 501
rect 2186 498 2278 501
rect 2282 498 2446 501
rect 2450 498 2726 501
rect 2738 498 2798 501
rect 2802 498 2878 501
rect 3178 498 3574 501
rect 3594 498 3718 501
rect 3722 498 3878 501
rect 3978 498 4006 501
rect 4010 498 4046 501
rect 4170 498 4470 501
rect 4474 498 4542 501
rect 4546 498 4918 501
rect 50 488 182 491
rect 314 488 342 491
rect 346 488 518 491
rect 746 488 817 491
rect 858 488 934 491
rect 1362 488 1438 491
rect 1442 488 1462 491
rect 1570 488 1574 491
rect 1634 488 1654 491
rect 1670 488 1726 491
rect 1738 488 1774 491
rect 1826 488 1926 491
rect 1934 491 1937 498
rect 1934 488 2030 491
rect 2142 491 2145 498
rect 2142 488 2174 491
rect 2178 488 2310 491
rect 2474 488 2734 491
rect 2738 488 2822 491
rect 2930 488 3014 491
rect 3026 488 3030 491
rect 3162 488 3182 491
rect 3298 488 3302 491
rect 3394 488 3542 491
rect 3546 488 4134 491
rect 4154 488 4510 491
rect 4514 488 4526 491
rect 4610 488 4622 491
rect 4922 488 5038 491
rect 5098 488 5102 491
rect 5186 488 5214 491
rect 814 482 817 488
rect 170 478 486 481
rect 778 478 806 481
rect 818 478 822 481
rect 914 478 966 481
rect 1150 481 1153 488
rect 1670 482 1673 488
rect 1150 478 1206 481
rect 1210 478 1217 481
rect 1698 478 1742 481
rect 1770 478 1777 481
rect 1994 478 2014 481
rect 2058 478 2070 481
rect 2578 478 2670 481
rect 2682 478 2838 481
rect 2842 478 3110 481
rect 3290 478 3310 481
rect 3314 478 3545 481
rect 3554 478 3734 481
rect 3738 478 3990 481
rect 3994 478 4030 481
rect 4034 478 4046 481
rect 4050 478 4166 481
rect 4170 478 4350 481
rect 4354 478 4358 481
rect 4362 478 4374 481
rect 4522 478 4534 481
rect 4538 478 4870 481
rect 4890 478 4894 481
rect 4930 478 4934 481
rect 4990 478 5046 481
rect 5262 481 5265 488
rect 5210 478 5265 481
rect 550 472 553 478
rect 1270 472 1273 478
rect 122 468 166 471
rect 170 468 174 471
rect 330 468 374 471
rect 522 468 542 471
rect 674 468 678 471
rect 738 468 886 471
rect 890 468 1038 471
rect 1306 468 1414 471
rect 1486 471 1489 478
rect 1434 468 1489 471
rect 1634 468 1718 471
rect 1722 468 1790 471
rect 1870 471 1873 478
rect 1826 468 1873 471
rect 1902 472 1905 478
rect 1942 468 2006 471
rect 2058 468 2062 471
rect 2110 471 2113 478
rect 2074 468 2113 471
rect 2330 468 2334 471
rect 2366 471 2369 478
rect 2338 468 2414 471
rect 2510 468 2534 471
rect 2690 468 2702 471
rect 2722 468 2870 471
rect 2954 468 2974 471
rect 2994 468 3078 471
rect 3106 468 3166 471
rect 3170 468 3177 471
rect 3210 468 3246 471
rect 3250 468 3326 471
rect 3330 468 3342 471
rect 3542 471 3545 478
rect 3538 468 3545 471
rect 18 458 198 461
rect 298 458 302 461
rect 374 461 377 468
rect 374 458 398 461
rect 402 458 422 461
rect 494 461 497 468
rect 490 458 497 461
rect 530 459 590 461
rect 530 458 593 459
rect 690 458 774 461
rect 778 458 950 461
rect 986 458 1054 461
rect 1130 459 1190 461
rect 1942 462 1945 468
rect 1130 458 1193 459
rect 1306 458 1318 461
rect 1338 458 1409 461
rect 1698 458 1926 461
rect 1970 458 2022 461
rect 2026 458 2134 461
rect 2138 458 2158 461
rect 2294 461 2297 468
rect 2242 459 2297 461
rect 2238 458 2297 459
rect 2338 458 2358 461
rect 2510 461 2513 468
rect 2426 458 2513 461
rect 2522 458 2609 461
rect 2634 459 2694 461
rect 2630 458 2694 459
rect 2898 458 2926 461
rect 3010 458 3030 461
rect 3114 458 3214 461
rect 3358 461 3361 468
rect 3542 462 3545 468
rect 3562 468 3702 471
rect 3714 468 3718 471
rect 3866 468 3894 471
rect 3898 468 3902 471
rect 3914 468 3934 471
rect 3978 468 3982 471
rect 4154 468 4174 471
rect 4202 468 4206 471
rect 4250 468 4334 471
rect 4386 468 4406 471
rect 4410 468 4574 471
rect 4690 468 4718 471
rect 4722 468 4750 471
rect 4958 471 4961 478
rect 4834 468 4961 471
rect 4990 472 4993 478
rect 5270 472 5273 478
rect 5030 468 5070 471
rect 5106 468 5222 471
rect 3550 462 3553 468
rect 3282 458 3382 461
rect 3474 458 3478 461
rect 3554 458 3566 461
rect 3658 458 3742 461
rect 3826 458 3830 461
rect 4102 461 4105 468
rect 4018 458 4105 461
rect 4122 458 4214 461
rect 4366 461 4369 468
rect 4298 459 4369 461
rect 4294 458 4369 459
rect 4394 458 4398 461
rect 4498 458 4566 461
rect 4834 458 4838 461
rect 4874 458 5014 461
rect 5030 461 5033 468
rect 5018 458 5033 461
rect 5042 458 5046 461
rect 5050 458 5054 461
rect 5074 458 5126 461
rect 5130 458 5166 461
rect 5186 458 5201 461
rect 5234 458 5278 461
rect 154 448 182 451
rect 202 448 406 451
rect 554 448 742 451
rect 754 448 806 451
rect 810 448 942 451
rect 954 448 998 451
rect 1302 451 1305 458
rect 1106 448 1305 451
rect 1406 452 1409 458
rect 2606 452 2609 458
rect 2782 452 2785 458
rect 3526 452 3529 458
rect 1666 448 1670 451
rect 1778 448 1862 451
rect 1898 448 1982 451
rect 2090 448 2142 451
rect 2282 448 2334 451
rect 2426 448 2433 451
rect 18 438 382 441
rect 386 438 390 441
rect 770 438 830 441
rect 946 438 1294 441
rect 1298 438 1302 441
rect 1570 438 1854 441
rect 1862 441 1865 448
rect 2430 442 2433 448
rect 2466 448 2526 451
rect 2610 448 2742 451
rect 2746 448 2766 451
rect 2838 448 2857 451
rect 1862 438 1918 441
rect 1954 438 2070 441
rect 2110 438 2286 441
rect 2290 438 2398 441
rect 2446 441 2449 448
rect 2838 442 2841 448
rect 2854 442 2857 448
rect 2914 448 3182 451
rect 3266 448 3294 451
rect 3354 448 3361 451
rect 3386 448 3526 451
rect 3546 448 3566 451
rect 3610 448 3686 451
rect 3706 448 3742 451
rect 3746 448 3774 451
rect 3786 448 3822 451
rect 3930 448 3942 451
rect 4186 448 4198 451
rect 4410 448 4494 451
rect 4498 448 4518 451
rect 4522 448 4529 451
rect 4538 448 4654 451
rect 4658 448 4678 451
rect 4682 448 4734 451
rect 4738 448 4758 451
rect 4762 448 4774 451
rect 4790 451 4793 458
rect 5198 452 5201 458
rect 4790 448 4894 451
rect 4962 448 4966 451
rect 4978 448 5006 451
rect 5082 448 5105 451
rect 2870 442 2873 448
rect 3358 442 3361 448
rect 2446 438 2470 441
rect 2562 438 2566 441
rect 2570 438 2814 441
rect 3018 438 3022 441
rect 3034 438 3110 441
rect 3114 438 3326 441
rect 3582 441 3585 448
rect 5102 442 5105 448
rect 3530 438 3585 441
rect 3602 438 3710 441
rect 4170 438 4686 441
rect 178 428 198 431
rect 882 428 1014 431
rect 1066 428 1374 431
rect 1538 428 1614 431
rect 1666 428 1918 431
rect 1922 428 1942 431
rect 2110 431 2113 438
rect 1946 428 2113 431
rect 2122 428 2142 431
rect 2474 428 2518 431
rect 2882 428 3118 431
rect 3122 428 3158 431
rect 3534 428 3694 431
rect 3762 428 3982 431
rect 4026 428 4126 431
rect 4130 428 4270 431
rect 4442 428 4542 431
rect 4626 428 4750 431
rect 770 418 942 421
rect 962 418 982 421
rect 1322 418 1662 421
rect 1786 418 2070 421
rect 2106 418 3278 421
rect 3326 421 3329 428
rect 3534 422 3537 428
rect 3326 418 3470 421
rect 3666 418 4022 421
rect 4034 418 4166 421
rect 4170 418 4598 421
rect 4690 418 4710 421
rect 4714 418 4878 421
rect 4882 418 4982 421
rect 5146 418 5198 421
rect 394 408 1214 411
rect 1610 408 1806 411
rect 1882 408 1958 411
rect 2114 408 2166 411
rect 2178 408 2206 411
rect 3530 408 3534 411
rect 3714 408 3774 411
rect 3874 408 4038 411
rect 4106 408 4190 411
rect 5146 408 5158 411
rect 328 403 330 407
rect 334 403 337 407
rect 342 403 344 407
rect 1352 403 1354 407
rect 1358 403 1361 407
rect 1366 403 1368 407
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2398 403 2400 407
rect 3400 403 3402 407
rect 3406 403 3409 407
rect 3414 403 3416 407
rect 4424 403 4426 407
rect 4430 403 4433 407
rect 4438 403 4440 407
rect 690 398 902 401
rect 938 398 1246 401
rect 1258 398 1342 401
rect 1642 398 1734 401
rect 1738 398 1766 401
rect 1866 398 2038 401
rect 2722 398 2758 401
rect 2962 398 2990 401
rect 3042 398 3134 401
rect 3442 398 3486 401
rect 3490 398 3662 401
rect 3690 398 3798 401
rect 3802 398 3934 401
rect 3938 398 4038 401
rect 4042 398 4182 401
rect 4602 398 4718 401
rect 5138 398 5238 401
rect 550 392 553 398
rect 5286 392 5289 398
rect 754 388 758 391
rect 810 388 838 391
rect 1306 388 1382 391
rect 1674 388 1854 391
rect 1858 388 1918 391
rect 1922 388 2702 391
rect 2874 388 3238 391
rect 3258 388 3262 391
rect 3266 388 3326 391
rect 3394 388 3598 391
rect 3610 388 3734 391
rect 4042 388 4142 391
rect 4242 388 4406 391
rect 4410 388 4646 391
rect 5170 388 5190 391
rect 418 378 678 381
rect 730 378 753 381
rect 1378 378 1438 381
rect 1442 378 1510 381
rect 1514 378 1702 381
rect 1706 378 1782 381
rect 1794 378 1950 381
rect 2042 378 2094 381
rect 2154 378 2614 381
rect 2658 378 2702 381
rect 3050 378 3054 381
rect 3346 378 3558 381
rect 3722 378 3790 381
rect 4050 378 4054 381
rect 4058 378 4166 381
rect 4578 378 4886 381
rect 4890 378 4910 381
rect 4914 378 5161 381
rect 5170 378 5198 381
rect 750 372 753 378
rect 354 368 406 371
rect 442 368 654 371
rect 762 368 910 371
rect 914 368 1278 371
rect 1386 368 1470 371
rect 1626 368 1830 371
rect 1978 368 2086 371
rect 2130 368 2174 371
rect 2178 368 2214 371
rect 2346 368 2398 371
rect 2850 368 3062 371
rect 3218 368 3494 371
rect 3738 368 3758 371
rect 3770 368 3886 371
rect 4034 368 4046 371
rect 4258 368 4342 371
rect 4642 368 4782 371
rect 4786 368 4990 371
rect 4994 368 5014 371
rect 5158 371 5161 378
rect 5158 368 5254 371
rect 5258 368 5262 371
rect 210 358 214 361
rect 258 358 406 361
rect 410 358 454 361
rect 458 358 798 361
rect 826 358 1006 361
rect 1018 358 1206 361
rect 1334 361 1337 368
rect 1350 361 1353 368
rect 2246 362 2249 368
rect 2702 362 2705 368
rect 1334 358 1353 361
rect 1538 358 1542 361
rect 1794 358 1814 361
rect 1882 358 1926 361
rect 2018 358 2182 361
rect 2266 358 2310 361
rect 2362 358 2382 361
rect 2418 358 2430 361
rect 2434 358 2462 361
rect 2818 358 2942 361
rect 3042 358 3158 361
rect 3514 358 3622 361
rect 3706 358 3726 361
rect 3746 358 3769 361
rect 3810 358 3814 361
rect 3986 358 4078 361
rect 4130 358 4206 361
rect 4246 361 4249 368
rect 4210 358 4249 361
rect 4394 358 4454 361
rect 4586 358 4878 361
rect 4882 358 4910 361
rect 5186 358 5190 361
rect 10 348 14 351
rect 226 348 326 351
rect 330 348 334 351
rect 1006 351 1009 358
rect 474 348 585 351
rect 86 341 89 348
rect 582 342 585 348
rect 710 348 817 351
rect 1006 348 1118 351
rect 1194 348 1222 351
rect 1226 348 1254 351
rect 1414 351 1417 358
rect 1330 348 1417 351
rect 1530 348 1542 351
rect 1594 348 1598 351
rect 1702 351 1705 358
rect 1650 348 1705 351
rect 1758 348 1809 351
rect 1818 348 1894 351
rect 1914 348 1982 351
rect 2122 348 2134 351
rect 2218 348 2286 351
rect 2378 348 2446 351
rect 2450 348 2590 351
rect 2594 348 2638 351
rect 2642 348 2726 351
rect 3050 348 3190 351
rect 3206 351 3209 358
rect 3766 352 3769 358
rect 3838 352 3841 358
rect 3206 348 3222 351
rect 3306 348 3382 351
rect 3546 348 3550 351
rect 3578 348 3582 351
rect 3626 348 3662 351
rect 3706 348 3750 351
rect 3930 348 4030 351
rect 4102 351 4105 358
rect 4102 348 4158 351
rect 4186 348 4198 351
rect 4286 351 4289 358
rect 4234 348 4289 351
rect 4362 348 4398 351
rect 4594 348 4638 351
rect 4682 348 4686 351
rect 4706 348 4710 351
rect 4722 348 4742 351
rect 4814 348 4902 351
rect 5002 348 5070 351
rect 5074 348 5081 351
rect 5154 348 5246 351
rect 710 342 713 348
rect 814 342 817 348
rect 1310 342 1313 348
rect 66 338 89 341
rect 202 338 206 341
rect 250 338 310 341
rect 370 338 398 341
rect 402 338 454 341
rect 818 338 926 341
rect 994 338 1078 341
rect 1122 338 1206 341
rect 1314 338 1326 341
rect 1354 338 1614 341
rect 1758 341 1761 348
rect 1618 338 1761 341
rect 1770 338 1782 341
rect 1806 341 1809 348
rect 2038 342 2041 348
rect 2094 342 2097 348
rect 2134 342 2137 348
rect 1806 338 1822 341
rect 1938 338 1966 341
rect 2058 338 2062 341
rect 2234 338 2262 341
rect 2314 338 2398 341
rect 2402 338 2406 341
rect 2458 338 2542 341
rect 2618 338 2630 341
rect 2634 338 2670 341
rect 2690 338 2758 341
rect 2902 341 2905 348
rect 4814 342 4817 348
rect 2770 338 2905 341
rect 2986 338 2998 341
rect 3050 338 3070 341
rect 3202 338 3294 341
rect 3302 338 3366 341
rect 3650 338 3654 341
rect 3714 338 3766 341
rect 3834 338 3846 341
rect 3890 338 4137 341
rect 4178 338 4182 341
rect 4226 338 4350 341
rect 4698 338 4750 341
rect 4978 338 4982 341
rect 5010 338 5014 341
rect 5170 338 5222 341
rect 5266 338 5278 341
rect 1798 332 1801 338
rect 266 328 310 331
rect 314 328 318 331
rect 642 328 1014 331
rect 1250 328 1342 331
rect 1510 328 1542 331
rect 1570 328 1574 331
rect 1846 328 1870 331
rect 2002 328 2030 331
rect 2034 328 2041 331
rect 2050 328 2062 331
rect 2158 331 2161 338
rect 2066 328 2161 331
rect 2218 328 2246 331
rect 2274 328 2286 331
rect 2322 328 2598 331
rect 2658 328 2662 331
rect 2670 331 2673 338
rect 3302 332 3305 338
rect 4134 332 4137 338
rect 2670 328 2694 331
rect 2866 328 3006 331
rect 3162 328 3302 331
rect 3394 328 3574 331
rect 3650 328 3686 331
rect 3746 328 3782 331
rect 3826 328 3830 331
rect 3898 328 4022 331
rect 4138 328 4182 331
rect 4490 328 4502 331
rect 4506 328 4790 331
rect 4874 328 4942 331
rect 4970 328 5134 331
rect 5162 328 5182 331
rect 5218 328 5294 331
rect 42 318 254 321
rect 366 321 369 328
rect 1510 322 1513 328
rect 1582 322 1585 328
rect 266 318 369 321
rect 506 318 649 321
rect 890 318 950 321
rect 994 318 1126 321
rect 1130 318 1334 321
rect 1846 321 1849 328
rect 1802 318 1849 321
rect 1858 318 2022 321
rect 2086 318 2094 321
rect 2098 318 2190 321
rect 2630 321 2633 328
rect 2386 318 2633 321
rect 2882 318 3030 321
rect 3474 318 3614 321
rect 3618 318 3678 321
rect 3754 318 3878 321
rect 4378 318 4510 321
rect 4546 318 4654 321
rect 4658 318 4734 321
rect 4770 318 4926 321
rect 4930 318 4950 321
rect 4962 318 5238 321
rect 5242 318 5270 321
rect 646 312 649 318
rect 5278 312 5281 318
rect 10 308 70 311
rect 74 308 94 311
rect 98 308 358 311
rect 370 308 486 311
rect 930 308 1094 311
rect 1474 308 1670 311
rect 1746 308 1750 311
rect 1922 308 2126 311
rect 2362 308 2422 311
rect 2442 308 2678 311
rect 2682 308 2846 311
rect 3090 308 3102 311
rect 3826 308 3886 311
rect 4114 308 4198 311
rect 4586 308 4662 311
rect 4682 308 4702 311
rect 5210 308 5214 311
rect 5234 308 5238 311
rect 848 303 850 307
rect 854 303 857 307
rect 862 303 864 307
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1886 303 1888 307
rect 2888 303 2890 307
rect 2894 303 2897 307
rect 2902 303 2904 307
rect 3920 303 3922 307
rect 3926 303 3929 307
rect 3934 303 3936 307
rect 4936 303 4938 307
rect 4942 303 4945 307
rect 4950 303 4952 307
rect 114 298 166 301
rect 170 298 286 301
rect 802 298 822 301
rect 954 298 982 301
rect 1074 298 1206 301
rect 1442 298 1518 301
rect 1538 298 1622 301
rect 1626 298 1774 301
rect 2002 298 2102 301
rect 2106 298 2126 301
rect 2154 298 2182 301
rect 2482 298 2830 301
rect 2834 298 2838 301
rect 2842 298 2862 301
rect 2962 298 3022 301
rect 3026 298 3054 301
rect 3066 298 3246 301
rect 3314 298 3438 301
rect 3442 298 3598 301
rect 3626 298 3678 301
rect 3682 298 3758 301
rect 3762 298 3862 301
rect 4650 298 4806 301
rect 5146 298 5246 301
rect 5250 298 5286 301
rect 26 288 190 291
rect 202 288 214 291
rect 218 288 382 291
rect 410 288 438 291
rect 754 288 958 291
rect 1050 288 1070 291
rect 1218 288 1278 291
rect 1298 288 1430 291
rect 1498 288 1526 291
rect 1530 288 1582 291
rect 1730 288 1769 291
rect 1786 288 1838 291
rect 1842 288 2158 291
rect 2250 288 2454 291
rect 2650 288 2710 291
rect 2938 288 3214 291
rect 3266 288 3278 291
rect 3282 288 3294 291
rect 3858 288 3913 291
rect 4026 288 4054 291
rect 4146 288 4230 291
rect 4338 288 4366 291
rect 4370 288 4398 291
rect 4402 288 4518 291
rect 4522 288 4542 291
rect 5002 288 5006 291
rect 5042 288 5094 291
rect 5098 288 5126 291
rect 5210 288 5214 291
rect 162 278 302 281
rect 306 278 350 281
rect 354 278 446 281
rect 450 278 606 281
rect 610 278 638 281
rect 882 278 886 281
rect 890 278 918 281
rect 1210 278 1382 281
rect 1386 278 1398 281
rect 1590 281 1593 288
rect 1766 282 1769 288
rect 1482 278 1593 281
rect 1666 278 1742 281
rect 1770 278 1806 281
rect 2170 278 2230 281
rect 2638 281 2641 288
rect 2490 278 2641 281
rect 2826 278 2849 281
rect 346 268 422 271
rect 458 268 486 271
rect 662 271 665 278
rect 806 272 809 278
rect 570 268 665 271
rect 690 268 774 271
rect 826 268 862 271
rect 866 268 878 271
rect 1042 268 1094 271
rect 1178 268 1238 271
rect 1242 268 1278 271
rect 1282 268 1310 271
rect 1338 268 1457 271
rect 1490 268 1542 271
rect 1730 268 1766 271
rect 1962 268 1966 271
rect 1986 268 2014 271
rect 2018 268 2110 271
rect 2302 271 2305 278
rect 2846 272 2849 278
rect 2926 281 2929 288
rect 3710 282 3713 288
rect 3910 282 3913 288
rect 2926 278 2990 281
rect 3074 278 3110 281
rect 3122 278 3222 281
rect 3226 278 3318 281
rect 3322 278 3342 281
rect 3482 278 3486 281
rect 3666 278 3670 281
rect 3794 278 3830 281
rect 4354 278 4382 281
rect 4538 278 4542 281
rect 4630 278 4670 281
rect 4674 278 4718 281
rect 4758 281 4761 288
rect 5246 282 5249 288
rect 4758 278 4782 281
rect 4930 278 4990 281
rect 4994 278 5142 281
rect 5146 278 5150 281
rect 5218 278 5222 281
rect 5282 278 5286 281
rect 2918 272 2921 278
rect 2302 268 2422 271
rect 2426 268 2470 271
rect 2530 268 2606 271
rect 2674 268 2678 271
rect 2722 268 2734 271
rect 2922 268 2942 271
rect 3026 268 3158 271
rect 3258 268 3278 271
rect 3518 271 3521 278
rect 4630 272 4633 278
rect 3386 268 3521 271
rect 3530 268 3534 271
rect 3570 268 3777 271
rect 3802 268 3838 271
rect 4002 268 4174 271
rect 4182 268 4209 271
rect 4218 268 4494 271
rect 4498 268 4582 271
rect 4746 268 4846 271
rect 4906 268 4926 271
rect 4978 268 5166 271
rect 5242 268 5254 271
rect 5282 268 5302 271
rect 142 262 145 268
rect 254 262 257 268
rect 290 258 390 261
rect 438 261 441 268
rect 1454 262 1457 268
rect 438 258 534 261
rect 538 258 686 261
rect 802 258 822 261
rect 1050 258 1078 261
rect 1082 258 1134 261
rect 1138 258 1302 261
rect 1310 258 1377 261
rect 1586 258 1598 261
rect 1602 258 1742 261
rect 2010 258 2065 261
rect 2222 261 2225 268
rect 2630 262 2633 268
rect 2154 258 2225 261
rect 2234 258 2254 261
rect 2282 258 2318 261
rect 2594 258 2614 261
rect 2662 258 2694 261
rect 2698 258 2718 261
rect 2730 258 2902 261
rect 2906 258 3174 261
rect 3186 258 3342 261
rect 3346 258 3478 261
rect 3482 258 3502 261
rect 3506 258 3742 261
rect 3774 261 3777 268
rect 3774 258 3806 261
rect 3882 258 3958 261
rect 4018 258 4046 261
rect 4182 261 4185 268
rect 4206 262 4209 268
rect 4162 258 4185 261
rect 4194 258 4198 261
rect 4218 258 4310 261
rect 4570 258 4606 261
rect 4698 258 4718 261
rect 4834 258 4902 261
rect 5002 258 5006 261
rect 5018 258 5022 261
rect 5066 258 5182 261
rect 5226 258 5286 261
rect 1310 252 1313 258
rect 1374 252 1377 258
rect 2062 252 2065 258
rect 66 248 214 251
rect 218 248 414 251
rect 426 248 454 251
rect 458 248 638 251
rect 650 248 942 251
rect 1170 248 1214 251
rect 1218 248 1286 251
rect 1522 248 1638 251
rect 1786 248 1806 251
rect 2178 248 2214 251
rect 2218 248 2246 251
rect 2338 248 2598 251
rect 2662 251 2665 258
rect 2602 248 2665 251
rect 2670 248 2678 251
rect 2702 248 2710 251
rect 2714 248 2774 251
rect 2890 248 3086 251
rect 3110 248 3118 251
rect 3122 248 3182 251
rect 3210 248 3222 251
rect 3258 248 3265 251
rect 602 238 894 241
rect 1026 238 1086 241
rect 1090 238 1110 241
rect 1114 238 1494 241
rect 1538 238 1670 241
rect 1834 238 2062 241
rect 2618 238 3022 241
rect 3086 241 3089 248
rect 3262 242 3265 248
rect 3334 248 3374 251
rect 3578 248 3694 251
rect 3782 248 3790 251
rect 4042 248 4102 251
rect 4174 248 4246 251
rect 4282 248 4366 251
rect 4422 251 4425 258
rect 4402 248 4534 251
rect 4570 248 4590 251
rect 4778 248 4782 251
rect 4786 248 4974 251
rect 5010 248 5070 251
rect 3334 242 3337 248
rect 3782 242 3785 248
rect 4174 242 4177 248
rect 3086 238 3118 241
rect 3386 238 3670 241
rect 3706 238 3750 241
rect 3818 238 4054 241
rect 4226 238 4294 241
rect 4546 238 4774 241
rect 1570 228 2126 231
rect 2482 228 2830 231
rect 2946 228 3230 231
rect 3458 228 3654 231
rect 4050 228 4510 231
rect 4530 228 4550 231
rect 4554 228 4806 231
rect 4810 228 5062 231
rect 722 218 1038 221
rect 1106 218 1566 221
rect 1578 218 1630 221
rect 1634 218 1670 221
rect 1674 218 1678 221
rect 1682 218 1910 221
rect 1914 218 2062 221
rect 2650 218 2918 221
rect 3010 218 3094 221
rect 3146 218 3425 221
rect 3554 218 3646 221
rect 3650 218 3726 221
rect 3730 218 3862 221
rect 3866 218 3902 221
rect 4386 218 4414 221
rect 4418 218 4430 221
rect 4810 218 4830 221
rect 4994 218 5086 221
rect 5090 218 5222 221
rect 1698 208 1790 211
rect 1890 208 2030 211
rect 2034 208 2102 211
rect 2114 208 2334 211
rect 2466 208 2870 211
rect 2918 211 2921 218
rect 2918 208 3214 211
rect 3422 211 3425 218
rect 3422 208 3622 211
rect 3898 208 3902 211
rect 4210 208 4406 211
rect 4658 208 5142 211
rect 328 203 330 207
rect 334 203 337 207
rect 342 203 344 207
rect 1352 203 1354 207
rect 1358 203 1361 207
rect 1366 203 1368 207
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2398 203 2400 207
rect 3400 203 3402 207
rect 3406 203 3409 207
rect 3414 203 3416 207
rect 3654 202 3657 208
rect 4424 203 4426 207
rect 4430 203 4433 207
rect 4438 203 4440 207
rect 1682 198 1982 201
rect 2634 198 2854 201
rect 2858 198 2894 201
rect 2898 198 3062 201
rect 3282 198 3390 201
rect 4082 198 4406 201
rect 5026 198 5198 201
rect 210 188 238 191
rect 1322 188 1665 191
rect 1978 188 1998 191
rect 2066 188 2662 191
rect 3162 188 3166 191
rect 3170 188 3462 191
rect 3498 188 3694 191
rect 3754 188 3766 191
rect 4146 188 4582 191
rect 5002 188 5062 191
rect 5082 188 5086 191
rect 1322 178 1582 181
rect 1662 181 1665 188
rect 1662 178 1702 181
rect 1706 178 1774 181
rect 1778 178 2270 181
rect 2274 178 2358 181
rect 2370 178 2401 181
rect 2834 178 3006 181
rect 3266 178 3734 181
rect 4058 178 4590 181
rect 4594 178 4686 181
rect 4930 178 5158 181
rect 5230 181 5233 188
rect 5162 178 5233 181
rect 2398 172 2401 178
rect 274 168 294 171
rect 698 168 718 171
rect 722 168 838 171
rect 842 168 1102 171
rect 1226 168 1326 171
rect 1466 168 1534 171
rect 1746 168 1894 171
rect 1978 168 2046 171
rect 2050 168 2094 171
rect 2098 168 2198 171
rect 2202 168 2398 171
rect 2730 168 2846 171
rect 3226 168 3318 171
rect 3426 168 3478 171
rect 3586 168 3678 171
rect 3682 168 3838 171
rect 4002 168 4126 171
rect 4366 168 4374 171
rect 4378 168 4414 171
rect 4450 168 4478 171
rect 4578 168 4598 171
rect 4602 168 4638 171
rect 4706 168 4718 171
rect 4722 168 4766 171
rect 4786 168 4990 171
rect 5018 168 5030 171
rect 5230 162 5233 168
rect 434 158 462 161
rect 1018 158 1278 161
rect 1346 158 1510 161
rect 2106 158 2310 161
rect 2818 158 2862 161
rect 3234 158 3334 161
rect 3474 158 3606 161
rect 3614 158 3654 161
rect 3826 158 3926 161
rect 4066 158 4102 161
rect 4122 158 4518 161
rect 4554 158 4710 161
rect 4754 158 4814 161
rect 4986 158 5030 161
rect 102 151 105 158
rect 90 148 105 151
rect 170 148 302 151
rect 306 148 390 151
rect 410 148 438 151
rect 442 148 550 151
rect 554 148 566 151
rect 634 148 662 151
rect 886 151 889 158
rect 886 148 902 151
rect 1034 148 1062 151
rect 1242 148 1246 151
rect 1474 148 1494 151
rect 1658 148 1686 151
rect 14 142 17 148
rect 1238 142 1241 148
rect 1770 148 1774 151
rect 1830 151 1833 158
rect 1818 148 1833 151
rect 1850 148 1854 151
rect 1942 151 1945 158
rect 1914 148 1945 151
rect 2038 151 2041 158
rect 2026 148 2041 151
rect 2090 148 2118 151
rect 2134 148 2150 151
rect 2242 148 2262 151
rect 2266 148 2286 151
rect 2338 148 2358 151
rect 2626 148 2638 151
rect 2654 151 2657 158
rect 2642 148 2657 151
rect 2666 148 2670 151
rect 2850 148 2934 151
rect 2986 148 2990 151
rect 3070 151 3073 158
rect 3058 148 3073 151
rect 3086 152 3089 158
rect 3110 152 3113 158
rect 3098 148 3102 151
rect 3218 148 3430 151
rect 3434 148 3462 151
rect 3490 148 3494 151
rect 3498 148 3518 151
rect 3614 151 3617 158
rect 3530 148 3617 151
rect 3650 148 3870 151
rect 4110 151 4113 158
rect 3922 148 4113 151
rect 4218 148 4270 151
rect 4306 148 4694 151
rect 4754 148 4758 151
rect 5038 151 5041 158
rect 5246 152 5249 158
rect 4882 148 5041 151
rect 5074 148 5126 151
rect 5274 148 5278 151
rect 2134 142 2137 148
rect 154 138 185 141
rect 394 138 446 141
rect 450 138 734 141
rect 738 138 1014 141
rect 1082 138 1182 141
rect 1186 138 1238 141
rect 1242 138 1358 141
rect 1362 138 1822 141
rect 2034 138 2134 141
rect 2194 138 2430 141
rect 2442 138 2518 141
rect 2542 141 2545 148
rect 2522 138 2545 141
rect 2570 138 2662 141
rect 2714 138 2742 141
rect 2754 138 2878 141
rect 2930 138 2934 141
rect 3066 138 3110 141
rect 3114 138 3158 141
rect 3178 138 3238 141
rect 3418 138 3462 141
rect 3610 138 3622 141
rect 3650 138 3654 141
rect 3690 138 3702 141
rect 3874 138 3918 141
rect 3978 138 3982 141
rect 4034 138 4054 141
rect 4074 138 4078 141
rect 4290 138 4310 141
rect 4314 138 4318 141
rect 4322 138 4638 141
rect 4738 138 4766 141
rect 4770 138 5022 141
rect 5114 138 5177 141
rect 182 132 185 138
rect 5174 132 5177 138
rect 5262 132 5265 138
rect 546 128 670 131
rect 962 128 1038 131
rect 1066 128 1078 131
rect 1402 128 1486 131
rect 1522 128 1534 131
rect 1586 128 1662 131
rect 1794 128 1926 131
rect 1934 128 2078 131
rect 2090 128 2318 131
rect 2370 128 2694 131
rect 2698 128 2718 131
rect 2890 128 3526 131
rect 3538 128 3630 131
rect 3642 128 3686 131
rect 3954 128 4041 131
rect 4370 128 4614 131
rect 4770 128 4870 131
rect 4890 128 4894 131
rect 458 118 518 121
rect 522 118 550 121
rect 602 118 606 121
rect 706 118 726 121
rect 834 118 838 121
rect 954 118 1078 121
rect 1082 118 1118 121
rect 1122 118 1254 121
rect 1258 118 1374 121
rect 1378 118 1486 121
rect 1934 121 1937 128
rect 1690 118 1937 121
rect 2350 121 2353 128
rect 1954 118 2353 121
rect 2786 118 2910 121
rect 2914 118 3566 121
rect 3886 121 3889 128
rect 3578 118 3889 121
rect 4038 122 4041 128
rect 4330 118 4598 121
rect 4790 118 4950 121
rect 58 108 542 111
rect 1018 108 1222 111
rect 1714 108 1806 111
rect 1898 108 2014 111
rect 2066 108 2286 111
rect 2306 108 2710 111
rect 3018 108 3454 111
rect 3466 108 3710 111
rect 3946 108 4150 111
rect 4250 108 4294 111
rect 4410 108 4430 111
rect 4790 111 4793 118
rect 4442 108 4793 111
rect 848 103 850 107
rect 854 103 857 107
rect 862 103 864 107
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1886 103 1888 107
rect 2888 103 2890 107
rect 2894 103 2897 107
rect 2902 103 2904 107
rect 3920 103 3922 107
rect 3926 103 3929 107
rect 3934 103 3936 107
rect 4798 102 4801 108
rect 4936 103 4938 107
rect 4942 103 4945 107
rect 4950 103 4952 107
rect 178 98 198 101
rect 202 98 222 101
rect 426 98 446 101
rect 450 98 710 101
rect 1010 98 1062 101
rect 1218 98 1462 101
rect 1570 98 1646 101
rect 2010 98 2086 101
rect 2154 98 2494 101
rect 2498 98 2646 101
rect 2650 98 2702 101
rect 2914 98 2926 101
rect 3114 98 3142 101
rect 3362 98 3534 101
rect 3538 98 3590 101
rect 3610 98 3870 101
rect 3946 98 4174 101
rect 4186 98 4254 101
rect 4338 98 4486 101
rect 18 88 102 91
rect 218 88 302 91
rect 306 88 446 91
rect 1274 88 1310 91
rect 1426 88 1798 91
rect 1866 88 1894 91
rect 1922 88 2094 91
rect 2114 88 2254 91
rect 2894 88 2918 91
rect 3130 88 3230 91
rect 3234 88 3382 91
rect 3394 88 3438 91
rect 3466 88 3470 91
rect 3490 88 3494 91
rect 3546 88 3574 91
rect 3626 88 3710 91
rect 3778 88 3854 91
rect 3858 88 3862 91
rect 3906 88 3942 91
rect 4018 88 4054 91
rect 4122 88 4126 91
rect 4250 88 4286 91
rect 4290 88 4374 91
rect 4418 88 4566 91
rect 4626 88 4782 91
rect 4834 88 4838 91
rect 4882 88 4934 91
rect 74 78 126 81
rect 562 78 662 81
rect 802 78 926 81
rect 1030 81 1033 88
rect 970 78 1033 81
rect 1114 78 1206 81
rect 1350 81 1353 88
rect 1350 78 1374 81
rect 1422 81 1425 88
rect 1386 78 1425 81
rect 1626 78 1670 81
rect 1674 78 1702 81
rect 1910 81 1913 88
rect 2894 82 2897 88
rect 1910 78 1974 81
rect 1982 78 2054 81
rect 2418 78 2518 81
rect 2746 78 2886 81
rect 3058 78 3134 81
rect 3202 78 3310 81
rect 3434 78 3494 81
rect 3506 78 3582 81
rect 3586 78 3606 81
rect 3690 78 3838 81
rect 3842 78 3966 81
rect 4098 78 4126 81
rect 4130 78 4262 81
rect 4266 78 4302 81
rect 4390 78 4398 81
rect 4402 78 4438 81
rect 4458 78 4526 81
rect 4594 78 4750 81
rect 4754 78 4790 81
rect 4826 78 4830 81
rect 4914 78 4918 81
rect 5034 78 5038 81
rect 122 68 150 71
rect 154 68 686 71
rect 722 68 814 71
rect 818 68 846 71
rect 882 68 894 71
rect 914 68 1046 71
rect 1106 68 1326 71
rect 1330 68 1542 71
rect 1650 68 1678 71
rect 1982 71 1985 78
rect 1818 68 1985 71
rect 2034 68 2118 71
rect 2562 68 2574 71
rect 2578 68 2646 71
rect 2746 68 2838 71
rect 2842 68 2958 71
rect 3030 71 3033 78
rect 2962 68 3033 71
rect 3186 68 3230 71
rect 3322 68 3430 71
rect 3434 68 3438 71
rect 3558 68 3622 71
rect 3738 68 3742 71
rect 3746 68 3758 71
rect 3898 68 3910 71
rect 3914 68 3918 71
rect 4030 71 4033 78
rect 4446 72 4449 78
rect 4030 68 4206 71
rect 4210 68 4289 71
rect 4410 68 4422 71
rect 4490 68 4550 71
rect 4642 68 5102 71
rect 5214 71 5217 78
rect 5146 68 5217 71
rect 5234 68 5286 71
rect 138 58 166 61
rect 194 58 249 61
rect 378 58 414 61
rect 634 58 638 61
rect 682 58 1014 61
rect 1026 58 1038 61
rect 1178 58 1193 61
rect 1242 59 1262 61
rect 1242 58 1265 59
rect 1418 58 1630 61
rect 1750 61 1753 68
rect 1750 58 1918 61
rect 2142 61 2145 68
rect 2142 58 2158 61
rect 2326 61 2329 68
rect 2326 58 2374 61
rect 2502 61 2505 68
rect 3558 62 3561 68
rect 4286 62 4289 68
rect 2490 58 2505 61
rect 2546 58 2550 61
rect 2570 58 2646 61
rect 2730 58 2734 61
rect 2826 58 2830 61
rect 2898 58 2934 61
rect 2962 58 2966 61
rect 3218 58 3254 61
rect 3314 58 3534 61
rect 3570 58 3582 61
rect 3610 58 3734 61
rect 3738 58 3886 61
rect 3890 58 4070 61
rect 4074 58 4150 61
rect 4250 58 4254 61
rect 4386 58 4414 61
rect 4426 58 4622 61
rect 4650 58 4710 61
rect 4730 58 4790 61
rect 4890 59 4958 61
rect 4886 58 4958 59
rect 5002 59 5126 61
rect 4998 58 5126 59
rect 5170 58 5174 61
rect 246 52 249 58
rect 1190 52 1193 58
rect 634 48 646 51
rect 786 48 894 51
rect 1194 48 1334 51
rect 1398 51 1401 58
rect 1398 48 1494 51
rect 2126 51 2129 58
rect 2126 48 2230 51
rect 3598 51 3601 58
rect 3598 48 3654 51
rect 3750 48 3806 51
rect 4098 48 4454 51
rect 4770 48 4774 51
rect 5026 48 5174 51
rect 5178 48 5182 51
rect 5334 51 5338 52
rect 5202 48 5338 51
rect 3750 42 3753 48
rect 714 38 822 41
rect 826 38 1350 41
rect 4090 38 4606 41
rect 4610 38 4982 41
rect 2226 8 2230 11
rect 4530 8 4534 11
rect 328 3 330 7
rect 334 3 337 7
rect 342 3 344 7
rect 1352 3 1354 7
rect 1358 3 1361 7
rect 1366 3 1368 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2398 3 2400 7
rect 3400 3 3402 7
rect 3406 3 3409 7
rect 3414 3 3416 7
rect 4424 3 4426 7
rect 4430 3 4433 7
rect 4438 3 4440 7
<< m4contact >>
rect 850 5103 854 5107
rect 858 5103 861 5107
rect 861 5103 862 5107
rect 1874 5103 1878 5107
rect 1882 5103 1885 5107
rect 1885 5103 1886 5107
rect 2890 5103 2894 5107
rect 2898 5103 2901 5107
rect 2901 5103 2902 5107
rect 3922 5103 3926 5107
rect 3930 5103 3933 5107
rect 3933 5103 3934 5107
rect 4938 5103 4942 5107
rect 4946 5103 4949 5107
rect 4949 5103 4950 5107
rect 318 5098 322 5102
rect 1654 5098 1658 5102
rect 2750 5088 2754 5092
rect 1134 5078 1138 5082
rect 4486 5078 4490 5082
rect 4494 5078 4498 5082
rect 5206 5078 5210 5082
rect 310 5068 314 5072
rect 1534 5068 1538 5072
rect 5166 5068 5170 5072
rect 174 5058 178 5062
rect 206 5058 210 5062
rect 462 5058 466 5062
rect 566 5058 570 5062
rect 838 5058 842 5062
rect 1782 5058 1786 5062
rect 4078 5058 4082 5062
rect 4574 5058 4578 5062
rect 4902 5058 4906 5062
rect 4926 5058 4930 5062
rect 5238 5058 5242 5062
rect 3278 5048 3282 5052
rect 3558 5048 3562 5052
rect 3950 5048 3954 5052
rect 4910 5048 4914 5052
rect 806 5038 810 5042
rect 5014 5038 5018 5042
rect 366 5028 370 5032
rect 950 5028 954 5032
rect 2438 5018 2442 5022
rect 3686 5018 3690 5022
rect 4134 5018 4138 5022
rect 4526 5018 4530 5022
rect 5054 5018 5058 5022
rect 5150 5018 5154 5022
rect 926 5008 930 5012
rect 330 5003 334 5007
rect 338 5003 341 5007
rect 341 5003 342 5007
rect 1354 5003 1358 5007
rect 1362 5003 1365 5007
rect 1365 5003 1366 5007
rect 2386 5003 2390 5007
rect 2394 5003 2397 5007
rect 2397 5003 2398 5007
rect 3402 5003 3406 5007
rect 3410 5003 3413 5007
rect 3413 5003 3414 5007
rect 4426 5003 4430 5007
rect 4434 5003 4437 5007
rect 4437 5003 4438 5007
rect 1662 4998 1666 5002
rect 3558 4998 3562 5002
rect 3550 4988 3554 4992
rect 4190 4978 4194 4982
rect 286 4968 290 4972
rect 438 4968 442 4972
rect 726 4968 730 4972
rect 742 4968 746 4972
rect 4614 4968 4618 4972
rect 4758 4968 4762 4972
rect 5118 4968 5122 4972
rect 374 4958 378 4962
rect 422 4958 426 4962
rect 478 4958 482 4962
rect 486 4958 490 4962
rect 2222 4958 2226 4962
rect 2630 4958 2634 4962
rect 182 4948 186 4952
rect 214 4948 218 4952
rect 246 4948 250 4952
rect 758 4948 762 4952
rect 1454 4948 1458 4952
rect 1734 4948 1738 4952
rect 366 4938 370 4942
rect 774 4938 778 4942
rect 806 4938 810 4942
rect 3574 4948 3578 4952
rect 3590 4948 3594 4952
rect 3702 4948 3706 4952
rect 3726 4948 3730 4952
rect 4094 4948 4098 4952
rect 4526 4948 4530 4952
rect 4126 4938 4130 4942
rect 206 4928 210 4932
rect 486 4928 490 4932
rect 758 4928 762 4932
rect 4190 4938 4194 4942
rect 4910 4938 4914 4942
rect 5014 4938 5018 4942
rect 5126 4938 5130 4942
rect 3846 4928 3850 4932
rect 5006 4928 5010 4932
rect 5094 4928 5098 4932
rect 374 4918 378 4922
rect 606 4918 610 4922
rect 934 4918 938 4922
rect 2158 4918 2162 4922
rect 4134 4918 4138 4922
rect 4182 4918 4186 4922
rect 4862 4918 4866 4922
rect 5030 4918 5034 4922
rect 5086 4918 5090 4922
rect 5230 4918 5234 4922
rect 462 4908 466 4912
rect 3590 4908 3594 4912
rect 4286 4908 4290 4912
rect 850 4903 854 4907
rect 858 4903 861 4907
rect 861 4903 862 4907
rect 1874 4903 1878 4907
rect 1882 4903 1885 4907
rect 1885 4903 1886 4907
rect 2890 4903 2894 4907
rect 2898 4903 2901 4907
rect 2901 4903 2902 4907
rect 3922 4903 3926 4907
rect 3930 4903 3933 4907
rect 3933 4903 3934 4907
rect 4938 4903 4942 4907
rect 4946 4903 4949 4907
rect 4949 4903 4950 4907
rect 870 4898 874 4902
rect 1318 4898 1322 4902
rect 2102 4898 2106 4902
rect 2878 4898 2882 4902
rect 4678 4898 4682 4902
rect 182 4888 186 4892
rect 2582 4888 2586 4892
rect 4094 4888 4098 4892
rect 5046 4888 5050 4892
rect 5190 4888 5194 4892
rect 550 4878 554 4882
rect 710 4878 714 4882
rect 1046 4878 1050 4882
rect 2454 4878 2458 4882
rect 3430 4878 3434 4882
rect 5030 4878 5034 4882
rect 5246 4878 5250 4882
rect 5262 4878 5266 4882
rect 126 4868 130 4872
rect 950 4868 954 4872
rect 1022 4868 1026 4872
rect 1174 4868 1178 4872
rect 2406 4868 2410 4872
rect 2726 4868 2730 4872
rect 3526 4868 3530 4872
rect 4406 4868 4410 4872
rect 5070 4868 5074 4872
rect 5110 4868 5114 4872
rect 5254 4868 5258 4872
rect 38 4858 42 4862
rect 798 4858 802 4862
rect 878 4858 882 4862
rect 1078 4858 1082 4862
rect 1462 4858 1466 4862
rect 2182 4858 2186 4862
rect 4134 4858 4138 4862
rect 4606 4858 4610 4862
rect 5134 4858 5138 4862
rect 166 4848 170 4852
rect 742 4848 746 4852
rect 2558 4848 2562 4852
rect 3254 4848 3258 4852
rect 3582 4848 3586 4852
rect 214 4838 218 4842
rect 566 4838 570 4842
rect 2630 4838 2634 4842
rect 2926 4838 2930 4842
rect 4214 4848 4218 4852
rect 5070 4848 5074 4852
rect 5254 4848 5258 4852
rect 4534 4838 4538 4842
rect 5270 4838 5274 4842
rect 4126 4828 4130 4832
rect 246 4818 250 4822
rect 550 4818 554 4822
rect 2350 4818 2354 4822
rect 3422 4818 3426 4822
rect 4214 4818 4218 4822
rect 4726 4818 4730 4822
rect 5278 4818 5282 4822
rect 414 4808 418 4812
rect 2262 4808 2266 4812
rect 2438 4808 2442 4812
rect 2566 4808 2570 4812
rect 5006 4808 5010 4812
rect 5286 4808 5290 4812
rect 330 4803 334 4807
rect 338 4803 341 4807
rect 341 4803 342 4807
rect 1354 4803 1358 4807
rect 1362 4803 1365 4807
rect 1365 4803 1366 4807
rect 2386 4803 2390 4807
rect 2394 4803 2397 4807
rect 2397 4803 2398 4807
rect 3402 4803 3406 4807
rect 3410 4803 3413 4807
rect 3413 4803 3414 4807
rect 4426 4803 4430 4807
rect 4434 4803 4437 4807
rect 4437 4803 4438 4807
rect 2190 4798 2194 4802
rect 2214 4798 2218 4802
rect 4150 4798 4154 4802
rect 4398 4798 4402 4802
rect 4558 4798 4562 4802
rect 4582 4798 4586 4802
rect 606 4788 610 4792
rect 742 4788 746 4792
rect 2158 4788 2162 4792
rect 2422 4788 2426 4792
rect 3686 4788 3690 4792
rect 4038 4788 4042 4792
rect 4078 4788 4082 4792
rect 4134 4788 4138 4792
rect 4502 4788 4506 4792
rect 4974 4788 4978 4792
rect 5302 4788 5306 4792
rect 430 4778 434 4782
rect 494 4778 498 4782
rect 638 4778 642 4782
rect 2358 4778 2362 4782
rect 438 4768 442 4772
rect 462 4768 466 4772
rect 662 4768 666 4772
rect 1342 4768 1346 4772
rect 1606 4768 1610 4772
rect 1854 4768 1858 4772
rect 3182 4768 3186 4772
rect 3422 4768 3426 4772
rect 4686 4768 4690 4772
rect 5078 4768 5082 4772
rect 86 4758 90 4762
rect 286 4758 290 4762
rect 734 4758 738 4762
rect 998 4758 1002 4762
rect 1038 4758 1042 4762
rect 1134 4758 1138 4762
rect 2094 4758 2098 4762
rect 2654 4758 2658 4762
rect 46 4748 50 4752
rect 414 4748 418 4752
rect 422 4748 426 4752
rect 854 4748 858 4752
rect 1254 4748 1258 4752
rect 1310 4748 1314 4752
rect 1446 4748 1450 4752
rect 1566 4748 1570 4752
rect 1710 4748 1714 4752
rect 2350 4748 2354 4752
rect 2486 4748 2490 4752
rect 2606 4748 2610 4752
rect 2878 4748 2882 4752
rect 3054 4748 3058 4752
rect 142 4738 146 4742
rect 214 4738 218 4742
rect 1134 4738 1138 4742
rect 3702 4748 3706 4752
rect 4150 4748 4154 4752
rect 4574 4748 4578 4752
rect 4782 4748 4786 4752
rect 5038 4748 5042 4752
rect 2870 4738 2874 4742
rect 3358 4738 3362 4742
rect 4030 4738 4034 4742
rect 4094 4738 4098 4742
rect 4766 4738 4770 4742
rect 630 4728 634 4732
rect 742 4728 746 4732
rect 854 4728 858 4732
rect 918 4728 922 4732
rect 1110 4728 1114 4732
rect 1174 4728 1178 4732
rect 1606 4728 1610 4732
rect 1614 4728 1618 4732
rect 1798 4728 1802 4732
rect 2182 4728 2186 4732
rect 2422 4728 2426 4732
rect 2598 4728 2602 4732
rect 2854 4728 2858 4732
rect 2886 4728 2890 4732
rect 3150 4728 3154 4732
rect 3742 4728 3746 4732
rect 4134 4728 4138 4732
rect 4446 4728 4450 4732
rect 4678 4728 4682 4732
rect 118 4718 122 4722
rect 1014 4718 1018 4722
rect 2006 4718 2010 4722
rect 2662 4718 2666 4722
rect 2846 4718 2850 4722
rect 3606 4718 3610 4722
rect 4206 4718 4210 4722
rect 5054 4718 5058 4722
rect 5174 4718 5178 4722
rect 38 4708 42 4712
rect 934 4708 938 4712
rect 2478 4708 2482 4712
rect 3190 4708 3194 4712
rect 3526 4708 3530 4712
rect 3670 4708 3674 4712
rect 3838 4708 3842 4712
rect 4926 4708 4930 4712
rect 5174 4708 5178 4712
rect 850 4703 854 4707
rect 858 4703 861 4707
rect 861 4703 862 4707
rect 1874 4703 1878 4707
rect 1882 4703 1885 4707
rect 1885 4703 1886 4707
rect 2890 4703 2894 4707
rect 2898 4703 2901 4707
rect 2901 4703 2902 4707
rect 3922 4703 3926 4707
rect 3930 4703 3933 4707
rect 3933 4703 3934 4707
rect 4938 4703 4942 4707
rect 4946 4703 4949 4707
rect 4949 4703 4950 4707
rect 726 4698 730 4702
rect 790 4698 794 4702
rect 918 4698 922 4702
rect 950 4698 954 4702
rect 1654 4698 1658 4702
rect 2374 4698 2378 4702
rect 3438 4698 3442 4702
rect 4030 4698 4034 4702
rect 4414 4698 4418 4702
rect 4638 4698 4642 4702
rect 5102 4698 5106 4702
rect 126 4688 130 4692
rect 3342 4688 3346 4692
rect 4070 4688 4074 4692
rect 4254 4688 4258 4692
rect 4854 4688 4858 4692
rect 4926 4688 4930 4692
rect 5158 4688 5162 4692
rect 326 4678 330 4682
rect 1342 4678 1346 4682
rect 2902 4678 2906 4682
rect 4230 4678 4234 4682
rect 4654 4678 4658 4682
rect 126 4668 130 4672
rect 342 4668 346 4672
rect 670 4668 674 4672
rect 1262 4668 1266 4672
rect 1534 4668 1538 4672
rect 2422 4668 2426 4672
rect 2750 4668 2754 4672
rect 3374 4668 3378 4672
rect 278 4658 282 4662
rect 742 4658 746 4662
rect 838 4658 842 4662
rect 1102 4658 1106 4662
rect 1318 4658 1322 4662
rect 2126 4658 2130 4662
rect 2934 4658 2938 4662
rect 3270 4658 3274 4662
rect 3278 4658 3282 4662
rect 3654 4658 3658 4662
rect 4550 4658 4554 4662
rect 4670 4658 4674 4662
rect 5142 4658 5146 4662
rect 222 4648 226 4652
rect 326 4648 330 4652
rect 342 4648 346 4652
rect 590 4648 594 4652
rect 774 4648 778 4652
rect 2054 4648 2058 4652
rect 3070 4648 3074 4652
rect 3550 4648 3554 4652
rect 214 4638 218 4642
rect 414 4638 418 4642
rect 486 4638 490 4642
rect 2846 4638 2850 4642
rect 3230 4638 3234 4642
rect 3630 4638 3634 4642
rect 5022 4638 5026 4642
rect 5150 4638 5154 4642
rect 2742 4628 2746 4632
rect 3230 4628 3234 4632
rect 3726 4628 3730 4632
rect 4478 4628 4482 4632
rect 214 4618 218 4622
rect 358 4618 362 4622
rect 582 4618 586 4622
rect 598 4618 602 4622
rect 822 4618 826 4622
rect 1606 4618 1610 4622
rect 2798 4618 2802 4622
rect 3782 4618 3786 4622
rect 4414 4618 4418 4622
rect 590 4608 594 4612
rect 694 4608 698 4612
rect 1894 4608 1898 4612
rect 2694 4608 2698 4612
rect 330 4603 334 4607
rect 338 4603 341 4607
rect 341 4603 342 4607
rect 1354 4603 1358 4607
rect 1362 4603 1365 4607
rect 1365 4603 1366 4607
rect 2386 4603 2390 4607
rect 2394 4603 2397 4607
rect 2397 4603 2398 4607
rect 3402 4603 3406 4607
rect 3410 4603 3413 4607
rect 3413 4603 3414 4607
rect 4426 4603 4430 4607
rect 4434 4603 4437 4607
rect 4437 4603 4438 4607
rect 94 4598 98 4602
rect 670 4598 674 4602
rect 4574 4598 4578 4602
rect 4646 4598 4650 4602
rect 726 4588 730 4592
rect 974 4588 978 4592
rect 1246 4588 1250 4592
rect 2734 4588 2738 4592
rect 3478 4588 3482 4592
rect 4054 4588 4058 4592
rect 4630 4588 4634 4592
rect 4654 4588 4658 4592
rect 4918 4588 4922 4592
rect 5230 4588 5234 4592
rect 134 4578 138 4582
rect 1158 4578 1162 4582
rect 2366 4578 2370 4582
rect 3886 4578 3890 4582
rect 4606 4578 4610 4582
rect 5046 4578 5050 4582
rect 414 4568 418 4572
rect 574 4568 578 4572
rect 694 4568 698 4572
rect 1470 4568 1474 4572
rect 2334 4568 2338 4572
rect 2358 4568 2362 4572
rect 3118 4568 3122 4572
rect 3518 4568 3522 4572
rect 4118 4568 4122 4572
rect 4206 4568 4210 4572
rect 4398 4568 4402 4572
rect 454 4558 458 4562
rect 470 4558 474 4562
rect 582 4558 586 4562
rect 1150 4558 1154 4562
rect 1462 4558 1466 4562
rect 1694 4558 1698 4562
rect 2102 4558 2106 4562
rect 2790 4558 2794 4562
rect 3214 4558 3218 4562
rect 3870 4558 3874 4562
rect 3886 4558 3890 4562
rect 4078 4558 4082 4562
rect 4142 4558 4146 4562
rect 4166 4558 4170 4562
rect 4214 4558 4218 4562
rect 4278 4558 4282 4562
rect 4414 4558 4418 4562
rect 4678 4558 4682 4562
rect 4710 4558 4714 4562
rect 4998 4558 5002 4562
rect 5214 4558 5218 4562
rect 494 4548 498 4552
rect 638 4548 642 4552
rect 1358 4548 1362 4552
rect 1454 4548 1458 4552
rect 1646 4548 1650 4552
rect 1958 4548 1962 4552
rect 2190 4548 2194 4552
rect 2414 4548 2418 4552
rect 2814 4548 2818 4552
rect 2958 4548 2962 4552
rect 3286 4548 3290 4552
rect 46 4538 50 4542
rect 174 4538 178 4542
rect 366 4538 370 4542
rect 446 4538 450 4542
rect 598 4538 602 4542
rect 1006 4538 1010 4542
rect 1030 4538 1034 4542
rect 1462 4538 1466 4542
rect 2734 4538 2738 4542
rect 2822 4538 2826 4542
rect 3358 4548 3362 4552
rect 3526 4548 3530 4552
rect 3734 4548 3738 4552
rect 3838 4548 3842 4552
rect 3942 4548 3946 4552
rect 3966 4548 3970 4552
rect 4406 4548 4410 4552
rect 4502 4548 4506 4552
rect 5150 4548 5154 4552
rect 5182 4548 5186 4552
rect 3342 4538 3346 4542
rect 3430 4538 3434 4542
rect 3462 4538 3466 4542
rect 3518 4538 3522 4542
rect 3958 4538 3962 4542
rect 4110 4538 4114 4542
rect 4238 4538 4242 4542
rect 4870 4538 4874 4542
rect 4998 4538 5002 4542
rect 662 4528 666 4532
rect 1038 4528 1042 4532
rect 1126 4528 1130 4532
rect 1662 4528 1666 4532
rect 1950 4528 1954 4532
rect 2734 4528 2738 4532
rect 2862 4528 2866 4532
rect 3470 4528 3474 4532
rect 3998 4528 4002 4532
rect 4142 4528 4146 4532
rect 4206 4528 4210 4532
rect 4662 4528 4666 4532
rect 5166 4528 5170 4532
rect 470 4518 474 4522
rect 542 4518 546 4522
rect 1046 4518 1050 4522
rect 2350 4518 2354 4522
rect 2638 4518 2642 4522
rect 3662 4518 3666 4522
rect 806 4508 810 4512
rect 998 4508 1002 4512
rect 1542 4508 1546 4512
rect 2662 4508 2666 4512
rect 3942 4508 3946 4512
rect 4734 4508 4738 4512
rect 4982 4508 4986 4512
rect 850 4503 854 4507
rect 858 4503 861 4507
rect 861 4503 862 4507
rect 1874 4503 1878 4507
rect 1882 4503 1885 4507
rect 1885 4503 1886 4507
rect 2890 4503 2894 4507
rect 2898 4503 2901 4507
rect 2901 4503 2902 4507
rect 1174 4498 1178 4502
rect 2758 4498 2762 4502
rect 3094 4498 3098 4502
rect 3686 4498 3690 4502
rect 3922 4503 3926 4507
rect 3930 4503 3933 4507
rect 3933 4503 3934 4507
rect 4938 4503 4942 4507
rect 4946 4503 4949 4507
rect 4949 4503 4950 4507
rect 4094 4498 4098 4502
rect 4990 4498 4994 4502
rect 678 4488 682 4492
rect 2750 4488 2754 4492
rect 2942 4488 2946 4492
rect 3934 4488 3938 4492
rect 142 4478 146 4482
rect 390 4478 394 4482
rect 974 4478 978 4482
rect 1070 4478 1074 4482
rect 1342 4478 1346 4482
rect 1662 4478 1666 4482
rect 2406 4478 2410 4482
rect 3590 4478 3594 4482
rect 3718 4478 3722 4482
rect 3942 4478 3946 4482
rect 4390 4478 4394 4482
rect 4966 4478 4970 4482
rect 502 4468 506 4472
rect 558 4468 562 4472
rect 710 4468 714 4472
rect 886 4468 890 4472
rect 942 4468 946 4472
rect 1846 4468 1850 4472
rect 2598 4468 2602 4472
rect 3118 4468 3122 4472
rect 3214 4468 3218 4472
rect 3734 4468 3738 4472
rect 4094 4468 4098 4472
rect 4910 4468 4914 4472
rect 5150 4468 5154 4472
rect 110 4458 114 4462
rect 1158 4458 1162 4462
rect 1310 4458 1314 4462
rect 1998 4458 2002 4462
rect 2078 4458 2082 4462
rect 2134 4458 2138 4462
rect 2342 4458 2346 4462
rect 2566 4458 2570 4462
rect 2686 4458 2690 4462
rect 3062 4458 3066 4462
rect 3086 4458 3090 4462
rect 3126 4458 3130 4462
rect 3838 4458 3842 4462
rect 4030 4458 4034 4462
rect 4038 4458 4042 4462
rect 4246 4458 4250 4462
rect 4630 4458 4634 4462
rect 4854 4458 4858 4462
rect 5182 4458 5186 4462
rect 574 4448 578 4452
rect 718 4448 722 4452
rect 1070 4448 1074 4452
rect 1198 4448 1202 4452
rect 1342 4448 1346 4452
rect 1462 4448 1466 4452
rect 1982 4448 1986 4452
rect 2014 4448 2018 4452
rect 2094 4448 2098 4452
rect 2662 4448 2666 4452
rect 3062 4448 3066 4452
rect 3222 4448 3226 4452
rect 3726 4448 3730 4452
rect 3974 4448 3978 4452
rect 4150 4448 4154 4452
rect 4654 4448 4658 4452
rect 86 4438 90 4442
rect 142 4438 146 4442
rect 774 4438 778 4442
rect 2086 4438 2090 4442
rect 2686 4438 2690 4442
rect 4006 4438 4010 4442
rect 4182 4438 4186 4442
rect 4606 4438 4610 4442
rect 4998 4438 5002 4442
rect 398 4428 402 4432
rect 582 4428 586 4432
rect 822 4428 826 4432
rect 1030 4428 1034 4432
rect 2438 4428 2442 4432
rect 2470 4428 2474 4432
rect 2686 4428 2690 4432
rect 790 4418 794 4422
rect 878 4418 882 4422
rect 1342 4418 1346 4422
rect 2326 4418 2330 4422
rect 3638 4418 3642 4422
rect 4166 4418 4170 4422
rect 4886 4418 4890 4422
rect 5142 4418 5146 4422
rect 5222 4418 5226 4422
rect 550 4408 554 4412
rect 726 4408 730 4412
rect 926 4408 930 4412
rect 1702 4408 1706 4412
rect 2070 4408 2074 4412
rect 3262 4408 3266 4412
rect 4502 4408 4506 4412
rect 330 4403 334 4407
rect 338 4403 341 4407
rect 341 4403 342 4407
rect 1354 4403 1358 4407
rect 1362 4403 1365 4407
rect 1365 4403 1366 4407
rect 2386 4403 2390 4407
rect 2394 4403 2397 4407
rect 2397 4403 2398 4407
rect 3402 4403 3406 4407
rect 3410 4403 3413 4407
rect 3413 4403 3414 4407
rect 4426 4403 4430 4407
rect 4434 4403 4437 4407
rect 4437 4403 4438 4407
rect 798 4398 802 4402
rect 1846 4398 1850 4402
rect 2574 4398 2578 4402
rect 3070 4398 3074 4402
rect 3710 4398 3714 4402
rect 3830 4398 3834 4402
rect 4350 4398 4354 4402
rect 4590 4398 4594 4402
rect 278 4388 282 4392
rect 46 4378 50 4382
rect 558 4378 562 4382
rect 726 4378 730 4382
rect 1214 4378 1218 4382
rect 2150 4378 2154 4382
rect 2446 4378 2450 4382
rect 398 4368 402 4372
rect 638 4368 642 4372
rect 798 4368 802 4372
rect 1078 4368 1082 4372
rect 1918 4368 1922 4372
rect 1926 4368 1930 4372
rect 1950 4368 1954 4372
rect 2422 4368 2426 4372
rect 3022 4368 3026 4372
rect 3662 4368 3666 4372
rect 4134 4368 4138 4372
rect 4294 4368 4298 4372
rect 5038 4368 5042 4372
rect 1190 4358 1194 4362
rect 1478 4358 1482 4362
rect 1830 4358 1834 4362
rect 2774 4358 2778 4362
rect 4086 4358 4090 4362
rect 4214 4358 4218 4362
rect 4454 4358 4458 4362
rect 4646 4358 4650 4362
rect 5118 4358 5122 4362
rect 5150 4358 5154 4362
rect 102 4348 106 4352
rect 382 4348 386 4352
rect 454 4348 458 4352
rect 702 4348 706 4352
rect 742 4348 746 4352
rect 806 4348 810 4352
rect 886 4348 890 4352
rect 1022 4348 1026 4352
rect 1262 4348 1266 4352
rect 1718 4348 1722 4352
rect 2414 4348 2418 4352
rect 2726 4348 2730 4352
rect 2838 4348 2842 4352
rect 86 4338 90 4342
rect 462 4338 466 4342
rect 566 4338 570 4342
rect 694 4338 698 4342
rect 2446 4338 2450 4342
rect 2518 4338 2522 4342
rect 2726 4338 2730 4342
rect 2798 4338 2802 4342
rect 3334 4348 3338 4352
rect 3406 4348 3410 4352
rect 3782 4348 3786 4352
rect 3854 4348 3858 4352
rect 3878 4348 3882 4352
rect 3934 4348 3938 4352
rect 4190 4348 4194 4352
rect 4206 4348 4210 4352
rect 4494 4348 4498 4352
rect 5102 4348 5106 4352
rect 5118 4348 5122 4352
rect 4062 4338 4066 4342
rect 4126 4338 4130 4342
rect 4182 4338 4186 4342
rect 4486 4338 4490 4342
rect 4622 4338 4626 4342
rect 4718 4338 4722 4342
rect 5102 4338 5106 4342
rect 5198 4338 5202 4342
rect 5246 4338 5250 4342
rect 486 4328 490 4332
rect 678 4328 682 4332
rect 702 4328 706 4332
rect 1262 4328 1266 4332
rect 1534 4328 1538 4332
rect 2574 4328 2578 4332
rect 2878 4328 2882 4332
rect 3518 4328 3522 4332
rect 3694 4328 3698 4332
rect 3838 4328 3842 4332
rect 254 4318 258 4322
rect 2014 4318 2018 4322
rect 3382 4318 3386 4322
rect 4910 4318 4914 4322
rect 5246 4318 5250 4322
rect 2262 4308 2266 4312
rect 3270 4308 3274 4312
rect 3830 4308 3834 4312
rect 4926 4308 4930 4312
rect 5182 4308 5186 4312
rect 850 4303 854 4307
rect 858 4303 861 4307
rect 861 4303 862 4307
rect 1874 4303 1878 4307
rect 1882 4303 1885 4307
rect 1885 4303 1886 4307
rect 2890 4303 2894 4307
rect 2898 4303 2901 4307
rect 2901 4303 2902 4307
rect 3922 4303 3926 4307
rect 3930 4303 3933 4307
rect 3933 4303 3934 4307
rect 4938 4303 4942 4307
rect 4946 4303 4949 4307
rect 4949 4303 4950 4307
rect 22 4298 26 4302
rect 414 4298 418 4302
rect 2270 4298 2274 4302
rect 3390 4298 3394 4302
rect 4078 4298 4082 4302
rect 4542 4298 4546 4302
rect 5158 4298 5162 4302
rect 5174 4298 5178 4302
rect 366 4288 370 4292
rect 774 4288 778 4292
rect 2462 4288 2466 4292
rect 2574 4288 2578 4292
rect 2590 4288 2594 4292
rect 2966 4288 2970 4292
rect 4110 4288 4114 4292
rect 4398 4288 4402 4292
rect 4414 4288 4418 4292
rect 4646 4288 4650 4292
rect 198 4278 202 4282
rect 214 4278 218 4282
rect 470 4278 474 4282
rect 1022 4278 1026 4282
rect 1190 4278 1194 4282
rect 2054 4278 2058 4282
rect 2470 4278 2474 4282
rect 2510 4278 2514 4282
rect 2638 4278 2642 4282
rect 2822 4278 2826 4282
rect 2894 4278 2898 4282
rect 3006 4278 3010 4282
rect 3174 4278 3178 4282
rect 4406 4278 4410 4282
rect 4478 4278 4482 4282
rect 4670 4278 4674 4282
rect 4750 4278 4754 4282
rect 5006 4278 5010 4282
rect 5030 4278 5034 4282
rect 5166 4278 5170 4282
rect 5182 4278 5186 4282
rect 254 4268 258 4272
rect 582 4268 586 4272
rect 742 4268 746 4272
rect 1302 4268 1306 4272
rect 1654 4268 1658 4272
rect 1686 4268 1690 4272
rect 1926 4268 1930 4272
rect 2022 4268 2026 4272
rect 2206 4268 2210 4272
rect 2358 4268 2362 4272
rect 2478 4268 2482 4272
rect 2726 4268 2730 4272
rect 2862 4268 2866 4272
rect 3166 4268 3170 4272
rect 3206 4268 3210 4272
rect 3742 4268 3746 4272
rect 4134 4268 4138 4272
rect 4158 4268 4162 4272
rect 4214 4268 4218 4272
rect 4254 4268 4258 4272
rect 4878 4268 4882 4272
rect 5054 4268 5058 4272
rect 94 4258 98 4262
rect 222 4258 226 4262
rect 590 4258 594 4262
rect 614 4258 618 4262
rect 622 4258 626 4262
rect 766 4258 770 4262
rect 790 4258 794 4262
rect 814 4258 818 4262
rect 878 4258 882 4262
rect 974 4258 978 4262
rect 1654 4258 1658 4262
rect 1822 4258 1826 4262
rect 2062 4258 2066 4262
rect 2198 4258 2202 4262
rect 2534 4258 2538 4262
rect 2566 4258 2570 4262
rect 2814 4258 2818 4262
rect 3270 4258 3274 4262
rect 3558 4258 3562 4262
rect 3598 4258 3602 4262
rect 3686 4258 3690 4262
rect 4118 4258 4122 4262
rect 4158 4258 4162 4262
rect 4566 4258 4570 4262
rect 4822 4258 4826 4262
rect 4838 4258 4842 4262
rect 5022 4258 5026 4262
rect 406 4248 410 4252
rect 638 4248 642 4252
rect 654 4248 658 4252
rect 1038 4248 1042 4252
rect 1670 4248 1674 4252
rect 1750 4248 1754 4252
rect 2126 4248 2130 4252
rect 2206 4248 2210 4252
rect 2830 4248 2834 4252
rect 2926 4248 2930 4252
rect 2958 4248 2962 4252
rect 3518 4248 3522 4252
rect 4070 4248 4074 4252
rect 4214 4248 4218 4252
rect 4550 4248 4554 4252
rect 4806 4248 4810 4252
rect 398 4238 402 4242
rect 830 4238 834 4242
rect 1966 4238 1970 4242
rect 2198 4238 2202 4242
rect 2486 4238 2490 4242
rect 2494 4238 2498 4242
rect 2854 4238 2858 4242
rect 2918 4238 2922 4242
rect 2950 4238 2954 4242
rect 3454 4238 3458 4242
rect 4734 4238 4738 4242
rect 4854 4238 4858 4242
rect 5142 4238 5146 4242
rect 2070 4228 2074 4232
rect 2766 4228 2770 4232
rect 2862 4228 2866 4232
rect 3014 4228 3018 4232
rect 3382 4228 3386 4232
rect 4350 4228 4354 4232
rect 470 4218 474 4222
rect 718 4218 722 4222
rect 1734 4218 1738 4222
rect 1774 4218 1778 4222
rect 2814 4218 2818 4222
rect 3454 4218 3458 4222
rect 3494 4218 3498 4222
rect 3670 4218 3674 4222
rect 4814 4218 4818 4222
rect 1966 4208 1970 4212
rect 4006 4208 4010 4212
rect 4094 4208 4098 4212
rect 4182 4208 4186 4212
rect 4478 4208 4482 4212
rect 5158 4208 5162 4212
rect 330 4203 334 4207
rect 338 4203 341 4207
rect 341 4203 342 4207
rect 1354 4203 1358 4207
rect 1362 4203 1365 4207
rect 1365 4203 1366 4207
rect 2386 4203 2390 4207
rect 2394 4203 2397 4207
rect 2397 4203 2398 4207
rect 3402 4203 3406 4207
rect 3410 4203 3413 4207
rect 3413 4203 3414 4207
rect 4426 4203 4430 4207
rect 4434 4203 4437 4207
rect 4437 4203 4438 4207
rect 726 4198 730 4202
rect 886 4198 890 4202
rect 1990 4198 1994 4202
rect 2238 4198 2242 4202
rect 2446 4198 2450 4202
rect 3022 4198 3026 4202
rect 3758 4198 3762 4202
rect 4398 4198 4402 4202
rect 4526 4198 4530 4202
rect 4838 4198 4842 4202
rect 142 4188 146 4192
rect 350 4188 354 4192
rect 630 4188 634 4192
rect 1390 4188 1394 4192
rect 1918 4188 1922 4192
rect 2214 4188 2218 4192
rect 2454 4188 2458 4192
rect 2774 4188 2778 4192
rect 2838 4188 2842 4192
rect 3702 4188 3706 4192
rect 3790 4188 3794 4192
rect 3822 4188 3826 4192
rect 4358 4188 4362 4192
rect 534 4178 538 4182
rect 2782 4178 2786 4182
rect 3078 4178 3082 4182
rect 3630 4178 3634 4182
rect 3662 4178 3666 4182
rect 3830 4178 3834 4182
rect 14 4168 18 4172
rect 686 4168 690 4172
rect 710 4168 714 4172
rect 1806 4168 1810 4172
rect 2206 4168 2210 4172
rect 3238 4168 3242 4172
rect 3638 4168 3642 4172
rect 4318 4168 4322 4172
rect 4670 4168 4674 4172
rect 5278 4168 5282 4172
rect 414 4158 418 4162
rect 510 4158 514 4162
rect 534 4158 538 4162
rect 694 4158 698 4162
rect 1174 4158 1178 4162
rect 1478 4158 1482 4162
rect 1830 4158 1834 4162
rect 2582 4158 2586 4162
rect 3038 4158 3042 4162
rect 3318 4158 3322 4162
rect 3494 4158 3498 4162
rect 3902 4158 3906 4162
rect 4342 4158 4346 4162
rect 4694 4158 4698 4162
rect 4886 4158 4890 4162
rect 1286 4148 1290 4152
rect 1718 4148 1722 4152
rect 2166 4148 2170 4152
rect 2190 4148 2194 4152
rect 2350 4148 2354 4152
rect 2438 4148 2442 4152
rect 2614 4148 2618 4152
rect 3286 4148 3290 4152
rect 4094 4148 4098 4152
rect 4190 4148 4194 4152
rect 4470 4148 4474 4152
rect 4734 4148 4738 4152
rect 502 4138 506 4142
rect 1206 4138 1210 4142
rect 1454 4138 1458 4142
rect 1854 4138 1858 4142
rect 1878 4138 1882 4142
rect 1910 4138 1914 4142
rect 2110 4138 2114 4142
rect 2134 4138 2138 4142
rect 2246 4138 2250 4142
rect 2782 4138 2786 4142
rect 2822 4138 2826 4142
rect 3038 4138 3042 4142
rect 3110 4138 3114 4142
rect 3742 4138 3746 4142
rect 3854 4138 3858 4142
rect 4166 4138 4170 4142
rect 4326 4138 4330 4142
rect 4486 4138 4490 4142
rect 4638 4138 4642 4142
rect 4926 4138 4930 4142
rect 478 4128 482 4132
rect 542 4128 546 4132
rect 638 4128 642 4132
rect 1294 4128 1298 4132
rect 2118 4128 2122 4132
rect 2318 4128 2322 4132
rect 2510 4128 2514 4132
rect 2646 4128 2650 4132
rect 2718 4128 2722 4132
rect 3006 4128 3010 4132
rect 3254 4128 3258 4132
rect 3286 4128 3290 4132
rect 4046 4128 4050 4132
rect 4398 4128 4402 4132
rect 4606 4128 4610 4132
rect 5094 4128 5098 4132
rect 366 4118 370 4122
rect 534 4118 538 4122
rect 550 4118 554 4122
rect 566 4118 570 4122
rect 1278 4118 1282 4122
rect 1742 4118 1746 4122
rect 1814 4118 1818 4122
rect 1950 4118 1954 4122
rect 2742 4118 2746 4122
rect 2934 4118 2938 4122
rect 3454 4118 3458 4122
rect 3902 4118 3906 4122
rect 3910 4118 3914 4122
rect 4254 4118 4258 4122
rect 4278 4118 4282 4122
rect 4662 4118 4666 4122
rect 158 4108 162 4112
rect 622 4108 626 4112
rect 638 4108 642 4112
rect 1686 4108 1690 4112
rect 2582 4108 2586 4112
rect 2670 4108 2674 4112
rect 3198 4108 3202 4112
rect 3518 4108 3522 4112
rect 4102 4108 4106 4112
rect 4710 4108 4714 4112
rect 5182 4108 5186 4112
rect 850 4103 854 4107
rect 858 4103 861 4107
rect 861 4103 862 4107
rect 1874 4103 1878 4107
rect 1882 4103 1885 4107
rect 1885 4103 1886 4107
rect 2890 4103 2894 4107
rect 2898 4103 2901 4107
rect 2901 4103 2902 4107
rect 3922 4103 3926 4107
rect 3930 4103 3933 4107
rect 3933 4103 3934 4107
rect 4938 4103 4942 4107
rect 4946 4103 4949 4107
rect 4949 4103 4950 4107
rect 254 4098 258 4102
rect 542 4098 546 4102
rect 1566 4098 1570 4102
rect 1646 4098 1650 4102
rect 2574 4098 2578 4102
rect 2614 4098 2618 4102
rect 3486 4098 3490 4102
rect 4262 4098 4266 4102
rect 4510 4098 4514 4102
rect 5126 4098 5130 4102
rect 5142 4098 5146 4102
rect 198 4088 202 4092
rect 566 4088 570 4092
rect 1926 4088 1930 4092
rect 1934 4088 1938 4092
rect 2846 4088 2850 4092
rect 3126 4088 3130 4092
rect 3646 4088 3650 4092
rect 4366 4088 4370 4092
rect 358 4078 362 4082
rect 558 4078 562 4082
rect 630 4078 634 4082
rect 838 4078 842 4082
rect 1718 4078 1722 4082
rect 1758 4078 1762 4082
rect 1782 4078 1786 4082
rect 1918 4078 1922 4082
rect 1942 4078 1946 4082
rect 2374 4078 2378 4082
rect 2502 4078 2506 4082
rect 3182 4078 3186 4082
rect 3342 4078 3346 4082
rect 3718 4078 3722 4082
rect 3894 4078 3898 4082
rect 3910 4078 3914 4082
rect 4054 4078 4058 4082
rect 5182 4078 5186 4082
rect 582 4068 586 4072
rect 726 4068 730 4072
rect 2126 4068 2130 4072
rect 2134 4068 2138 4072
rect 2454 4068 2458 4072
rect 3014 4068 3018 4072
rect 3054 4068 3058 4072
rect 4230 4068 4234 4072
rect 4238 4068 4242 4072
rect 4286 4068 4290 4072
rect 4414 4068 4418 4072
rect 4646 4068 4650 4072
rect 5046 4068 5050 4072
rect 414 4058 418 4062
rect 566 4058 570 4062
rect 1502 4058 1506 4062
rect 1654 4058 1658 4062
rect 1710 4058 1714 4062
rect 1846 4058 1850 4062
rect 1966 4058 1970 4062
rect 2014 4058 2018 4062
rect 2078 4058 2082 4062
rect 2238 4058 2242 4062
rect 2606 4058 2610 4062
rect 3094 4058 3098 4062
rect 3438 4058 3442 4062
rect 3630 4058 3634 4062
rect 4078 4058 4082 4062
rect 4086 4058 4090 4062
rect 4294 4058 4298 4062
rect 158 4048 162 4052
rect 278 4048 282 4052
rect 494 4048 498 4052
rect 1390 4048 1394 4052
rect 1446 4048 1450 4052
rect 1846 4048 1850 4052
rect 2046 4048 2050 4052
rect 2054 4048 2058 4052
rect 3158 4048 3162 4052
rect 3198 4048 3202 4052
rect 3310 4048 3314 4052
rect 3710 4048 3714 4052
rect 3774 4048 3778 4052
rect 4070 4048 4074 4052
rect 4238 4048 4242 4052
rect 4286 4048 4290 4052
rect 5166 4048 5170 4052
rect 110 4038 114 4042
rect 638 4038 642 4042
rect 1678 4038 1682 4042
rect 2078 4038 2082 4042
rect 2470 4038 2474 4042
rect 2734 4038 2738 4042
rect 3726 4038 3730 4042
rect 4246 4038 4250 4042
rect 4462 4038 4466 4042
rect 510 4028 514 4032
rect 566 4028 570 4032
rect 1294 4028 1298 4032
rect 2142 4028 2146 4032
rect 2854 4028 2858 4032
rect 2870 4028 2874 4032
rect 3854 4028 3858 4032
rect 3974 4028 3978 4032
rect 1662 4018 1666 4022
rect 1742 4018 1746 4022
rect 2550 4018 2554 4022
rect 2822 4018 2826 4022
rect 3510 4018 3514 4022
rect 3702 4018 3706 4022
rect 4158 4018 4162 4022
rect 4494 4018 4498 4022
rect 494 4008 498 4012
rect 1374 4008 1378 4012
rect 2078 4008 2082 4012
rect 2326 4008 2330 4012
rect 2510 4008 2514 4012
rect 2878 4008 2882 4012
rect 4358 4008 4362 4012
rect 5198 4008 5202 4012
rect 330 4003 334 4007
rect 338 4003 341 4007
rect 341 4003 342 4007
rect 1354 4003 1358 4007
rect 1362 4003 1365 4007
rect 1365 4003 1366 4007
rect 2386 4003 2390 4007
rect 2394 4003 2397 4007
rect 2397 4003 2398 4007
rect 3402 4003 3406 4007
rect 3410 4003 3413 4007
rect 3413 4003 3414 4007
rect 4426 4003 4430 4007
rect 4434 4003 4437 4007
rect 4437 4003 4438 4007
rect 350 3998 354 4002
rect 1838 3998 1842 4002
rect 1854 3998 1858 4002
rect 1974 3998 1978 4002
rect 2206 3998 2210 4002
rect 3470 3998 3474 4002
rect 4358 3998 4362 4002
rect 142 3988 146 3992
rect 414 3988 418 3992
rect 1710 3988 1714 3992
rect 3526 3988 3530 3992
rect 3614 3988 3618 3992
rect 5110 3988 5114 3992
rect 5134 3988 5138 3992
rect 78 3978 82 3982
rect 582 3978 586 3982
rect 590 3978 594 3982
rect 1694 3978 1698 3982
rect 2134 3978 2138 3982
rect 4302 3978 4306 3982
rect 4726 3978 4730 3982
rect 38 3968 42 3972
rect 350 3968 354 3972
rect 574 3968 578 3972
rect 2494 3968 2498 3972
rect 3574 3968 3578 3972
rect 3678 3968 3682 3972
rect 4038 3968 4042 3972
rect 4758 3968 4762 3972
rect 142 3958 146 3962
rect 310 3958 314 3962
rect 446 3958 450 3962
rect 1110 3958 1114 3962
rect 2326 3958 2330 3962
rect 2950 3958 2954 3962
rect 3390 3958 3394 3962
rect 3638 3958 3642 3962
rect 3862 3958 3866 3962
rect 4126 3958 4130 3962
rect 4342 3958 4346 3962
rect 4494 3958 4498 3962
rect 4918 3958 4922 3962
rect 5038 3958 5042 3962
rect 5158 3958 5162 3962
rect 390 3948 394 3952
rect 502 3948 506 3952
rect 558 3948 562 3952
rect 734 3948 738 3952
rect 1286 3948 1290 3952
rect 1670 3948 1674 3952
rect 1894 3948 1898 3952
rect 2006 3948 2010 3952
rect 2038 3948 2042 3952
rect 2086 3948 2090 3952
rect 2134 3948 2138 3952
rect 2174 3948 2178 3952
rect 2430 3948 2434 3952
rect 2438 3948 2442 3952
rect 2862 3948 2866 3952
rect 2878 3948 2882 3952
rect 3182 3948 3186 3952
rect 3374 3948 3378 3952
rect 3494 3948 3498 3952
rect 3502 3948 3506 3952
rect 3646 3948 3650 3952
rect 3718 3948 3722 3952
rect 3790 3948 3794 3952
rect 4022 3948 4026 3952
rect 4086 3948 4090 3952
rect 4270 3948 4274 3952
rect 4510 3948 4514 3952
rect 4606 3948 4610 3952
rect 4886 3948 4890 3952
rect 4982 3948 4986 3952
rect 4998 3948 5002 3952
rect 5046 3948 5050 3952
rect 382 3938 386 3942
rect 1374 3938 1378 3942
rect 1790 3938 1794 3942
rect 1934 3938 1938 3942
rect 1942 3938 1946 3942
rect 2014 3938 2018 3942
rect 2030 3938 2034 3942
rect 2206 3938 2210 3942
rect 2326 3938 2330 3942
rect 2854 3938 2858 3942
rect 3382 3938 3386 3942
rect 3398 3938 3402 3942
rect 3566 3938 3570 3942
rect 3614 3938 3618 3942
rect 3654 3938 3658 3942
rect 5118 3948 5122 3952
rect 4806 3938 4810 3942
rect 4894 3938 4898 3942
rect 198 3928 202 3932
rect 1270 3928 1274 3932
rect 1414 3928 1418 3932
rect 1574 3928 1578 3932
rect 1742 3928 1746 3932
rect 1750 3928 1754 3932
rect 1822 3928 1826 3932
rect 1982 3928 1986 3932
rect 2182 3928 2186 3932
rect 2198 3928 2202 3932
rect 2438 3928 2442 3932
rect 3230 3928 3234 3932
rect 3734 3928 3738 3932
rect 4990 3938 4994 3942
rect 5046 3938 5050 3942
rect 5166 3938 5170 3942
rect 4070 3928 4074 3932
rect 4118 3928 4122 3932
rect 4390 3928 4394 3932
rect 4606 3928 4610 3932
rect 4998 3928 5002 3932
rect 5270 3928 5274 3932
rect 870 3918 874 3922
rect 1662 3918 1666 3922
rect 2230 3918 2234 3922
rect 2326 3918 2330 3922
rect 3654 3918 3658 3922
rect 4102 3918 4106 3922
rect 4958 3918 4962 3922
rect 5022 3918 5026 3922
rect 198 3908 202 3912
rect 542 3908 546 3912
rect 838 3908 842 3912
rect 1222 3908 1226 3912
rect 1390 3908 1394 3912
rect 2718 3908 2722 3912
rect 3582 3908 3586 3912
rect 4126 3908 4130 3912
rect 4134 3908 4138 3912
rect 4502 3908 4506 3912
rect 4534 3908 4538 3912
rect 850 3903 854 3907
rect 858 3903 861 3907
rect 861 3903 862 3907
rect 1874 3903 1878 3907
rect 1882 3903 1885 3907
rect 1885 3903 1886 3907
rect 2890 3903 2894 3907
rect 2898 3903 2901 3907
rect 2901 3903 2902 3907
rect 3922 3903 3926 3907
rect 3930 3903 3933 3907
rect 3933 3903 3934 3907
rect 4938 3903 4942 3907
rect 4946 3903 4949 3907
rect 4949 3903 4950 3907
rect 510 3898 514 3902
rect 870 3898 874 3902
rect 1206 3898 1210 3902
rect 1790 3898 1794 3902
rect 2830 3898 2834 3902
rect 3382 3898 3386 3902
rect 3574 3898 3578 3902
rect 3694 3898 3698 3902
rect 4030 3898 4034 3902
rect 4590 3898 4594 3902
rect 550 3888 554 3892
rect 2134 3888 2138 3892
rect 2334 3888 2338 3892
rect 2614 3888 2618 3892
rect 3230 3888 3234 3892
rect 3622 3888 3626 3892
rect 3646 3888 3650 3892
rect 118 3878 122 3882
rect 966 3878 970 3882
rect 1158 3878 1162 3882
rect 1174 3878 1178 3882
rect 1222 3878 1226 3882
rect 1230 3878 1234 3882
rect 1350 3878 1354 3882
rect 1486 3878 1490 3882
rect 1774 3878 1778 3882
rect 2422 3878 2426 3882
rect 2910 3878 2914 3882
rect 3686 3878 3690 3882
rect 3694 3878 3698 3882
rect 3998 3878 4002 3882
rect 4454 3878 4458 3882
rect 4590 3878 4594 3882
rect 1302 3868 1306 3872
rect 1326 3868 1330 3872
rect 1814 3868 1818 3872
rect 1822 3868 1826 3872
rect 1838 3868 1842 3872
rect 1918 3868 1922 3872
rect 2054 3868 2058 3872
rect 2086 3868 2090 3872
rect 2102 3868 2106 3872
rect 2134 3868 2138 3872
rect 2406 3868 2410 3872
rect 2670 3868 2674 3872
rect 2686 3868 2690 3872
rect 2742 3868 2746 3872
rect 2950 3868 2954 3872
rect 3118 3868 3122 3872
rect 3174 3868 3178 3872
rect 3430 3868 3434 3872
rect 3494 3868 3498 3872
rect 3798 3868 3802 3872
rect 4206 3868 4210 3872
rect 4998 3868 5002 3872
rect 5030 3868 5034 3872
rect 5174 3868 5178 3872
rect 118 3858 122 3862
rect 382 3858 386 3862
rect 934 3858 938 3862
rect 998 3858 1002 3862
rect 1062 3858 1066 3862
rect 1086 3858 1090 3862
rect 1094 3858 1098 3862
rect 1302 3858 1306 3862
rect 1310 3858 1314 3862
rect 1374 3858 1378 3862
rect 1742 3858 1746 3862
rect 1894 3858 1898 3862
rect 2006 3858 2010 3862
rect 2150 3858 2154 3862
rect 2854 3858 2858 3862
rect 3302 3858 3306 3862
rect 3630 3858 3634 3862
rect 3718 3858 3722 3862
rect 4246 3858 4250 3862
rect 4334 3858 4338 3862
rect 4462 3858 4466 3862
rect 5166 3858 5170 3862
rect 5198 3858 5202 3862
rect 5246 3858 5250 3862
rect 222 3848 226 3852
rect 702 3848 706 3852
rect 1798 3848 1802 3852
rect 1838 3848 1842 3852
rect 2038 3848 2042 3852
rect 2062 3848 2066 3852
rect 2342 3848 2346 3852
rect 2358 3848 2362 3852
rect 2934 3848 2938 3852
rect 3070 3848 3074 3852
rect 3102 3848 3106 3852
rect 3374 3848 3378 3852
rect 3590 3848 3594 3852
rect 3806 3848 3810 3852
rect 3886 3848 3890 3852
rect 4374 3848 4378 3852
rect 4894 3848 4898 3852
rect 4982 3848 4986 3852
rect 5038 3848 5042 3852
rect 94 3838 98 3842
rect 102 3838 106 3842
rect 446 3838 450 3842
rect 470 3838 474 3842
rect 1030 3838 1034 3842
rect 2006 3838 2010 3842
rect 2446 3838 2450 3842
rect 2870 3838 2874 3842
rect 3094 3838 3098 3842
rect 3446 3838 3450 3842
rect 4894 3838 4898 3842
rect 5150 3838 5154 3842
rect 126 3828 130 3832
rect 1494 3828 1498 3832
rect 2094 3828 2098 3832
rect 3214 3828 3218 3832
rect 3462 3828 3466 3832
rect 102 3818 106 3822
rect 310 3818 314 3822
rect 478 3818 482 3822
rect 2670 3818 2674 3822
rect 3070 3818 3074 3822
rect 3270 3818 3274 3822
rect 3686 3818 3690 3822
rect 4854 3818 4858 3822
rect 4870 3818 4874 3822
rect 5126 3818 5130 3822
rect 126 3808 130 3812
rect 318 3808 322 3812
rect 1694 3808 1698 3812
rect 2294 3808 2298 3812
rect 3342 3808 3346 3812
rect 3462 3808 3466 3812
rect 4302 3808 4306 3812
rect 330 3803 334 3807
rect 338 3803 341 3807
rect 341 3803 342 3807
rect 1354 3803 1358 3807
rect 1362 3803 1365 3807
rect 1365 3803 1366 3807
rect 2386 3803 2390 3807
rect 2394 3803 2397 3807
rect 2397 3803 2398 3807
rect 3402 3803 3406 3807
rect 3410 3803 3413 3807
rect 3413 3803 3414 3807
rect 4426 3803 4430 3807
rect 4434 3803 4437 3807
rect 4437 3803 4438 3807
rect 1014 3798 1018 3802
rect 1534 3798 1538 3802
rect 2510 3798 2514 3802
rect 3086 3798 3090 3802
rect 3526 3798 3530 3802
rect 4718 3798 4722 3802
rect 5118 3798 5122 3802
rect 1446 3788 1450 3792
rect 1582 3788 1586 3792
rect 2398 3788 2402 3792
rect 2878 3788 2882 3792
rect 3150 3788 3154 3792
rect 4110 3788 4114 3792
rect 4366 3788 4370 3792
rect 1502 3778 1506 3782
rect 1558 3778 1562 3782
rect 2022 3778 2026 3782
rect 2110 3778 2114 3782
rect 2806 3778 2810 3782
rect 3094 3778 3098 3782
rect 3134 3778 3138 3782
rect 3438 3778 3442 3782
rect 4542 3778 4546 3782
rect 46 3768 50 3772
rect 86 3768 90 3772
rect 134 3768 138 3772
rect 646 3768 650 3772
rect 1422 3768 1426 3772
rect 1934 3768 1938 3772
rect 2838 3768 2842 3772
rect 3118 3768 3122 3772
rect 3758 3768 3762 3772
rect 4382 3768 4386 3772
rect 4414 3768 4418 3772
rect 5110 3768 5114 3772
rect 206 3758 210 3762
rect 1150 3758 1154 3762
rect 2222 3758 2226 3762
rect 2302 3758 2306 3762
rect 2438 3758 2442 3762
rect 2526 3758 2530 3762
rect 3038 3758 3042 3762
rect 3142 3758 3146 3762
rect 3190 3758 3194 3762
rect 3262 3758 3266 3762
rect 3462 3758 3466 3762
rect 3470 3758 3474 3762
rect 3998 3758 4002 3762
rect 4006 3758 4010 3762
rect 4054 3758 4058 3762
rect 4334 3758 4338 3762
rect 4542 3758 4546 3762
rect 4630 3758 4634 3762
rect 4990 3758 4994 3762
rect 5134 3758 5138 3762
rect 46 3748 50 3752
rect 78 3748 82 3752
rect 94 3748 98 3752
rect 1302 3748 1306 3752
rect 1510 3748 1514 3752
rect 1598 3748 1602 3752
rect 1726 3748 1730 3752
rect 1934 3748 1938 3752
rect 2406 3748 2410 3752
rect 2790 3748 2794 3752
rect 3214 3748 3218 3752
rect 3366 3748 3370 3752
rect 3382 3748 3386 3752
rect 4374 3748 4378 3752
rect 4630 3748 4634 3752
rect 4846 3748 4850 3752
rect 4926 3748 4930 3752
rect 4982 3748 4986 3752
rect 102 3738 106 3742
rect 510 3738 514 3742
rect 1230 3738 1234 3742
rect 1246 3738 1250 3742
rect 1478 3738 1482 3742
rect 1582 3738 1586 3742
rect 1614 3738 1618 3742
rect 1638 3738 1642 3742
rect 1686 3738 1690 3742
rect 1694 3738 1698 3742
rect 1902 3738 1906 3742
rect 1950 3738 1954 3742
rect 2078 3738 2082 3742
rect 2438 3738 2442 3742
rect 2486 3738 2490 3742
rect 2494 3738 2498 3742
rect 2710 3738 2714 3742
rect 3358 3738 3362 3742
rect 4758 3738 4762 3742
rect 5110 3738 5114 3742
rect 5190 3738 5194 3742
rect 134 3728 138 3732
rect 878 3728 882 3732
rect 926 3728 930 3732
rect 1934 3728 1938 3732
rect 2126 3728 2130 3732
rect 2158 3728 2162 3732
rect 2350 3728 2354 3732
rect 2782 3728 2786 3732
rect 2822 3728 2826 3732
rect 2862 3728 2866 3732
rect 2942 3728 2946 3732
rect 3134 3728 3138 3732
rect 3294 3728 3298 3732
rect 3734 3728 3738 3732
rect 3766 3728 3770 3732
rect 3998 3728 4002 3732
rect 4350 3728 4354 3732
rect 5134 3728 5138 3732
rect 1662 3718 1666 3722
rect 1950 3718 1954 3722
rect 2270 3718 2274 3722
rect 2942 3718 2946 3722
rect 2982 3718 2986 3722
rect 3982 3718 3986 3722
rect 4958 3718 4962 3722
rect 2590 3708 2594 3712
rect 2654 3708 2658 3712
rect 2710 3708 2714 3712
rect 2926 3708 2930 3712
rect 3206 3708 3210 3712
rect 3534 3708 3538 3712
rect 3550 3708 3554 3712
rect 3894 3708 3898 3712
rect 3998 3708 4002 3712
rect 4014 3708 4018 3712
rect 4774 3708 4778 3712
rect 5166 3708 5170 3712
rect 850 3703 854 3707
rect 858 3703 861 3707
rect 861 3703 862 3707
rect 1874 3703 1878 3707
rect 1882 3703 1885 3707
rect 1885 3703 1886 3707
rect 1110 3698 1114 3702
rect 2070 3698 2074 3702
rect 2094 3698 2098 3702
rect 2102 3698 2106 3702
rect 2890 3703 2894 3707
rect 2898 3703 2901 3707
rect 2901 3703 2902 3707
rect 3922 3703 3926 3707
rect 3930 3703 3933 3707
rect 3933 3703 3934 3707
rect 4938 3703 4942 3707
rect 4946 3703 4949 3707
rect 4949 3703 4950 3707
rect 2254 3698 2258 3702
rect 2726 3698 2730 3702
rect 2782 3698 2786 3702
rect 2814 3698 2818 3702
rect 2998 3698 3002 3702
rect 3454 3698 3458 3702
rect 3758 3698 3762 3702
rect 4190 3698 4194 3702
rect 5126 3698 5130 3702
rect 2110 3688 2114 3692
rect 2414 3688 2418 3692
rect 2654 3688 2658 3692
rect 3334 3688 3338 3692
rect 3598 3688 3602 3692
rect 3942 3688 3946 3692
rect 4214 3688 4218 3692
rect 4358 3688 4362 3692
rect 4950 3688 4954 3692
rect 4958 3688 4962 3692
rect 206 3678 210 3682
rect 982 3678 986 3682
rect 1350 3678 1354 3682
rect 1374 3678 1378 3682
rect 1838 3678 1842 3682
rect 1862 3678 1866 3682
rect 2190 3678 2194 3682
rect 2206 3678 2210 3682
rect 2414 3678 2418 3682
rect 2438 3678 2442 3682
rect 2846 3678 2850 3682
rect 2974 3678 2978 3682
rect 3030 3678 3034 3682
rect 3894 3678 3898 3682
rect 5118 3678 5122 3682
rect 5174 3678 5178 3682
rect 5278 3678 5282 3682
rect 118 3668 122 3672
rect 846 3668 850 3672
rect 1118 3668 1122 3672
rect 1214 3668 1218 3672
rect 1238 3668 1242 3672
rect 1486 3668 1490 3672
rect 1590 3668 1594 3672
rect 3134 3668 3138 3672
rect 3238 3668 3242 3672
rect 3278 3668 3282 3672
rect 3350 3668 3354 3672
rect 3510 3668 3514 3672
rect 3662 3668 3666 3672
rect 4166 3668 4170 3672
rect 4630 3668 4634 3672
rect 630 3658 634 3662
rect 710 3658 714 3662
rect 750 3658 754 3662
rect 1590 3658 1594 3662
rect 2054 3658 2058 3662
rect 2438 3658 2442 3662
rect 2686 3658 2690 3662
rect 2758 3658 2762 3662
rect 510 3648 514 3652
rect 630 3648 634 3652
rect 1174 3648 1178 3652
rect 1238 3648 1242 3652
rect 1318 3648 1322 3652
rect 1550 3648 1554 3652
rect 1798 3648 1802 3652
rect 2230 3648 2234 3652
rect 2446 3648 2450 3652
rect 2950 3658 2954 3662
rect 3030 3658 3034 3662
rect 3046 3658 3050 3662
rect 3214 3658 3218 3662
rect 3310 3658 3314 3662
rect 3558 3658 3562 3662
rect 3702 3658 3706 3662
rect 4006 3658 4010 3662
rect 4094 3658 4098 3662
rect 4278 3658 4282 3662
rect 4366 3658 4370 3662
rect 4398 3658 4402 3662
rect 4606 3658 4610 3662
rect 4774 3658 4778 3662
rect 4910 3658 4914 3662
rect 5038 3658 5042 3662
rect 5198 3658 5202 3662
rect 2934 3648 2938 3652
rect 2942 3648 2946 3652
rect 4254 3648 4258 3652
rect 1094 3638 1098 3642
rect 1494 3638 1498 3642
rect 1630 3638 1634 3642
rect 2678 3638 2682 3642
rect 2846 3638 2850 3642
rect 2854 3638 2858 3642
rect 2982 3638 2986 3642
rect 3422 3638 3426 3642
rect 3534 3638 3538 3642
rect 4198 3638 4202 3642
rect 4206 3638 4210 3642
rect 4374 3638 4378 3642
rect 4670 3638 4674 3642
rect 4694 3638 4698 3642
rect 4886 3638 4890 3642
rect 5270 3638 5274 3642
rect 1126 3628 1130 3632
rect 1174 3628 1178 3632
rect 1694 3628 1698 3632
rect 1798 3628 1802 3632
rect 2342 3628 2346 3632
rect 2974 3628 2978 3632
rect 3326 3628 3330 3632
rect 4222 3628 4226 3632
rect 4310 3628 4314 3632
rect 294 3618 298 3622
rect 1102 3618 1106 3622
rect 2102 3618 2106 3622
rect 3166 3618 3170 3622
rect 4086 3618 4090 3622
rect 4174 3618 4178 3622
rect 5046 3618 5050 3622
rect 646 3608 650 3612
rect 1334 3608 1338 3612
rect 2606 3608 2610 3612
rect 2734 3608 2738 3612
rect 2758 3608 2762 3612
rect 2934 3608 2938 3612
rect 3214 3608 3218 3612
rect 3638 3608 3642 3612
rect 4414 3608 4418 3612
rect 330 3603 334 3607
rect 338 3603 341 3607
rect 341 3603 342 3607
rect 1354 3603 1358 3607
rect 1362 3603 1365 3607
rect 1365 3603 1366 3607
rect 2386 3603 2390 3607
rect 2394 3603 2397 3607
rect 2397 3603 2398 3607
rect 3402 3603 3406 3607
rect 3410 3603 3413 3607
rect 3413 3603 3414 3607
rect 4426 3603 4430 3607
rect 4434 3603 4437 3607
rect 4437 3603 4438 3607
rect 974 3598 978 3602
rect 918 3588 922 3592
rect 1038 3588 1042 3592
rect 1270 3588 1274 3592
rect 1734 3588 1738 3592
rect 1838 3588 1842 3592
rect 2286 3588 2290 3592
rect 2606 3588 2610 3592
rect 3190 3588 3194 3592
rect 3550 3588 3554 3592
rect 3694 3588 3698 3592
rect 3990 3588 3994 3592
rect 4446 3588 4450 3592
rect 206 3578 210 3582
rect 502 3578 506 3582
rect 734 3578 738 3582
rect 870 3578 874 3582
rect 1014 3578 1018 3582
rect 1670 3578 1674 3582
rect 1830 3578 1834 3582
rect 2254 3578 2258 3582
rect 2670 3578 2674 3582
rect 2838 3578 2842 3582
rect 3278 3578 3282 3582
rect 4566 3578 4570 3582
rect 5006 3578 5010 3582
rect 462 3568 466 3572
rect 2478 3568 2482 3572
rect 2502 3568 2506 3572
rect 2574 3568 2578 3572
rect 3118 3568 3122 3572
rect 3678 3568 3682 3572
rect 4006 3568 4010 3572
rect 4014 3568 4018 3572
rect 4582 3568 4586 3572
rect 150 3558 154 3562
rect 406 3558 410 3562
rect 782 3558 786 3562
rect 822 3558 826 3562
rect 1174 3558 1178 3562
rect 1526 3558 1530 3562
rect 1782 3558 1786 3562
rect 2246 3558 2250 3562
rect 2726 3558 2730 3562
rect 2950 3558 2954 3562
rect 3294 3558 3298 3562
rect 3462 3558 3466 3562
rect 3702 3558 3706 3562
rect 3734 3558 3738 3562
rect 3758 3558 3762 3562
rect 4062 3558 4066 3562
rect 4278 3558 4282 3562
rect 4334 3558 4338 3562
rect 5174 3558 5178 3562
rect 5238 3558 5242 3562
rect 5270 3558 5274 3562
rect 622 3548 626 3552
rect 638 3548 642 3552
rect 830 3548 834 3552
rect 1054 3548 1058 3552
rect 1478 3548 1482 3552
rect 1486 3548 1490 3552
rect 1582 3548 1586 3552
rect 1614 3548 1618 3552
rect 1646 3548 1650 3552
rect 1662 3548 1666 3552
rect 1694 3548 1698 3552
rect 1766 3548 1770 3552
rect 1790 3548 1794 3552
rect 1822 3548 1826 3552
rect 2166 3548 2170 3552
rect 2342 3548 2346 3552
rect 846 3538 850 3542
rect 862 3538 866 3542
rect 1014 3538 1018 3542
rect 1278 3538 1282 3542
rect 1446 3538 1450 3542
rect 2062 3538 2066 3542
rect 2150 3538 2154 3542
rect 3318 3548 3322 3552
rect 3494 3548 3498 3552
rect 3526 3548 3530 3552
rect 4070 3548 4074 3552
rect 4158 3548 4162 3552
rect 4310 3548 4314 3552
rect 4366 3548 4370 3552
rect 4398 3548 4402 3552
rect 4526 3548 4530 3552
rect 4638 3548 4642 3552
rect 4662 3548 4666 3552
rect 4926 3548 4930 3552
rect 4966 3548 4970 3552
rect 2406 3538 2410 3542
rect 2510 3538 2514 3542
rect 2590 3538 2594 3542
rect 2710 3538 2714 3542
rect 2910 3538 2914 3542
rect 2966 3538 2970 3542
rect 3022 3538 3026 3542
rect 3150 3538 3154 3542
rect 3166 3538 3170 3542
rect 3230 3538 3234 3542
rect 3254 3538 3258 3542
rect 3286 3538 3290 3542
rect 4206 3538 4210 3542
rect 4470 3538 4474 3542
rect 4822 3538 4826 3542
rect 5174 3538 5178 3542
rect 5294 3538 5298 3542
rect 462 3528 466 3532
rect 558 3528 562 3532
rect 590 3528 594 3532
rect 1182 3528 1186 3532
rect 1622 3528 1626 3532
rect 1750 3528 1754 3532
rect 2038 3528 2042 3532
rect 2350 3528 2354 3532
rect 2862 3528 2866 3532
rect 3382 3528 3386 3532
rect 3438 3528 3442 3532
rect 3694 3528 3698 3532
rect 3806 3528 3810 3532
rect 3942 3528 3946 3532
rect 4030 3528 4034 3532
rect 4190 3528 4194 3532
rect 4286 3528 4290 3532
rect 4318 3528 4322 3532
rect 4382 3528 4386 3532
rect 4494 3528 4498 3532
rect 4502 3528 4506 3532
rect 5278 3528 5282 3532
rect 654 3518 658 3522
rect 1534 3518 1538 3522
rect 2206 3518 2210 3522
rect 3094 3518 3098 3522
rect 3198 3518 3202 3522
rect 3214 3518 3218 3522
rect 3310 3518 3314 3522
rect 3318 3518 3322 3522
rect 3678 3518 3682 3522
rect 4158 3518 4162 3522
rect 4206 3518 4210 3522
rect 5198 3518 5202 3522
rect 5246 3518 5250 3522
rect 638 3508 642 3512
rect 1438 3508 1442 3512
rect 1446 3508 1450 3512
rect 1606 3508 1610 3512
rect 1614 3508 1618 3512
rect 1774 3508 1778 3512
rect 2326 3508 2330 3512
rect 2910 3508 2914 3512
rect 3430 3508 3434 3512
rect 3966 3508 3970 3512
rect 4558 3508 4562 3512
rect 5246 3508 5250 3512
rect 850 3503 854 3507
rect 858 3503 861 3507
rect 861 3503 862 3507
rect 1874 3503 1878 3507
rect 1882 3503 1885 3507
rect 1885 3503 1886 3507
rect 2890 3503 2894 3507
rect 2898 3503 2901 3507
rect 2901 3503 2902 3507
rect 3922 3503 3926 3507
rect 3930 3503 3933 3507
rect 3933 3503 3934 3507
rect 4938 3503 4942 3507
rect 4946 3503 4949 3507
rect 4949 3503 4950 3507
rect 390 3498 394 3502
rect 1582 3498 1586 3502
rect 2230 3498 2234 3502
rect 2334 3498 2338 3502
rect 2766 3498 2770 3502
rect 3206 3498 3210 3502
rect 3502 3498 3506 3502
rect 3518 3498 3522 3502
rect 3958 3498 3962 3502
rect 4310 3498 4314 3502
rect 398 3488 402 3492
rect 1302 3488 1306 3492
rect 1334 3488 1338 3492
rect 1422 3488 1426 3492
rect 1606 3488 1610 3492
rect 2318 3488 2322 3492
rect 2374 3488 2378 3492
rect 2726 3488 2730 3492
rect 3486 3488 3490 3492
rect 3718 3488 3722 3492
rect 4054 3488 4058 3492
rect 4742 3488 4746 3492
rect 5038 3488 5042 3492
rect 510 3478 514 3482
rect 822 3478 826 3482
rect 966 3478 970 3482
rect 1342 3478 1346 3482
rect 1438 3478 1442 3482
rect 1590 3478 1594 3482
rect 2134 3478 2138 3482
rect 2822 3478 2826 3482
rect 3174 3478 3178 3482
rect 3278 3478 3282 3482
rect 3566 3478 3570 3482
rect 3694 3478 3698 3482
rect 3774 3478 3778 3482
rect 3998 3478 4002 3482
rect 894 3468 898 3472
rect 982 3468 986 3472
rect 1206 3468 1210 3472
rect 1270 3468 1274 3472
rect 1534 3468 1538 3472
rect 30 3458 34 3462
rect 1798 3468 1802 3472
rect 2182 3468 2186 3472
rect 2686 3468 2690 3472
rect 2982 3468 2986 3472
rect 3182 3468 3186 3472
rect 3574 3468 3578 3472
rect 3726 3468 3730 3472
rect 4046 3468 4050 3472
rect 4470 3468 4474 3472
rect 4998 3468 5002 3472
rect 510 3458 514 3462
rect 830 3458 834 3462
rect 910 3458 914 3462
rect 1278 3458 1282 3462
rect 1454 3458 1458 3462
rect 1742 3458 1746 3462
rect 1790 3458 1794 3462
rect 1814 3458 1818 3462
rect 1846 3458 1850 3462
rect 2830 3458 2834 3462
rect 3142 3458 3146 3462
rect 3198 3458 3202 3462
rect 3486 3458 3490 3462
rect 3750 3458 3754 3462
rect 4310 3458 4314 3462
rect 4518 3458 4522 3462
rect 4598 3458 4602 3462
rect 4614 3458 4618 3462
rect 4654 3458 4658 3462
rect 4678 3458 4682 3462
rect 4686 3458 4690 3462
rect 5126 3458 5130 3462
rect 5238 3458 5242 3462
rect 710 3448 714 3452
rect 1270 3448 1274 3452
rect 1342 3448 1346 3452
rect 1494 3448 1498 3452
rect 2702 3448 2706 3452
rect 3150 3448 3154 3452
rect 3230 3448 3234 3452
rect 4006 3448 4010 3452
rect 4486 3448 4490 3452
rect 4678 3448 4682 3452
rect 4958 3448 4962 3452
rect 1086 3438 1090 3442
rect 1198 3438 1202 3442
rect 1518 3438 1522 3442
rect 2014 3438 2018 3442
rect 3086 3438 3090 3442
rect 4654 3438 4658 3442
rect 5094 3438 5098 3442
rect 5134 3438 5138 3442
rect 1166 3428 1170 3432
rect 2318 3428 2322 3432
rect 4094 3428 4098 3432
rect 4142 3428 4146 3432
rect 4190 3428 4194 3432
rect 4790 3428 4794 3432
rect 782 3418 786 3422
rect 3302 3418 3306 3422
rect 3510 3418 3514 3422
rect 3590 3418 3594 3422
rect 4190 3418 4194 3422
rect 4510 3418 4514 3422
rect 4630 3418 4634 3422
rect 5230 3418 5234 3422
rect 2246 3408 2250 3412
rect 2366 3408 2370 3412
rect 2790 3408 2794 3412
rect 3062 3408 3066 3412
rect 3174 3408 3178 3412
rect 3446 3408 3450 3412
rect 3598 3408 3602 3412
rect 4470 3408 4474 3412
rect 4982 3408 4986 3412
rect 330 3403 334 3407
rect 338 3403 341 3407
rect 341 3403 342 3407
rect 1354 3403 1358 3407
rect 1362 3403 1365 3407
rect 1365 3403 1366 3407
rect 2386 3403 2390 3407
rect 2394 3403 2397 3407
rect 2397 3403 2398 3407
rect 3402 3403 3406 3407
rect 3410 3403 3413 3407
rect 3413 3403 3414 3407
rect 4426 3403 4430 3407
rect 4434 3403 4437 3407
rect 4437 3403 4438 3407
rect 1750 3398 1754 3402
rect 2030 3398 2034 3402
rect 2694 3398 2698 3402
rect 3214 3398 3218 3402
rect 4702 3398 4706 3402
rect 4982 3398 4986 3402
rect 4990 3398 4994 3402
rect 2966 3388 2970 3392
rect 3518 3388 3522 3392
rect 3542 3388 3546 3392
rect 4758 3388 4762 3392
rect 1294 3378 1298 3382
rect 1766 3378 1770 3382
rect 1806 3378 1810 3382
rect 2878 3378 2882 3382
rect 4550 3378 4554 3382
rect 4662 3378 4666 3382
rect 5046 3378 5050 3382
rect 502 3368 506 3372
rect 1494 3368 1498 3372
rect 2022 3368 2026 3372
rect 2134 3368 2138 3372
rect 2638 3368 2642 3372
rect 2670 3368 2674 3372
rect 2974 3368 2978 3372
rect 3054 3368 3058 3372
rect 3158 3368 3162 3372
rect 3214 3368 3218 3372
rect 4478 3368 4482 3372
rect 4926 3368 4930 3372
rect 430 3358 434 3362
rect 558 3358 562 3362
rect 878 3358 882 3362
rect 1150 3358 1154 3362
rect 1486 3358 1490 3362
rect 1774 3358 1778 3362
rect 2134 3358 2138 3362
rect 2166 3358 2170 3362
rect 2934 3358 2938 3362
rect 3422 3358 3426 3362
rect 3574 3358 3578 3362
rect 4462 3358 4466 3362
rect 4486 3358 4490 3362
rect 4518 3358 4522 3362
rect 4726 3358 4730 3362
rect 4854 3358 4858 3362
rect 5126 3358 5130 3362
rect 1958 3348 1962 3352
rect 2166 3348 2170 3352
rect 2438 3348 2442 3352
rect 2518 3348 2522 3352
rect 2670 3348 2674 3352
rect 3278 3348 3282 3352
rect 3902 3348 3906 3352
rect 4830 3348 4834 3352
rect 134 3338 138 3342
rect 630 3338 634 3342
rect 806 3338 810 3342
rect 830 3338 834 3342
rect 878 3338 882 3342
rect 1142 3338 1146 3342
rect 1318 3338 1322 3342
rect 1598 3338 1602 3342
rect 1782 3338 1786 3342
rect 2070 3338 2074 3342
rect 2094 3338 2098 3342
rect 2118 3338 2122 3342
rect 2614 3338 2618 3342
rect 2910 3338 2914 3342
rect 3038 3338 3042 3342
rect 3054 3338 3058 3342
rect 3358 3338 3362 3342
rect 3606 3338 3610 3342
rect 3718 3338 3722 3342
rect 4070 3338 4074 3342
rect 4374 3338 4378 3342
rect 4494 3338 4498 3342
rect 5134 3338 5138 3342
rect 590 3328 594 3332
rect 630 3328 634 3332
rect 806 3328 810 3332
rect 886 3328 890 3332
rect 1150 3328 1154 3332
rect 1486 3328 1490 3332
rect 1934 3328 1938 3332
rect 302 3318 306 3322
rect 582 3318 586 3322
rect 646 3318 650 3322
rect 742 3318 746 3322
rect 1566 3318 1570 3322
rect 2710 3328 2714 3332
rect 3214 3328 3218 3332
rect 3390 3328 3394 3332
rect 3678 3328 3682 3332
rect 3790 3328 3794 3332
rect 4214 3328 4218 3332
rect 2318 3318 2322 3322
rect 2614 3318 2618 3322
rect 3686 3318 3690 3322
rect 4102 3318 4106 3322
rect 4574 3318 4578 3322
rect 590 3308 594 3312
rect 734 3308 738 3312
rect 806 3308 810 3312
rect 1542 3308 1546 3312
rect 1574 3308 1578 3312
rect 1590 3308 1594 3312
rect 2110 3308 2114 3312
rect 2342 3308 2346 3312
rect 2598 3308 2602 3312
rect 2742 3308 2746 3312
rect 2838 3308 2842 3312
rect 3166 3308 3170 3312
rect 3734 3308 3738 3312
rect 3982 3308 3986 3312
rect 850 3303 854 3307
rect 858 3303 861 3307
rect 861 3303 862 3307
rect 1874 3303 1878 3307
rect 1882 3303 1885 3307
rect 1885 3303 1886 3307
rect 2890 3303 2894 3307
rect 2898 3303 2901 3307
rect 2901 3303 2902 3307
rect 3922 3303 3926 3307
rect 3930 3303 3933 3307
rect 3933 3303 3934 3307
rect 4938 3303 4942 3307
rect 4946 3303 4949 3307
rect 4949 3303 4950 3307
rect 2254 3298 2258 3302
rect 2734 3298 2738 3302
rect 2942 3298 2946 3302
rect 3374 3298 3378 3302
rect 4838 3298 4842 3302
rect 1942 3288 1946 3292
rect 2270 3288 2274 3292
rect 2566 3288 2570 3292
rect 2830 3288 2834 3292
rect 3334 3288 3338 3292
rect 3502 3288 3506 3292
rect 3710 3288 3714 3292
rect 4886 3288 4890 3292
rect 102 3278 106 3282
rect 446 3278 450 3282
rect 766 3278 770 3282
rect 878 3278 882 3282
rect 1174 3278 1178 3282
rect 1486 3278 1490 3282
rect 1742 3278 1746 3282
rect 2062 3278 2066 3282
rect 2446 3278 2450 3282
rect 2718 3278 2722 3282
rect 2726 3278 2730 3282
rect 2782 3278 2786 3282
rect 3350 3278 3354 3282
rect 4310 3278 4314 3282
rect 4846 3278 4850 3282
rect 4910 3278 4914 3282
rect 758 3268 762 3272
rect 1334 3268 1338 3272
rect 1430 3268 1434 3272
rect 1814 3268 1818 3272
rect 2182 3268 2186 3272
rect 2542 3268 2546 3272
rect 2734 3268 2738 3272
rect 3134 3268 3138 3272
rect 3294 3268 3298 3272
rect 3726 3268 3730 3272
rect 4030 3268 4034 3272
rect 4086 3268 4090 3272
rect 4334 3268 4338 3272
rect 4454 3268 4458 3272
rect 4494 3268 4498 3272
rect 4510 3268 4514 3272
rect 4798 3268 4802 3272
rect 4878 3268 4882 3272
rect 5214 3268 5218 3272
rect 5294 3268 5298 3272
rect 470 3258 474 3262
rect 734 3258 738 3262
rect 918 3258 922 3262
rect 1158 3258 1162 3262
rect 1286 3258 1290 3262
rect 1526 3258 1530 3262
rect 2038 3258 2042 3262
rect 2478 3258 2482 3262
rect 2494 3258 2498 3262
rect 2742 3258 2746 3262
rect 3526 3258 3530 3262
rect 4062 3258 4066 3262
rect 4158 3258 4162 3262
rect 4486 3258 4490 3262
rect 4526 3258 4530 3262
rect 4582 3258 4586 3262
rect 4814 3258 4818 3262
rect 5294 3258 5298 3262
rect 990 3248 994 3252
rect 1454 3248 1458 3252
rect 1478 3248 1482 3252
rect 1526 3248 1530 3252
rect 1582 3248 1586 3252
rect 1606 3248 1610 3252
rect 1614 3248 1618 3252
rect 2478 3248 2482 3252
rect 2806 3248 2810 3252
rect 2830 3248 2834 3252
rect 2854 3248 2858 3252
rect 3862 3248 3866 3252
rect 4214 3248 4218 3252
rect 4534 3248 4538 3252
rect 4838 3248 4842 3252
rect 4870 3248 4874 3252
rect 670 3238 674 3242
rect 1502 3238 1506 3242
rect 2022 3238 2026 3242
rect 2102 3238 2106 3242
rect 2686 3238 2690 3242
rect 2758 3238 2762 3242
rect 2774 3238 2778 3242
rect 2894 3238 2898 3242
rect 2966 3238 2970 3242
rect 3302 3238 3306 3242
rect 3558 3238 3562 3242
rect 3814 3238 3818 3242
rect 4270 3238 4274 3242
rect 4558 3238 4562 3242
rect 4862 3238 4866 3242
rect 4870 3238 4874 3242
rect 726 3228 730 3232
rect 1510 3228 1514 3232
rect 2678 3228 2682 3232
rect 2718 3228 2722 3232
rect 2766 3228 2770 3232
rect 3190 3228 3194 3232
rect 3606 3228 3610 3232
rect 4198 3228 4202 3232
rect 5038 3228 5042 3232
rect 966 3218 970 3222
rect 1710 3218 1714 3222
rect 1998 3218 2002 3222
rect 2070 3218 2074 3222
rect 2102 3218 2106 3222
rect 2710 3218 2714 3222
rect 4558 3218 4562 3222
rect 718 3208 722 3212
rect 926 3208 930 3212
rect 2254 3208 2258 3212
rect 2310 3208 2314 3212
rect 2550 3208 2554 3212
rect 4110 3208 4114 3212
rect 4366 3208 4370 3212
rect 5102 3208 5106 3212
rect 5134 3208 5138 3212
rect 330 3203 334 3207
rect 338 3203 341 3207
rect 341 3203 342 3207
rect 1354 3203 1358 3207
rect 1362 3203 1365 3207
rect 1365 3203 1366 3207
rect 2386 3203 2390 3207
rect 2394 3203 2397 3207
rect 2397 3203 2398 3207
rect 3402 3203 3406 3207
rect 3410 3203 3413 3207
rect 3413 3203 3414 3207
rect 4426 3203 4430 3207
rect 4434 3203 4437 3207
rect 4437 3203 4438 3207
rect 894 3198 898 3202
rect 942 3198 946 3202
rect 1654 3198 1658 3202
rect 2190 3198 2194 3202
rect 3134 3198 3138 3202
rect 4518 3198 4522 3202
rect 4870 3198 4874 3202
rect 4990 3198 4994 3202
rect 1262 3188 1266 3192
rect 1590 3188 1594 3192
rect 2782 3188 2786 3192
rect 3078 3188 3082 3192
rect 3382 3188 3386 3192
rect 4118 3188 4122 3192
rect 4182 3188 4186 3192
rect 4326 3188 4330 3192
rect 4790 3188 4794 3192
rect 1478 3178 1482 3182
rect 2046 3178 2050 3182
rect 2694 3178 2698 3182
rect 2950 3178 2954 3182
rect 3038 3178 3042 3182
rect 3158 3178 3162 3182
rect 3790 3178 3794 3182
rect 1374 3168 1378 3172
rect 4526 3178 4530 3182
rect 1398 3168 1402 3172
rect 1454 3168 1458 3172
rect 1734 3168 1738 3172
rect 2486 3168 2490 3172
rect 3606 3168 3610 3172
rect 3742 3168 3746 3172
rect 4134 3168 4138 3172
rect 4342 3168 4346 3172
rect 4518 3168 4522 3172
rect 4566 3168 4570 3172
rect 638 3158 642 3162
rect 1166 3158 1170 3162
rect 1190 3158 1194 3162
rect 1494 3158 1498 3162
rect 2438 3158 2442 3162
rect 2486 3158 2490 3162
rect 2622 3158 2626 3162
rect 2822 3158 2826 3162
rect 2838 3158 2842 3162
rect 3446 3158 3450 3162
rect 4150 3158 4154 3162
rect 294 3148 298 3152
rect 654 3148 658 3152
rect 686 3148 690 3152
rect 710 3148 714 3152
rect 726 3148 730 3152
rect 798 3148 802 3152
rect 1054 3148 1058 3152
rect 1174 3148 1178 3152
rect 1542 3148 1546 3152
rect 1622 3148 1626 3152
rect 1670 3148 1674 3152
rect 1694 3148 1698 3152
rect 1838 3148 1842 3152
rect 1966 3148 1970 3152
rect 2110 3148 2114 3152
rect 2270 3148 2274 3152
rect 2550 3148 2554 3152
rect 2654 3148 2658 3152
rect 2934 3148 2938 3152
rect 3030 3148 3034 3152
rect 4558 3158 4562 3162
rect 4606 3158 4610 3162
rect 4822 3158 4826 3162
rect 4886 3158 4890 3162
rect 4910 3158 4914 3162
rect 3150 3148 3154 3152
rect 3198 3148 3202 3152
rect 3678 3148 3682 3152
rect 3734 3148 3738 3152
rect 3846 3148 3850 3152
rect 3894 3148 3898 3152
rect 4062 3148 4066 3152
rect 4126 3148 4130 3152
rect 4414 3148 4418 3152
rect 4446 3148 4450 3152
rect 4526 3148 4530 3152
rect 4534 3148 4538 3152
rect 4574 3148 4578 3152
rect 4726 3148 4730 3152
rect 4870 3148 4874 3152
rect 5118 3148 5122 3152
rect 726 3138 730 3142
rect 734 3138 738 3142
rect 1174 3138 1178 3142
rect 1214 3138 1218 3142
rect 1566 3138 1570 3142
rect 1622 3138 1626 3142
rect 1646 3138 1650 3142
rect 1686 3138 1690 3142
rect 2238 3138 2242 3142
rect 2278 3138 2282 3142
rect 2310 3138 2314 3142
rect 2630 3138 2634 3142
rect 2678 3138 2682 3142
rect 2822 3138 2826 3142
rect 2942 3138 2946 3142
rect 2998 3138 3002 3142
rect 3110 3138 3114 3142
rect 4742 3138 4746 3142
rect 4758 3138 4762 3142
rect 4798 3138 4802 3142
rect 4862 3138 4866 3142
rect 598 3128 602 3132
rect 798 3128 802 3132
rect 822 3128 826 3132
rect 846 3128 850 3132
rect 1126 3128 1130 3132
rect 1398 3128 1402 3132
rect 1462 3128 1466 3132
rect 1478 3128 1482 3132
rect 1782 3128 1786 3132
rect 2350 3128 2354 3132
rect 2478 3128 2482 3132
rect 2854 3128 2858 3132
rect 3054 3128 3058 3132
rect 3166 3128 3170 3132
rect 4414 3128 4418 3132
rect 5014 3128 5018 3132
rect 5198 3128 5202 3132
rect 5230 3128 5234 3132
rect 582 3118 586 3122
rect 734 3118 738 3122
rect 742 3118 746 3122
rect 1462 3118 1466 3122
rect 1926 3118 1930 3122
rect 2022 3118 2026 3122
rect 2342 3118 2346 3122
rect 2558 3118 2562 3122
rect 2686 3118 2690 3122
rect 3150 3118 3154 3122
rect 3430 3118 3434 3122
rect 4518 3118 4522 3122
rect 614 3108 618 3112
rect 678 3108 682 3112
rect 1238 3108 1242 3112
rect 1438 3108 1442 3112
rect 1622 3108 1626 3112
rect 2646 3108 2650 3112
rect 3470 3108 3474 3112
rect 3630 3108 3634 3112
rect 4062 3108 4066 3112
rect 4086 3108 4090 3112
rect 4758 3108 4762 3112
rect 850 3103 854 3107
rect 858 3103 861 3107
rect 861 3103 862 3107
rect 366 3098 370 3102
rect 838 3098 842 3102
rect 1470 3098 1474 3102
rect 1874 3103 1878 3107
rect 1882 3103 1885 3107
rect 1885 3103 1886 3107
rect 1894 3098 1898 3102
rect 2126 3098 2130 3102
rect 2486 3098 2490 3102
rect 2494 3098 2498 3102
rect 2890 3103 2894 3107
rect 2898 3103 2901 3107
rect 2901 3103 2902 3107
rect 3922 3103 3926 3107
rect 3930 3103 3933 3107
rect 3933 3103 3934 3107
rect 4938 3103 4942 3107
rect 4946 3103 4949 3107
rect 4949 3103 4950 3107
rect 2878 3098 2882 3102
rect 2918 3098 2922 3102
rect 2942 3098 2946 3102
rect 3174 3098 3178 3102
rect 3942 3098 3946 3102
rect 4462 3098 4466 3102
rect 4470 3098 4474 3102
rect 5110 3098 5114 3102
rect 1206 3088 1210 3092
rect 1382 3088 1386 3092
rect 2158 3088 2162 3092
rect 3430 3088 3434 3092
rect 606 3078 610 3082
rect 1374 3078 1378 3082
rect 4022 3088 4026 3092
rect 4262 3088 4266 3092
rect 4630 3088 4634 3092
rect 4910 3088 4914 3092
rect 5230 3088 5234 3092
rect 1542 3078 1546 3082
rect 1566 3078 1570 3082
rect 1622 3078 1626 3082
rect 1670 3078 1674 3082
rect 1718 3078 1722 3082
rect 1894 3078 1898 3082
rect 1982 3078 1986 3082
rect 2126 3078 2130 3082
rect 2838 3078 2842 3082
rect 3126 3078 3130 3082
rect 3238 3078 3242 3082
rect 3662 3078 3666 3082
rect 4310 3078 4314 3082
rect 4358 3078 4362 3082
rect 4374 3078 4378 3082
rect 4574 3078 4578 3082
rect 670 3068 674 3072
rect 990 3068 994 3072
rect 1326 3068 1330 3072
rect 1334 3068 1338 3072
rect 1638 3068 1642 3072
rect 1654 3068 1658 3072
rect 1838 3068 1842 3072
rect 1870 3068 1874 3072
rect 2358 3068 2362 3072
rect 2558 3068 2562 3072
rect 2630 3068 2634 3072
rect 3038 3068 3042 3072
rect 3086 3068 3090 3072
rect 3430 3068 3434 3072
rect 3678 3068 3682 3072
rect 3694 3068 3698 3072
rect 3862 3068 3866 3072
rect 3902 3068 3906 3072
rect 3942 3068 3946 3072
rect 4174 3068 4178 3072
rect 158 3058 162 3062
rect 198 3058 202 3062
rect 558 3058 562 3062
rect 1198 3058 1202 3062
rect 1222 3058 1226 3062
rect 1446 3058 1450 3062
rect 1486 3058 1490 3062
rect 1646 3058 1650 3062
rect 1862 3058 1866 3062
rect 2510 3058 2514 3062
rect 2598 3058 2602 3062
rect 2654 3058 2658 3062
rect 2830 3058 2834 3062
rect 3622 3058 3626 3062
rect 3646 3058 3650 3062
rect 3742 3058 3746 3062
rect 3910 3058 3914 3062
rect 4022 3058 4026 3062
rect 4038 3058 4042 3062
rect 4150 3058 4154 3062
rect 1374 3048 1378 3052
rect 1382 3048 1386 3052
rect 1446 3048 1450 3052
rect 1598 3048 1602 3052
rect 4262 3058 4266 3062
rect 4374 3058 4378 3062
rect 4606 3058 4610 3062
rect 4702 3058 4706 3062
rect 4958 3058 4962 3062
rect 1862 3048 1866 3052
rect 1894 3048 1898 3052
rect 1902 3048 1906 3052
rect 2502 3048 2506 3052
rect 2526 3048 2530 3052
rect 2542 3048 2546 3052
rect 2790 3048 2794 3052
rect 2934 3048 2938 3052
rect 3118 3048 3122 3052
rect 3150 3048 3154 3052
rect 3334 3048 3338 3052
rect 4254 3048 4258 3052
rect 4574 3048 4578 3052
rect 4646 3048 4650 3052
rect 4710 3048 4714 3052
rect 4758 3048 4762 3052
rect 4982 3048 4986 3052
rect 1582 3038 1586 3042
rect 1638 3038 1642 3042
rect 1894 3038 1898 3042
rect 2134 3038 2138 3042
rect 2310 3038 2314 3042
rect 2486 3038 2490 3042
rect 2990 3038 2994 3042
rect 3302 3038 3306 3042
rect 3382 3038 3386 3042
rect 1854 3028 1858 3032
rect 2918 3028 2922 3032
rect 3038 3028 3042 3032
rect 3046 3028 3050 3032
rect 3150 3028 3154 3032
rect 3358 3028 3362 3032
rect 4198 3028 4202 3032
rect 4398 3028 4402 3032
rect 4910 3028 4914 3032
rect 5190 3028 5194 3032
rect 1078 3018 1082 3022
rect 1598 3018 1602 3022
rect 1950 3018 1954 3022
rect 2718 3018 2722 3022
rect 3086 3018 3090 3022
rect 3390 3018 3394 3022
rect 3958 3018 3962 3022
rect 4142 3018 4146 3022
rect 4694 3018 4698 3022
rect 5110 3018 5114 3022
rect 5190 3018 5194 3022
rect 5230 3018 5234 3022
rect 1478 3008 1482 3012
rect 1742 3008 1746 3012
rect 1822 3008 1826 3012
rect 1910 3008 1914 3012
rect 2654 3008 2658 3012
rect 3198 3008 3202 3012
rect 4190 3008 4194 3012
rect 4406 3008 4410 3012
rect 4478 3008 4482 3012
rect 5022 3008 5026 3012
rect 5230 3008 5234 3012
rect 330 3003 334 3007
rect 338 3003 341 3007
rect 341 3003 342 3007
rect 1354 3003 1358 3007
rect 1362 3003 1365 3007
rect 1365 3003 1366 3007
rect 2386 3003 2390 3007
rect 2394 3003 2397 3007
rect 2397 3003 2398 3007
rect 3402 3003 3406 3007
rect 3410 3003 3413 3007
rect 3413 3003 3414 3007
rect 4426 3003 4430 3007
rect 4434 3003 4437 3007
rect 4437 3003 4438 3007
rect 1294 2998 1298 3002
rect 2366 2998 2370 3002
rect 2662 2998 2666 3002
rect 3030 2998 3034 3002
rect 3286 2998 3290 3002
rect 3302 2998 3306 3002
rect 4022 2998 4026 3002
rect 4166 2998 4170 3002
rect 286 2988 290 2992
rect 1206 2988 1210 2992
rect 1270 2988 1274 2992
rect 1702 2988 1706 2992
rect 2462 2988 2466 2992
rect 3062 2988 3066 2992
rect 3254 2988 3258 2992
rect 3886 2988 3890 2992
rect 3894 2988 3898 2992
rect 4582 2988 4586 2992
rect 5134 2988 5138 2992
rect 310 2978 314 2982
rect 638 2978 642 2982
rect 1062 2978 1066 2982
rect 1086 2978 1090 2982
rect 1622 2978 1626 2982
rect 3174 2978 3178 2982
rect 3206 2978 3210 2982
rect 3350 2978 3354 2982
rect 3582 2978 3586 2982
rect 3686 2978 3690 2982
rect 3702 2978 3706 2982
rect 4414 2978 4418 2982
rect 4702 2978 4706 2982
rect 518 2968 522 2972
rect 1534 2968 1538 2972
rect 3142 2968 3146 2972
rect 3310 2968 3314 2972
rect 3566 2968 3570 2972
rect 3798 2968 3802 2972
rect 4334 2968 4338 2972
rect 4390 2968 4394 2972
rect 4446 2968 4450 2972
rect 4662 2968 4666 2972
rect 4734 2968 4738 2972
rect 5134 2968 5138 2972
rect 2478 2958 2482 2962
rect 2518 2958 2522 2962
rect 3990 2958 3994 2962
rect 4078 2958 4082 2962
rect 4406 2958 4410 2962
rect 4422 2958 4426 2962
rect 4486 2958 4490 2962
rect 606 2948 610 2952
rect 662 2948 666 2952
rect 678 2948 682 2952
rect 718 2948 722 2952
rect 814 2948 818 2952
rect 910 2948 914 2952
rect 1030 2948 1034 2952
rect 1134 2948 1138 2952
rect 1166 2948 1170 2952
rect 1254 2948 1258 2952
rect 1654 2948 1658 2952
rect 1734 2948 1738 2952
rect 1806 2948 1810 2952
rect 1950 2948 1954 2952
rect 2254 2948 2258 2952
rect 2358 2948 2362 2952
rect 2414 2948 2418 2952
rect 2502 2948 2506 2952
rect 2990 2948 2994 2952
rect 2998 2948 3002 2952
rect 3382 2948 3386 2952
rect 3390 2948 3394 2952
rect 4046 2948 4050 2952
rect 4310 2948 4314 2952
rect 4350 2948 4354 2952
rect 4366 2948 4370 2952
rect 4390 2948 4394 2952
rect 4862 2948 4866 2952
rect 5150 2948 5154 2952
rect 5214 2948 5218 2952
rect 5294 2948 5298 2952
rect 1094 2938 1098 2942
rect 1262 2938 1266 2942
rect 1638 2938 1642 2942
rect 1822 2938 1826 2942
rect 1838 2938 1842 2942
rect 1974 2938 1978 2942
rect 2254 2938 2258 2942
rect 2534 2938 2538 2942
rect 2558 2938 2562 2942
rect 2582 2938 2586 2942
rect 2750 2938 2754 2942
rect 3030 2938 3034 2942
rect 3982 2938 3986 2942
rect 4174 2938 4178 2942
rect 4190 2938 4194 2942
rect 4302 2938 4306 2942
rect 4494 2938 4498 2942
rect 4510 2938 4514 2942
rect 4870 2938 4874 2942
rect 5038 2938 5042 2942
rect 5254 2938 5258 2942
rect 694 2928 698 2932
rect 1814 2928 1818 2932
rect 1830 2928 1834 2932
rect 2230 2928 2234 2932
rect 2486 2928 2490 2932
rect 2598 2928 2602 2932
rect 2606 2928 2610 2932
rect 3422 2928 3426 2932
rect 3430 2928 3434 2932
rect 3446 2928 3450 2932
rect 3638 2928 3642 2932
rect 4142 2928 4146 2932
rect 4318 2928 4322 2932
rect 4526 2928 4530 2932
rect 502 2918 506 2922
rect 638 2918 642 2922
rect 974 2918 978 2922
rect 1918 2918 1922 2922
rect 2750 2918 2754 2922
rect 3198 2918 3202 2922
rect 3230 2918 3234 2922
rect 3294 2918 3298 2922
rect 3646 2918 3650 2922
rect 4814 2918 4818 2922
rect 4854 2918 4858 2922
rect 4862 2918 4866 2922
rect 5006 2918 5010 2922
rect 454 2908 458 2912
rect 1766 2908 1770 2912
rect 1910 2908 1914 2912
rect 2198 2908 2202 2912
rect 3054 2908 3058 2912
rect 3326 2908 3330 2912
rect 3358 2908 3362 2912
rect 3902 2908 3906 2912
rect 4838 2908 4842 2912
rect 850 2903 854 2907
rect 858 2903 861 2907
rect 861 2903 862 2907
rect 814 2898 818 2902
rect 1874 2903 1878 2907
rect 1882 2903 1885 2907
rect 1885 2903 1886 2907
rect 2890 2903 2894 2907
rect 2898 2903 2901 2907
rect 2901 2903 2902 2907
rect 3922 2903 3926 2907
rect 3930 2903 3933 2907
rect 3933 2903 3934 2907
rect 4938 2903 4942 2907
rect 4946 2903 4949 2907
rect 4949 2903 4950 2907
rect 1262 2898 1266 2902
rect 1478 2898 1482 2902
rect 1710 2898 1714 2902
rect 1854 2898 1858 2902
rect 2574 2898 2578 2902
rect 2606 2898 2610 2902
rect 2910 2898 2914 2902
rect 3870 2898 3874 2902
rect 4654 2898 4658 2902
rect 4854 2898 4858 2902
rect 1046 2888 1050 2892
rect 1070 2888 1074 2892
rect 1334 2888 1338 2892
rect 2142 2888 2146 2892
rect 2294 2888 2298 2892
rect 2342 2888 2346 2892
rect 2582 2888 2586 2892
rect 2942 2888 2946 2892
rect 3030 2888 3034 2892
rect 4294 2888 4298 2892
rect 4950 2888 4954 2892
rect 5166 2888 5170 2892
rect 206 2878 210 2882
rect 614 2878 618 2882
rect 1590 2878 1594 2882
rect 1750 2878 1754 2882
rect 2430 2878 2434 2882
rect 2654 2878 2658 2882
rect 3654 2878 3658 2882
rect 3686 2878 3690 2882
rect 4286 2878 4290 2882
rect 110 2868 114 2872
rect 270 2868 274 2872
rect 526 2868 530 2872
rect 878 2868 882 2872
rect 1294 2868 1298 2872
rect 1310 2868 1314 2872
rect 1782 2868 1786 2872
rect 2030 2868 2034 2872
rect 2254 2868 2258 2872
rect 2302 2868 2306 2872
rect 3006 2868 3010 2872
rect 3206 2868 3210 2872
rect 4526 2868 4530 2872
rect 38 2858 42 2862
rect 142 2858 146 2862
rect 198 2858 202 2862
rect 558 2858 562 2862
rect 1054 2858 1058 2862
rect 1590 2858 1594 2862
rect 1766 2858 1770 2862
rect 2150 2858 2154 2862
rect 2582 2858 2586 2862
rect 2630 2858 2634 2862
rect 2654 2858 2658 2862
rect 3174 2858 3178 2862
rect 3542 2858 3546 2862
rect 4046 2858 4050 2862
rect 4190 2858 4194 2862
rect 4326 2858 4330 2862
rect 4486 2858 4490 2862
rect 4542 2858 4546 2862
rect 4830 2858 4834 2862
rect 4846 2858 4850 2862
rect 4886 2858 4890 2862
rect 5142 2858 5146 2862
rect 262 2848 266 2852
rect 518 2848 522 2852
rect 646 2848 650 2852
rect 734 2848 738 2852
rect 926 2848 930 2852
rect 1086 2848 1090 2852
rect 1102 2848 1106 2852
rect 1118 2848 1122 2852
rect 1286 2848 1290 2852
rect 1310 2848 1314 2852
rect 1566 2848 1570 2852
rect 2766 2848 2770 2852
rect 2926 2848 2930 2852
rect 3070 2848 3074 2852
rect 3142 2848 3146 2852
rect 3190 2848 3194 2852
rect 3262 2848 3266 2852
rect 3558 2848 3562 2852
rect 3830 2848 3834 2852
rect 4246 2848 4250 2852
rect 4790 2848 4794 2852
rect 5206 2848 5210 2852
rect 5222 2848 5226 2852
rect 246 2838 250 2842
rect 390 2838 394 2842
rect 510 2838 514 2842
rect 902 2838 906 2842
rect 1158 2838 1162 2842
rect 1942 2838 1946 2842
rect 2310 2838 2314 2842
rect 3366 2838 3370 2842
rect 3622 2838 3626 2842
rect 3854 2838 3858 2842
rect 4118 2838 4122 2842
rect 4718 2838 4722 2842
rect 5086 2838 5090 2842
rect 598 2828 602 2832
rect 822 2828 826 2832
rect 1134 2828 1138 2832
rect 1206 2828 1210 2832
rect 1686 2828 1690 2832
rect 2846 2828 2850 2832
rect 3166 2828 3170 2832
rect 3334 2828 3338 2832
rect 4206 2828 4210 2832
rect 4246 2828 4250 2832
rect 534 2818 538 2822
rect 686 2818 690 2822
rect 1542 2818 1546 2822
rect 2094 2818 2098 2822
rect 2470 2818 2474 2822
rect 2654 2818 2658 2822
rect 2686 2818 2690 2822
rect 3118 2818 3122 2822
rect 4134 2818 4138 2822
rect 5022 2818 5026 2822
rect 5198 2818 5202 2822
rect 5286 2818 5290 2822
rect 686 2808 690 2812
rect 1334 2808 1338 2812
rect 1742 2808 1746 2812
rect 2086 2808 2090 2812
rect 2134 2808 2138 2812
rect 2406 2808 2410 2812
rect 2534 2808 2538 2812
rect 3102 2808 3106 2812
rect 3966 2808 3970 2812
rect 330 2803 334 2807
rect 338 2803 341 2807
rect 341 2803 342 2807
rect 470 2798 474 2802
rect 1354 2803 1358 2807
rect 1362 2803 1365 2807
rect 1365 2803 1366 2807
rect 902 2798 906 2802
rect 1142 2798 1146 2802
rect 1214 2798 1218 2802
rect 2386 2803 2390 2807
rect 2394 2803 2397 2807
rect 2397 2803 2398 2807
rect 3402 2803 3406 2807
rect 3410 2803 3413 2807
rect 3413 2803 3414 2807
rect 1926 2798 1930 2802
rect 2502 2798 2506 2802
rect 2702 2798 2706 2802
rect 2966 2798 2970 2802
rect 3014 2798 3018 2802
rect 4426 2803 4430 2807
rect 4434 2803 4437 2807
rect 4437 2803 4438 2807
rect 3998 2798 4002 2802
rect 5174 2798 5178 2802
rect 702 2788 706 2792
rect 822 2788 826 2792
rect 1086 2788 1090 2792
rect 1598 2788 1602 2792
rect 2454 2788 2458 2792
rect 2958 2788 2962 2792
rect 2990 2788 2994 2792
rect 3286 2788 3290 2792
rect 4574 2788 4578 2792
rect 1398 2778 1402 2782
rect 1574 2778 1578 2782
rect 2110 2778 2114 2782
rect 2262 2778 2266 2782
rect 2270 2778 2274 2782
rect 2998 2778 3002 2782
rect 3070 2778 3074 2782
rect 3638 2778 3642 2782
rect 4030 2778 4034 2782
rect 4222 2778 4226 2782
rect 4598 2778 4602 2782
rect 1510 2768 1514 2772
rect 1582 2768 1586 2772
rect 2478 2768 2482 2772
rect 3718 2768 3722 2772
rect 3782 2768 3786 2772
rect 4238 2768 4242 2772
rect 4350 2768 4354 2772
rect 4582 2768 4586 2772
rect 4710 2768 4714 2772
rect 4870 2768 4874 2772
rect 5086 2768 5090 2772
rect 950 2758 954 2762
rect 966 2758 970 2762
rect 990 2758 994 2762
rect 1126 2758 1130 2762
rect 1158 2758 1162 2762
rect 2086 2758 2090 2762
rect 2870 2758 2874 2762
rect 2878 2758 2882 2762
rect 2966 2758 2970 2762
rect 3166 2758 3170 2762
rect 3758 2758 3762 2762
rect 3846 2758 3850 2762
rect 3862 2758 3866 2762
rect 4758 2758 4762 2762
rect 4894 2758 4898 2762
rect 254 2748 258 2752
rect 590 2748 594 2752
rect 614 2748 618 2752
rect 718 2748 722 2752
rect 734 2748 738 2752
rect 1502 2748 1506 2752
rect 1558 2748 1562 2752
rect 1662 2748 1666 2752
rect 1718 2748 1722 2752
rect 1958 2748 1962 2752
rect 2150 2748 2154 2752
rect 2246 2748 2250 2752
rect 2494 2748 2498 2752
rect 2790 2748 2794 2752
rect 2958 2748 2962 2752
rect 4086 2748 4090 2752
rect 4102 2748 4106 2752
rect 4110 2748 4114 2752
rect 4174 2748 4178 2752
rect 4390 2748 4394 2752
rect 4782 2748 4786 2752
rect 4910 2748 4914 2752
rect 4918 2748 4922 2752
rect 5166 2748 5170 2752
rect 310 2738 314 2742
rect 694 2738 698 2742
rect 734 2738 738 2742
rect 878 2738 882 2742
rect 1070 2738 1074 2742
rect 1102 2738 1106 2742
rect 1694 2738 1698 2742
rect 1758 2738 1762 2742
rect 1830 2738 1834 2742
rect 2246 2738 2250 2742
rect 2262 2738 2266 2742
rect 2446 2738 2450 2742
rect 2790 2738 2794 2742
rect 3102 2738 3106 2742
rect 3150 2738 3154 2742
rect 3166 2738 3170 2742
rect 3358 2738 3362 2742
rect 3574 2738 3578 2742
rect 3718 2738 3722 2742
rect 4662 2738 4666 2742
rect 4686 2738 4690 2742
rect 1110 2728 1114 2732
rect 1174 2728 1178 2732
rect 1454 2728 1458 2732
rect 1990 2728 1994 2732
rect 2254 2728 2258 2732
rect 2574 2728 2578 2732
rect 2614 2728 2618 2732
rect 2734 2728 2738 2732
rect 2974 2728 2978 2732
rect 3798 2728 3802 2732
rect 3886 2728 3890 2732
rect 4454 2728 4458 2732
rect 4950 2728 4954 2732
rect 5038 2728 5042 2732
rect 1118 2718 1122 2722
rect 1150 2718 1154 2722
rect 1158 2718 1162 2722
rect 1422 2718 1426 2722
rect 1486 2718 1490 2722
rect 1566 2718 1570 2722
rect 1590 2718 1594 2722
rect 1694 2718 1698 2722
rect 2070 2718 2074 2722
rect 2182 2718 2186 2722
rect 2590 2718 2594 2722
rect 2606 2718 2610 2722
rect 3742 2718 3746 2722
rect 3758 2718 3762 2722
rect 4334 2718 4338 2722
rect 4742 2718 4746 2722
rect 5062 2718 5066 2722
rect 246 2708 250 2712
rect 590 2708 594 2712
rect 1174 2708 1178 2712
rect 1422 2708 1426 2712
rect 1534 2708 1538 2712
rect 1598 2708 1602 2712
rect 2222 2708 2226 2712
rect 2518 2708 2522 2712
rect 2582 2708 2586 2712
rect 2878 2708 2882 2712
rect 3134 2708 3138 2712
rect 3974 2708 3978 2712
rect 4078 2708 4082 2712
rect 4302 2708 4306 2712
rect 4406 2708 4410 2712
rect 4470 2708 4474 2712
rect 4862 2708 4866 2712
rect 850 2703 854 2707
rect 858 2703 861 2707
rect 861 2703 862 2707
rect 1874 2703 1878 2707
rect 1882 2703 1885 2707
rect 1885 2703 1886 2707
rect 2890 2703 2894 2707
rect 2898 2703 2901 2707
rect 2901 2703 2902 2707
rect 3922 2703 3926 2707
rect 3930 2703 3933 2707
rect 3933 2703 3934 2707
rect 4938 2703 4942 2707
rect 4946 2703 4949 2707
rect 4949 2703 4950 2707
rect 2070 2698 2074 2702
rect 2614 2698 2618 2702
rect 2678 2698 2682 2702
rect 3030 2698 3034 2702
rect 3150 2698 3154 2702
rect 3246 2698 3250 2702
rect 3590 2698 3594 2702
rect 3854 2698 3858 2702
rect 4126 2698 4130 2702
rect 4142 2698 4146 2702
rect 4918 2698 4922 2702
rect 486 2688 490 2692
rect 630 2688 634 2692
rect 926 2688 930 2692
rect 1166 2688 1170 2692
rect 1654 2688 1658 2692
rect 1838 2688 1842 2692
rect 2606 2688 2610 2692
rect 3326 2688 3330 2692
rect 3494 2688 3498 2692
rect 3766 2688 3770 2692
rect 3886 2688 3890 2692
rect 4470 2688 4474 2692
rect 254 2678 258 2682
rect 1126 2678 1130 2682
rect 2046 2678 2050 2682
rect 2062 2678 2066 2682
rect 2182 2678 2186 2682
rect 2238 2678 2242 2682
rect 2286 2678 2290 2682
rect 2518 2678 2522 2682
rect 2990 2678 2994 2682
rect 3670 2678 3674 2682
rect 3798 2678 3802 2682
rect 3862 2678 3866 2682
rect 4190 2678 4194 2682
rect 4262 2678 4266 2682
rect 4582 2678 4586 2682
rect 5086 2678 5090 2682
rect 126 2668 130 2672
rect 518 2668 522 2672
rect 534 2668 538 2672
rect 710 2668 714 2672
rect 966 2668 970 2672
rect 1118 2668 1122 2672
rect 1334 2668 1338 2672
rect 2046 2668 2050 2672
rect 2150 2668 2154 2672
rect 2982 2668 2986 2672
rect 3606 2668 3610 2672
rect 3654 2668 3658 2672
rect 3726 2668 3730 2672
rect 4350 2668 4354 2672
rect 4358 2668 4362 2672
rect 4390 2668 4394 2672
rect 4830 2668 4834 2672
rect 86 2658 90 2662
rect 110 2658 114 2662
rect 582 2658 586 2662
rect 590 2658 594 2662
rect 758 2658 762 2662
rect 814 2658 818 2662
rect 830 2658 834 2662
rect 846 2658 850 2662
rect 1086 2658 1090 2662
rect 1102 2658 1106 2662
rect 1414 2658 1418 2662
rect 1814 2658 1818 2662
rect 2054 2658 2058 2662
rect 2102 2658 2106 2662
rect 2118 2658 2122 2662
rect 2166 2658 2170 2662
rect 2238 2658 2242 2662
rect 3534 2658 3538 2662
rect 3638 2658 3642 2662
rect 3662 2658 3666 2662
rect 3782 2658 3786 2662
rect 3790 2658 3794 2662
rect 4214 2658 4218 2662
rect 4366 2658 4370 2662
rect 4454 2658 4458 2662
rect 4502 2658 4506 2662
rect 4534 2658 4538 2662
rect 4774 2658 4778 2662
rect 4878 2658 4882 2662
rect 5014 2658 5018 2662
rect 550 2648 554 2652
rect 758 2648 762 2652
rect 1070 2648 1074 2652
rect 1710 2648 1714 2652
rect 2158 2648 2162 2652
rect 2198 2648 2202 2652
rect 2254 2648 2258 2652
rect 2798 2648 2802 2652
rect 3454 2648 3458 2652
rect 3470 2648 3474 2652
rect 4134 2648 4138 2652
rect 4318 2648 4322 2652
rect 4342 2648 4346 2652
rect 4414 2648 4418 2652
rect 4686 2648 4690 2652
rect 4814 2648 4818 2652
rect 5246 2648 5250 2652
rect 1790 2638 1794 2642
rect 1998 2638 2002 2642
rect 3038 2638 3042 2642
rect 3534 2638 3538 2642
rect 3606 2638 3610 2642
rect 3750 2638 3754 2642
rect 4302 2638 4306 2642
rect 694 2628 698 2632
rect 1110 2628 1114 2632
rect 1782 2628 1786 2632
rect 1790 2628 1794 2632
rect 2094 2628 2098 2632
rect 2150 2628 2154 2632
rect 2310 2628 2314 2632
rect 2566 2628 2570 2632
rect 2598 2628 2602 2632
rect 3222 2628 3226 2632
rect 3830 2628 3834 2632
rect 4022 2628 4026 2632
rect 614 2618 618 2622
rect 1902 2618 1906 2622
rect 1966 2618 1970 2622
rect 2214 2618 2218 2622
rect 2622 2618 2626 2622
rect 2766 2618 2770 2622
rect 2886 2618 2890 2622
rect 2950 2618 2954 2622
rect 3366 2618 3370 2622
rect 3422 2618 3426 2622
rect 3734 2618 3738 2622
rect 4358 2618 4362 2622
rect 4374 2618 4378 2622
rect 1070 2608 1074 2612
rect 1774 2608 1778 2612
rect 2174 2608 2178 2612
rect 2222 2608 2226 2612
rect 2574 2608 2578 2612
rect 2582 2608 2586 2612
rect 2822 2608 2826 2612
rect 3494 2608 3498 2612
rect 3782 2608 3786 2612
rect 3814 2608 3818 2612
rect 4470 2608 4474 2612
rect 4526 2608 4530 2612
rect 330 2603 334 2607
rect 338 2603 341 2607
rect 341 2603 342 2607
rect 1354 2603 1358 2607
rect 1362 2603 1365 2607
rect 1365 2603 1366 2607
rect 2386 2603 2390 2607
rect 2394 2603 2397 2607
rect 2397 2603 2398 2607
rect 3402 2603 3406 2607
rect 3410 2603 3413 2607
rect 3413 2603 3414 2607
rect 4426 2603 4430 2607
rect 4434 2603 4437 2607
rect 4437 2603 4438 2607
rect 846 2598 850 2602
rect 1398 2598 1402 2602
rect 1622 2598 1626 2602
rect 1686 2598 1690 2602
rect 2078 2598 2082 2602
rect 2174 2598 2178 2602
rect 2782 2598 2786 2602
rect 3054 2598 3058 2602
rect 3062 2598 3066 2602
rect 3390 2598 3394 2602
rect 3558 2598 3562 2602
rect 3718 2598 3722 2602
rect 3750 2598 3754 2602
rect 4502 2598 4506 2602
rect 4838 2598 4842 2602
rect 4990 2598 4994 2602
rect 262 2588 266 2592
rect 294 2588 298 2592
rect 2598 2588 2602 2592
rect 3214 2588 3218 2592
rect 3222 2588 3226 2592
rect 3686 2588 3690 2592
rect 3710 2588 3714 2592
rect 4038 2588 4042 2592
rect 4382 2588 4386 2592
rect 4398 2588 4402 2592
rect 4798 2588 4802 2592
rect 5086 2588 5090 2592
rect 718 2578 722 2582
rect 1094 2578 1098 2582
rect 1982 2578 1986 2582
rect 4614 2578 4618 2582
rect 734 2568 738 2572
rect 838 2568 842 2572
rect 870 2568 874 2572
rect 926 2568 930 2572
rect 1142 2568 1146 2572
rect 1222 2568 1226 2572
rect 1526 2568 1530 2572
rect 1702 2568 1706 2572
rect 2094 2568 2098 2572
rect 2134 2568 2138 2572
rect 2438 2568 2442 2572
rect 2926 2568 2930 2572
rect 3478 2568 3482 2572
rect 3550 2568 3554 2572
rect 3774 2568 3778 2572
rect 4614 2568 4618 2572
rect 5166 2568 5170 2572
rect 374 2558 378 2562
rect 470 2558 474 2562
rect 1142 2558 1146 2562
rect 1526 2558 1530 2562
rect 1566 2558 1570 2562
rect 1758 2558 1762 2562
rect 1918 2558 1922 2562
rect 2078 2558 2082 2562
rect 2182 2558 2186 2562
rect 2206 2558 2210 2562
rect 2238 2558 2242 2562
rect 2254 2558 2258 2562
rect 2406 2558 2410 2562
rect 2422 2558 2426 2562
rect 2558 2558 2562 2562
rect 2766 2558 2770 2562
rect 2894 2558 2898 2562
rect 3070 2558 3074 2562
rect 3254 2558 3258 2562
rect 3414 2558 3418 2562
rect 4134 2558 4138 2562
rect 4486 2558 4490 2562
rect 4590 2558 4594 2562
rect 5118 2558 5122 2562
rect 5190 2558 5194 2562
rect 110 2548 114 2552
rect 270 2548 274 2552
rect 654 2548 658 2552
rect 662 2548 666 2552
rect 1326 2548 1330 2552
rect 1422 2548 1426 2552
rect 1726 2548 1730 2552
rect 2782 2548 2786 2552
rect 2790 2548 2794 2552
rect 2950 2548 2954 2552
rect 2982 2548 2986 2552
rect 3014 2548 3018 2552
rect 3022 2548 3026 2552
rect 3086 2548 3090 2552
rect 3246 2548 3250 2552
rect 3790 2548 3794 2552
rect 3822 2548 3826 2552
rect 3910 2548 3914 2552
rect 4054 2548 4058 2552
rect 4118 2548 4122 2552
rect 4454 2548 4458 2552
rect 4878 2548 4882 2552
rect 5246 2548 5250 2552
rect 254 2538 258 2542
rect 1054 2538 1058 2542
rect 2422 2538 2426 2542
rect 2718 2538 2722 2542
rect 2990 2538 2994 2542
rect 3030 2538 3034 2542
rect 3078 2538 3082 2542
rect 3102 2538 3106 2542
rect 3126 2538 3130 2542
rect 3166 2538 3170 2542
rect 3550 2538 3554 2542
rect 3774 2538 3778 2542
rect 4422 2538 4426 2542
rect 4606 2538 4610 2542
rect 5238 2538 5242 2542
rect 1334 2528 1338 2532
rect 1446 2528 1450 2532
rect 1630 2528 1634 2532
rect 1942 2528 1946 2532
rect 2102 2528 2106 2532
rect 2262 2528 2266 2532
rect 2382 2528 2386 2532
rect 2750 2528 2754 2532
rect 3094 2528 3098 2532
rect 3134 2528 3138 2532
rect 3486 2528 3490 2532
rect 3502 2528 3506 2532
rect 3590 2528 3594 2532
rect 3982 2528 3986 2532
rect 4278 2528 4282 2532
rect 4342 2528 4346 2532
rect 4462 2528 4466 2532
rect 1454 2518 1458 2522
rect 1462 2518 1466 2522
rect 2134 2518 2138 2522
rect 2230 2518 2234 2522
rect 2654 2518 2658 2522
rect 2670 2518 2674 2522
rect 2878 2518 2882 2522
rect 2934 2518 2938 2522
rect 3166 2518 3170 2522
rect 3294 2518 3298 2522
rect 3470 2518 3474 2522
rect 4030 2518 4034 2522
rect 4038 2518 4042 2522
rect 4310 2518 4314 2522
rect 5086 2518 5090 2522
rect 5254 2518 5258 2522
rect 686 2508 690 2512
rect 2342 2508 2346 2512
rect 2350 2508 2354 2512
rect 2726 2508 2730 2512
rect 2806 2508 2810 2512
rect 2942 2508 2946 2512
rect 2950 2508 2954 2512
rect 3270 2508 3274 2512
rect 3366 2508 3370 2512
rect 3782 2508 3786 2512
rect 3910 2508 3914 2512
rect 850 2503 854 2507
rect 858 2503 861 2507
rect 861 2503 862 2507
rect 1874 2503 1878 2507
rect 1882 2503 1885 2507
rect 1885 2503 1886 2507
rect 1502 2498 1506 2502
rect 1518 2498 1522 2502
rect 2078 2498 2082 2502
rect 2158 2498 2162 2502
rect 2174 2498 2178 2502
rect 2890 2503 2894 2507
rect 2898 2503 2901 2507
rect 2901 2503 2902 2507
rect 3922 2503 3926 2507
rect 3930 2503 3933 2507
rect 3933 2503 3934 2507
rect 2630 2498 2634 2502
rect 3046 2498 3050 2502
rect 3222 2498 3226 2502
rect 3302 2498 3306 2502
rect 3342 2498 3346 2502
rect 3350 2498 3354 2502
rect 3646 2498 3650 2502
rect 4078 2498 4082 2502
rect 4230 2498 4234 2502
rect 5190 2508 5194 2512
rect 4938 2503 4942 2507
rect 4946 2503 4949 2507
rect 4949 2503 4950 2507
rect 822 2488 826 2492
rect 1990 2488 1994 2492
rect 2022 2488 2026 2492
rect 2054 2488 2058 2492
rect 2094 2488 2098 2492
rect 2374 2488 2378 2492
rect 2782 2488 2786 2492
rect 2798 2488 2802 2492
rect 2942 2488 2946 2492
rect 3022 2488 3026 2492
rect 3286 2488 3290 2492
rect 4758 2488 4762 2492
rect 5190 2488 5194 2492
rect 1902 2478 1906 2482
rect 1918 2478 1922 2482
rect 2086 2478 2090 2482
rect 2102 2478 2106 2482
rect 2382 2478 2386 2482
rect 2558 2478 2562 2482
rect 2662 2478 2666 2482
rect 3078 2478 3082 2482
rect 3230 2478 3234 2482
rect 3614 2478 3618 2482
rect 3630 2478 3634 2482
rect 862 2468 866 2472
rect 1022 2468 1026 2472
rect 1494 2468 1498 2472
rect 1622 2468 1626 2472
rect 1830 2468 1834 2472
rect 1886 2468 1890 2472
rect 2022 2468 2026 2472
rect 2358 2468 2362 2472
rect 278 2458 282 2462
rect 614 2458 618 2462
rect 702 2458 706 2462
rect 878 2458 882 2462
rect 974 2458 978 2462
rect 1198 2458 1202 2462
rect 1526 2458 1530 2462
rect 1542 2458 1546 2462
rect 1582 2458 1586 2462
rect 2718 2468 2722 2472
rect 2750 2468 2754 2472
rect 3206 2468 3210 2472
rect 3286 2468 3290 2472
rect 3334 2468 3338 2472
rect 4142 2478 4146 2482
rect 4190 2478 4194 2482
rect 4326 2478 4330 2482
rect 3518 2468 3522 2472
rect 3726 2468 3730 2472
rect 3838 2468 3842 2472
rect 3878 2468 3882 2472
rect 4110 2468 4114 2472
rect 4198 2468 4202 2472
rect 4214 2468 4218 2472
rect 4270 2468 4274 2472
rect 4294 2468 4298 2472
rect 4350 2468 4354 2472
rect 4390 2468 4394 2472
rect 4414 2468 4418 2472
rect 4430 2468 4434 2472
rect 4518 2468 4522 2472
rect 1798 2458 1802 2462
rect 1838 2458 1842 2462
rect 1894 2458 1898 2462
rect 1934 2458 1938 2462
rect 2078 2458 2082 2462
rect 2110 2458 2114 2462
rect 2126 2458 2130 2462
rect 2286 2458 2290 2462
rect 2334 2458 2338 2462
rect 2446 2458 2450 2462
rect 2462 2458 2466 2462
rect 2510 2458 2514 2462
rect 2542 2458 2546 2462
rect 2694 2458 2698 2462
rect 2710 2458 2714 2462
rect 2726 2458 2730 2462
rect 2846 2458 2850 2462
rect 2966 2458 2970 2462
rect 3014 2458 3018 2462
rect 3166 2458 3170 2462
rect 3182 2458 3186 2462
rect 3326 2458 3330 2462
rect 3542 2458 3546 2462
rect 3574 2458 3578 2462
rect 3886 2458 3890 2462
rect 4094 2458 4098 2462
rect 4254 2458 4258 2462
rect 4638 2458 4642 2462
rect 646 2448 650 2452
rect 894 2448 898 2452
rect 1454 2448 1458 2452
rect 1646 2448 1650 2452
rect 1822 2448 1826 2452
rect 1926 2448 1930 2452
rect 1966 2448 1970 2452
rect 2086 2448 2090 2452
rect 2142 2448 2146 2452
rect 2454 2448 2458 2452
rect 2838 2448 2842 2452
rect 2934 2448 2938 2452
rect 3246 2448 3250 2452
rect 3310 2448 3314 2452
rect 3734 2448 3738 2452
rect 4046 2448 4050 2452
rect 4286 2448 4290 2452
rect 4414 2448 4418 2452
rect 4542 2448 4546 2452
rect 4734 2448 4738 2452
rect 4742 2448 4746 2452
rect 4782 2448 4786 2452
rect 4798 2448 4802 2452
rect 5022 2448 5026 2452
rect 142 2438 146 2442
rect 1014 2438 1018 2442
rect 1158 2438 1162 2442
rect 1302 2438 1306 2442
rect 2086 2438 2090 2442
rect 2534 2438 2538 2442
rect 3366 2438 3370 2442
rect 3966 2438 3970 2442
rect 4270 2438 4274 2442
rect 4558 2438 4562 2442
rect 4638 2438 4642 2442
rect 4790 2438 4794 2442
rect 4966 2438 4970 2442
rect 710 2428 714 2432
rect 902 2428 906 2432
rect 934 2428 938 2432
rect 1230 2428 1234 2432
rect 1342 2428 1346 2432
rect 2358 2428 2362 2432
rect 2814 2428 2818 2432
rect 2902 2428 2906 2432
rect 2958 2428 2962 2432
rect 3062 2428 3066 2432
rect 3190 2428 3194 2432
rect 3646 2428 3650 2432
rect 4246 2428 4250 2432
rect 4294 2428 4298 2432
rect 4710 2428 4714 2432
rect 1558 2418 1562 2422
rect 1750 2418 1754 2422
rect 1942 2418 1946 2422
rect 2158 2418 2162 2422
rect 3222 2418 3226 2422
rect 3734 2418 3738 2422
rect 4070 2418 4074 2422
rect 5294 2418 5298 2422
rect 1046 2408 1050 2412
rect 1062 2408 1066 2412
rect 1406 2408 1410 2412
rect 1470 2408 1474 2412
rect 1550 2408 1554 2412
rect 2086 2408 2090 2412
rect 2094 2408 2098 2412
rect 2326 2408 2330 2412
rect 2446 2408 2450 2412
rect 2558 2408 2562 2412
rect 2790 2408 2794 2412
rect 2862 2408 2866 2412
rect 2950 2408 2954 2412
rect 3574 2408 3578 2412
rect 3894 2408 3898 2412
rect 3902 2408 3906 2412
rect 4542 2408 4546 2412
rect 5286 2408 5290 2412
rect 330 2403 334 2407
rect 338 2403 341 2407
rect 341 2403 342 2407
rect 1354 2403 1358 2407
rect 1362 2403 1365 2407
rect 1365 2403 1366 2407
rect 2386 2403 2390 2407
rect 2394 2403 2397 2407
rect 2397 2403 2398 2407
rect 278 2398 282 2402
rect 574 2398 578 2402
rect 1382 2398 1386 2402
rect 1398 2398 1402 2402
rect 1774 2398 1778 2402
rect 2118 2398 2122 2402
rect 3402 2403 3406 2407
rect 3410 2403 3413 2407
rect 3413 2403 3414 2407
rect 4426 2403 4430 2407
rect 4434 2403 4437 2407
rect 4437 2403 4438 2407
rect 2686 2398 2690 2402
rect 2718 2398 2722 2402
rect 3094 2398 3098 2402
rect 3142 2398 3146 2402
rect 3734 2398 3738 2402
rect 4406 2398 4410 2402
rect 4686 2398 4690 2402
rect 1230 2388 1234 2392
rect 1382 2388 1386 2392
rect 1638 2388 1642 2392
rect 2478 2388 2482 2392
rect 2574 2388 2578 2392
rect 3342 2388 3346 2392
rect 3822 2388 3826 2392
rect 4158 2388 4162 2392
rect 2158 2378 2162 2382
rect 2310 2378 2314 2382
rect 4614 2388 4618 2392
rect 5030 2388 5034 2392
rect 5102 2388 5106 2392
rect 3166 2378 3170 2382
rect 3310 2378 3314 2382
rect 3982 2378 3986 2382
rect 4710 2378 4714 2382
rect 4894 2378 4898 2382
rect 5158 2378 5162 2382
rect 526 2368 530 2372
rect 1846 2368 1850 2372
rect 1878 2368 1882 2372
rect 1926 2368 1930 2372
rect 2230 2368 2234 2372
rect 2270 2368 2274 2372
rect 2278 2368 2282 2372
rect 2494 2368 2498 2372
rect 2502 2368 2506 2372
rect 2974 2368 2978 2372
rect 3030 2368 3034 2372
rect 3486 2368 3490 2372
rect 3502 2368 3506 2372
rect 3598 2368 3602 2372
rect 4238 2368 4242 2372
rect 5054 2368 5058 2372
rect 5286 2368 5290 2372
rect 662 2358 666 2362
rect 1310 2358 1314 2362
rect 1542 2358 1546 2362
rect 1774 2358 1778 2362
rect 1806 2358 1810 2362
rect 2094 2358 2098 2362
rect 2206 2358 2210 2362
rect 2270 2358 2274 2362
rect 2518 2358 2522 2362
rect 2622 2358 2626 2362
rect 2646 2358 2650 2362
rect 3014 2358 3018 2362
rect 3118 2358 3122 2362
rect 3318 2358 3322 2362
rect 3614 2358 3618 2362
rect 3894 2358 3898 2362
rect 4070 2358 4074 2362
rect 4102 2358 4106 2362
rect 4630 2358 4634 2362
rect 4790 2358 4794 2362
rect 494 2348 498 2352
rect 526 2348 530 2352
rect 614 2348 618 2352
rect 654 2348 658 2352
rect 702 2348 706 2352
rect 742 2348 746 2352
rect 926 2348 930 2352
rect 1366 2348 1370 2352
rect 1430 2348 1434 2352
rect 1462 2348 1466 2352
rect 1526 2348 1530 2352
rect 1670 2348 1674 2352
rect 1742 2348 1746 2352
rect 1838 2348 1842 2352
rect 1926 2348 1930 2352
rect 2070 2348 2074 2352
rect 2134 2348 2138 2352
rect 2406 2348 2410 2352
rect 2430 2348 2434 2352
rect 2542 2348 2546 2352
rect 2822 2348 2826 2352
rect 2862 2348 2866 2352
rect 3046 2348 3050 2352
rect 3062 2348 3066 2352
rect 3094 2348 3098 2352
rect 3190 2348 3194 2352
rect 3326 2348 3330 2352
rect 3438 2348 3442 2352
rect 3646 2348 3650 2352
rect 3678 2348 3682 2352
rect 3982 2348 3986 2352
rect 4310 2348 4314 2352
rect 4350 2348 4354 2352
rect 4614 2348 4618 2352
rect 4958 2348 4962 2352
rect 4966 2348 4970 2352
rect 5158 2348 5162 2352
rect 5294 2348 5298 2352
rect 462 2338 466 2342
rect 518 2338 522 2342
rect 1126 2338 1130 2342
rect 1502 2338 1506 2342
rect 1630 2338 1634 2342
rect 1694 2338 1698 2342
rect 1750 2338 1754 2342
rect 2246 2338 2250 2342
rect 2510 2338 2514 2342
rect 2766 2338 2770 2342
rect 2846 2338 2850 2342
rect 2894 2338 2898 2342
rect 2958 2338 2962 2342
rect 2990 2338 2994 2342
rect 3006 2338 3010 2342
rect 3022 2338 3026 2342
rect 3334 2338 3338 2342
rect 4102 2338 4106 2342
rect 4806 2338 4810 2342
rect 5174 2338 5178 2342
rect 5246 2338 5250 2342
rect 814 2328 818 2332
rect 934 2328 938 2332
rect 1614 2328 1618 2332
rect 2038 2328 2042 2332
rect 2110 2328 2114 2332
rect 2318 2328 2322 2332
rect 2670 2328 2674 2332
rect 2806 2328 2810 2332
rect 3134 2328 3138 2332
rect 3214 2328 3218 2332
rect 3390 2328 3394 2332
rect 3758 2328 3762 2332
rect 3886 2328 3890 2332
rect 4318 2328 4322 2332
rect 838 2318 842 2322
rect 1518 2318 1522 2322
rect 1558 2318 1562 2322
rect 1606 2318 1610 2322
rect 1686 2318 1690 2322
rect 1758 2318 1762 2322
rect 2062 2318 2066 2322
rect 2190 2318 2194 2322
rect 2526 2318 2530 2322
rect 3142 2318 3146 2322
rect 3342 2318 3346 2322
rect 3374 2318 3378 2322
rect 3414 2318 3418 2322
rect 3486 2318 3490 2322
rect 3614 2318 3618 2322
rect 3846 2318 3850 2322
rect 4022 2318 4026 2322
rect 4286 2318 4290 2322
rect 4302 2318 4306 2322
rect 742 2308 746 2312
rect 974 2308 978 2312
rect 1862 2308 1866 2312
rect 1974 2308 1978 2312
rect 1990 2308 1994 2312
rect 2038 2308 2042 2312
rect 2198 2308 2202 2312
rect 2318 2308 2322 2312
rect 2918 2308 2922 2312
rect 3190 2308 3194 2312
rect 3406 2308 3410 2312
rect 3518 2308 3522 2312
rect 3582 2308 3586 2312
rect 3790 2308 3794 2312
rect 3910 2308 3914 2312
rect 3990 2308 3994 2312
rect 3998 2308 4002 2312
rect 5126 2308 5130 2312
rect 5270 2308 5274 2312
rect 850 2303 854 2307
rect 858 2303 861 2307
rect 861 2303 862 2307
rect 1874 2303 1878 2307
rect 1882 2303 1885 2307
rect 1885 2303 1886 2307
rect 2890 2303 2894 2307
rect 2898 2303 2901 2307
rect 2901 2303 2902 2307
rect 3922 2303 3926 2307
rect 3930 2303 3933 2307
rect 3933 2303 3934 2307
rect 4938 2303 4942 2307
rect 4946 2303 4949 2307
rect 4949 2303 4950 2307
rect 1022 2298 1026 2302
rect 1438 2298 1442 2302
rect 1990 2298 1994 2302
rect 2278 2298 2282 2302
rect 2718 2298 2722 2302
rect 2806 2298 2810 2302
rect 2950 2298 2954 2302
rect 3222 2298 3226 2302
rect 3230 2298 3234 2302
rect 3982 2298 3986 2302
rect 5014 2298 5018 2302
rect 654 2288 658 2292
rect 974 2288 978 2292
rect 1958 2288 1962 2292
rect 2006 2288 2010 2292
rect 2054 2288 2058 2292
rect 2510 2288 2514 2292
rect 2574 2288 2578 2292
rect 2662 2288 2666 2292
rect 2670 2288 2674 2292
rect 2710 2288 2714 2292
rect 2942 2288 2946 2292
rect 3470 2288 3474 2292
rect 3558 2288 3562 2292
rect 3694 2288 3698 2292
rect 4334 2288 4338 2292
rect 4438 2288 4442 2292
rect 5254 2288 5258 2292
rect 366 2278 370 2282
rect 798 2278 802 2282
rect 1270 2278 1274 2282
rect 1374 2278 1378 2282
rect 1390 2278 1394 2282
rect 1414 2278 1418 2282
rect 2062 2278 2066 2282
rect 2270 2278 2274 2282
rect 2790 2278 2794 2282
rect 3526 2278 3530 2282
rect 3590 2278 3594 2282
rect 3678 2278 3682 2282
rect 3998 2278 4002 2282
rect 4230 2278 4234 2282
rect 4558 2278 4562 2282
rect 286 2268 290 2272
rect 1006 2268 1010 2272
rect 1206 2268 1210 2272
rect 1286 2268 1290 2272
rect 1550 2268 1554 2272
rect 1998 2268 2002 2272
rect 2046 2268 2050 2272
rect 2070 2268 2074 2272
rect 2158 2268 2162 2272
rect 2254 2268 2258 2272
rect 2302 2268 2306 2272
rect 2478 2268 2482 2272
rect 2574 2268 2578 2272
rect 2646 2268 2650 2272
rect 2846 2268 2850 2272
rect 3014 2268 3018 2272
rect 3126 2268 3130 2272
rect 3134 2268 3138 2272
rect 3206 2268 3210 2272
rect 3262 2268 3266 2272
rect 3318 2268 3322 2272
rect 3366 2268 3370 2272
rect 214 2258 218 2262
rect 278 2258 282 2262
rect 526 2258 530 2262
rect 718 2258 722 2262
rect 766 2258 770 2262
rect 974 2258 978 2262
rect 990 2258 994 2262
rect 1486 2258 1490 2262
rect 1894 2258 1898 2262
rect 1942 2258 1946 2262
rect 3438 2268 3442 2272
rect 3470 2268 3474 2272
rect 3486 2268 3490 2272
rect 3502 2268 3506 2272
rect 3526 2268 3530 2272
rect 3574 2268 3578 2272
rect 3630 2268 3634 2272
rect 3726 2268 3730 2272
rect 3830 2268 3834 2272
rect 4134 2268 4138 2272
rect 4462 2268 4466 2272
rect 4742 2268 4746 2272
rect 4766 2268 4770 2272
rect 5150 2268 5154 2272
rect 5302 2268 5306 2272
rect 2198 2258 2202 2262
rect 2446 2258 2450 2262
rect 2462 2258 2466 2262
rect 2566 2258 2570 2262
rect 2574 2258 2578 2262
rect 2662 2258 2666 2262
rect 2726 2258 2730 2262
rect 326 2248 330 2252
rect 1302 2248 1306 2252
rect 1342 2248 1346 2252
rect 1422 2248 1426 2252
rect 2142 2248 2146 2252
rect 2814 2258 2818 2262
rect 2998 2258 3002 2262
rect 3662 2258 3666 2262
rect 3774 2258 3778 2262
rect 3814 2258 3818 2262
rect 4030 2258 4034 2262
rect 4038 2258 4042 2262
rect 4190 2258 4194 2262
rect 4462 2258 4466 2262
rect 4534 2258 4538 2262
rect 4582 2258 4586 2262
rect 4806 2258 4810 2262
rect 2342 2248 2346 2252
rect 2350 2248 2354 2252
rect 2422 2248 2426 2252
rect 2558 2248 2562 2252
rect 2686 2248 2690 2252
rect 2718 2248 2722 2252
rect 2782 2248 2786 2252
rect 2910 2248 2914 2252
rect 3374 2248 3378 2252
rect 3390 2248 3394 2252
rect 3550 2248 3554 2252
rect 3566 2248 3570 2252
rect 4614 2248 4618 2252
rect 5078 2248 5082 2252
rect 5302 2248 5306 2252
rect 2366 2238 2370 2242
rect 2422 2238 2426 2242
rect 2454 2238 2458 2242
rect 2534 2238 2538 2242
rect 3358 2238 3362 2242
rect 4054 2238 4058 2242
rect 4878 2238 4882 2242
rect 5086 2238 5090 2242
rect 246 2228 250 2232
rect 966 2228 970 2232
rect 2318 2228 2322 2232
rect 2358 2228 2362 2232
rect 2638 2228 2642 2232
rect 2694 2228 2698 2232
rect 2750 2228 2754 2232
rect 2774 2228 2778 2232
rect 4358 2228 4362 2232
rect 4438 2228 4442 2232
rect 4758 2228 4762 2232
rect 4926 2228 4930 2232
rect 1486 2218 1490 2222
rect 1494 2218 1498 2222
rect 1750 2218 1754 2222
rect 2022 2218 2026 2222
rect 2374 2218 2378 2222
rect 2878 2218 2882 2222
rect 3262 2218 3266 2222
rect 3462 2218 3466 2222
rect 3486 2218 3490 2222
rect 4086 2218 4090 2222
rect 4710 2218 4714 2222
rect 4966 2218 4970 2222
rect 5198 2218 5202 2222
rect 5246 2218 5250 2222
rect 1334 2208 1338 2212
rect 1646 2208 1650 2212
rect 1726 2208 1730 2212
rect 2286 2208 2290 2212
rect 2358 2208 2362 2212
rect 2406 2208 2410 2212
rect 2950 2208 2954 2212
rect 3206 2208 3210 2212
rect 3470 2208 3474 2212
rect 4262 2208 4266 2212
rect 4446 2208 4450 2212
rect 4886 2208 4890 2212
rect 5262 2208 5266 2212
rect 330 2203 334 2207
rect 338 2203 341 2207
rect 341 2203 342 2207
rect 1354 2203 1358 2207
rect 1362 2203 1365 2207
rect 1365 2203 1366 2207
rect 2386 2203 2390 2207
rect 2394 2203 2397 2207
rect 2397 2203 2398 2207
rect 3402 2203 3406 2207
rect 3410 2203 3413 2207
rect 3413 2203 3414 2207
rect 4426 2203 4430 2207
rect 4434 2203 4437 2207
rect 4437 2203 4438 2207
rect 750 2198 754 2202
rect 1278 2198 1282 2202
rect 1830 2198 1834 2202
rect 2086 2198 2090 2202
rect 2206 2198 2210 2202
rect 2374 2198 2378 2202
rect 2534 2198 2538 2202
rect 2998 2198 3002 2202
rect 3886 2198 3890 2202
rect 3966 2198 3970 2202
rect 5278 2198 5282 2202
rect 734 2188 738 2192
rect 806 2188 810 2192
rect 942 2188 946 2192
rect 1654 2188 1658 2192
rect 1742 2188 1746 2192
rect 1942 2188 1946 2192
rect 2534 2188 2538 2192
rect 2822 2188 2826 2192
rect 3838 2188 3842 2192
rect 3894 2188 3898 2192
rect 4390 2188 4394 2192
rect 5182 2188 5186 2192
rect 1222 2178 1226 2182
rect 1566 2178 1570 2182
rect 1590 2178 1594 2182
rect 2270 2178 2274 2182
rect 2326 2178 2330 2182
rect 2798 2178 2802 2182
rect 3174 2178 3178 2182
rect 3254 2178 3258 2182
rect 3438 2178 3442 2182
rect 3710 2178 3714 2182
rect 686 2168 690 2172
rect 1246 2168 1250 2172
rect 1686 2168 1690 2172
rect 1718 2168 1722 2172
rect 1742 2168 1746 2172
rect 2182 2168 2186 2172
rect 2302 2168 2306 2172
rect 2334 2168 2338 2172
rect 2550 2168 2554 2172
rect 2614 2168 2618 2172
rect 3718 2168 3722 2172
rect 3822 2168 3826 2172
rect 5014 2168 5018 2172
rect 5030 2168 5034 2172
rect 5094 2168 5098 2172
rect 5286 2168 5290 2172
rect 302 2158 306 2162
rect 718 2158 722 2162
rect 742 2158 746 2162
rect 1254 2158 1258 2162
rect 1670 2158 1674 2162
rect 1966 2158 1970 2162
rect 2030 2158 2034 2162
rect 2206 2158 2210 2162
rect 2246 2158 2250 2162
rect 2478 2158 2482 2162
rect 3246 2158 3250 2162
rect 3262 2158 3266 2162
rect 4094 2158 4098 2162
rect 4894 2158 4898 2162
rect 4990 2158 4994 2162
rect 5094 2158 5098 2162
rect 1750 2148 1754 2152
rect 1870 2148 1874 2152
rect 2094 2148 2098 2152
rect 2302 2148 2306 2152
rect 2870 2148 2874 2152
rect 2918 2148 2922 2152
rect 3302 2148 3306 2152
rect 3310 2148 3314 2152
rect 3358 2148 3362 2152
rect 3734 2148 3738 2152
rect 3838 2148 3842 2152
rect 3942 2148 3946 2152
rect 4286 2148 4290 2152
rect 4302 2148 4306 2152
rect 4374 2148 4378 2152
rect 4446 2148 4450 2152
rect 4782 2148 4786 2152
rect 4814 2148 4818 2152
rect 4918 2148 4922 2152
rect 5022 2148 5026 2152
rect 5182 2148 5186 2152
rect 566 2138 570 2142
rect 662 2138 666 2142
rect 1214 2138 1218 2142
rect 1238 2138 1242 2142
rect 1542 2138 1546 2142
rect 1638 2138 1642 2142
rect 1670 2138 1674 2142
rect 1934 2138 1938 2142
rect 2054 2138 2058 2142
rect 2270 2138 2274 2142
rect 2286 2138 2290 2142
rect 2342 2138 2346 2142
rect 2494 2138 2498 2142
rect 2542 2138 2546 2142
rect 3222 2138 3226 2142
rect 3286 2138 3290 2142
rect 3302 2138 3306 2142
rect 3830 2138 3834 2142
rect 3878 2138 3882 2142
rect 4190 2138 4194 2142
rect 4406 2138 4410 2142
rect 5142 2138 5146 2142
rect 110 2128 114 2132
rect 286 2128 290 2132
rect 734 2128 738 2132
rect 1430 2128 1434 2132
rect 1518 2128 1522 2132
rect 1606 2128 1610 2132
rect 1694 2128 1698 2132
rect 1758 2128 1762 2132
rect 2334 2128 2338 2132
rect 2366 2128 2370 2132
rect 3334 2128 3338 2132
rect 3590 2128 3594 2132
rect 4254 2128 4258 2132
rect 4454 2128 4458 2132
rect 4766 2128 4770 2132
rect 5046 2128 5050 2132
rect 5182 2128 5186 2132
rect 670 2118 674 2122
rect 750 2118 754 2122
rect 766 2118 770 2122
rect 1030 2118 1034 2122
rect 1526 2118 1530 2122
rect 2750 2118 2754 2122
rect 2942 2118 2946 2122
rect 3062 2118 3066 2122
rect 3070 2118 3074 2122
rect 3166 2118 3170 2122
rect 3198 2118 3202 2122
rect 3254 2118 3258 2122
rect 446 2108 450 2112
rect 838 2108 842 2112
rect 1494 2108 1498 2112
rect 1894 2108 1898 2112
rect 2214 2108 2218 2112
rect 2294 2108 2298 2112
rect 2318 2108 2322 2112
rect 3670 2108 3674 2112
rect 3694 2108 3698 2112
rect 3942 2108 3946 2112
rect 4382 2108 4386 2112
rect 5110 2108 5114 2112
rect 5222 2108 5226 2112
rect 850 2103 854 2107
rect 858 2103 861 2107
rect 861 2103 862 2107
rect 1874 2103 1878 2107
rect 1882 2103 1885 2107
rect 1885 2103 1886 2107
rect 2890 2103 2894 2107
rect 2898 2103 2901 2107
rect 2901 2103 2902 2107
rect 302 2098 306 2102
rect 1638 2098 1642 2102
rect 2406 2098 2410 2102
rect 2430 2098 2434 2102
rect 2582 2098 2586 2102
rect 2758 2098 2762 2102
rect 2830 2098 2834 2102
rect 3006 2098 3010 2102
rect 3922 2103 3926 2107
rect 3930 2103 3933 2107
rect 3933 2103 3934 2107
rect 4938 2103 4942 2107
rect 4946 2103 4949 2107
rect 4949 2103 4950 2107
rect 3462 2098 3466 2102
rect 3758 2098 3762 2102
rect 3806 2098 3810 2102
rect 4094 2098 4098 2102
rect 4246 2098 4250 2102
rect 4454 2098 4458 2102
rect 4494 2098 4498 2102
rect 5102 2098 5106 2102
rect 542 2088 546 2092
rect 1022 2088 1026 2092
rect 1526 2088 1530 2092
rect 2958 2088 2962 2092
rect 3142 2088 3146 2092
rect 3150 2088 3154 2092
rect 3422 2088 3426 2092
rect 3894 2088 3898 2092
rect 4366 2088 4370 2092
rect 1006 2078 1010 2082
rect 1014 2078 1018 2082
rect 1198 2078 1202 2082
rect 1214 2078 1218 2082
rect 1566 2078 1570 2082
rect 1582 2078 1586 2082
rect 1758 2078 1762 2082
rect 1934 2078 1938 2082
rect 2230 2078 2234 2082
rect 2270 2078 2274 2082
rect 2470 2078 2474 2082
rect 2694 2078 2698 2082
rect 3174 2078 3178 2082
rect 3430 2078 3434 2082
rect 3614 2078 3618 2082
rect 3686 2078 3690 2082
rect 3766 2078 3770 2082
rect 3774 2078 3778 2082
rect 4062 2078 4066 2082
rect 4414 2078 4418 2082
rect 4478 2078 4482 2082
rect 4510 2078 4514 2082
rect 1174 2068 1178 2072
rect 1318 2068 1322 2072
rect 1558 2068 1562 2072
rect 1886 2068 1890 2072
rect 1918 2068 1922 2072
rect 1998 2068 2002 2072
rect 2158 2068 2162 2072
rect 2366 2068 2370 2072
rect 2502 2068 2506 2072
rect 2638 2068 2642 2072
rect 2750 2068 2754 2072
rect 3374 2068 3378 2072
rect 3406 2068 3410 2072
rect 3534 2068 3538 2072
rect 4038 2068 4042 2072
rect 4142 2068 4146 2072
rect 4174 2068 4178 2072
rect 4222 2068 4226 2072
rect 4342 2068 4346 2072
rect 4678 2068 4682 2072
rect 4734 2068 4738 2072
rect 5038 2068 5042 2072
rect 5190 2068 5194 2072
rect 5278 2068 5282 2072
rect 774 2058 778 2062
rect 902 2058 906 2062
rect 950 2058 954 2062
rect 1206 2058 1210 2062
rect 1230 2058 1234 2062
rect 1246 2058 1250 2062
rect 1326 2058 1330 2062
rect 1374 2058 1378 2062
rect 1422 2058 1426 2062
rect 1494 2058 1498 2062
rect 1694 2058 1698 2062
rect 1782 2058 1786 2062
rect 1854 2058 1858 2062
rect 2414 2058 2418 2062
rect 2702 2058 2706 2062
rect 2710 2058 2714 2062
rect 3286 2058 3290 2062
rect 3598 2058 3602 2062
rect 3726 2058 3730 2062
rect 3766 2058 3770 2062
rect 3894 2058 3898 2062
rect 4014 2058 4018 2062
rect 4094 2058 4098 2062
rect 4190 2058 4194 2062
rect 4614 2058 4618 2062
rect 4638 2058 4642 2062
rect 4670 2058 4674 2062
rect 4718 2058 4722 2062
rect 4990 2058 4994 2062
rect 5054 2058 5058 2062
rect 5078 2058 5082 2062
rect 246 2048 250 2052
rect 502 2048 506 2052
rect 630 2048 634 2052
rect 694 2048 698 2052
rect 902 2048 906 2052
rect 1182 2048 1186 2052
rect 1214 2048 1218 2052
rect 1918 2048 1922 2052
rect 1934 2048 1938 2052
rect 2014 2048 2018 2052
rect 2406 2048 2410 2052
rect 2958 2048 2962 2052
rect 3062 2048 3066 2052
rect 3222 2048 3226 2052
rect 3238 2048 3242 2052
rect 3366 2048 3370 2052
rect 3694 2048 3698 2052
rect 3726 2048 3730 2052
rect 3806 2048 3810 2052
rect 4238 2048 4242 2052
rect 558 2038 562 2042
rect 1142 2038 1146 2042
rect 4502 2048 4506 2052
rect 4510 2048 4514 2052
rect 4582 2048 4586 2052
rect 5014 2048 5018 2052
rect 2526 2038 2530 2042
rect 2926 2038 2930 2042
rect 3022 2038 3026 2042
rect 3070 2038 3074 2042
rect 3742 2038 3746 2042
rect 3854 2038 3858 2042
rect 3886 2038 3890 2042
rect 4142 2038 4146 2042
rect 4382 2038 4386 2042
rect 4518 2038 4522 2042
rect 374 2028 378 2032
rect 1102 2028 1106 2032
rect 1518 2028 1522 2032
rect 1942 2028 1946 2032
rect 2102 2028 2106 2032
rect 2254 2028 2258 2032
rect 2342 2028 2346 2032
rect 2574 2028 2578 2032
rect 4054 2028 4058 2032
rect 686 2018 690 2022
rect 1094 2018 1098 2022
rect 1334 2018 1338 2022
rect 1582 2018 1586 2022
rect 2294 2018 2298 2022
rect 2518 2018 2522 2022
rect 2854 2018 2858 2022
rect 2966 2018 2970 2022
rect 3390 2018 3394 2022
rect 5030 2018 5034 2022
rect 230 2008 234 2012
rect 1470 2008 1474 2012
rect 1686 2008 1690 2012
rect 2094 2008 2098 2012
rect 2126 2008 2130 2012
rect 2814 2008 2818 2012
rect 3102 2008 3106 2012
rect 3470 2008 3474 2012
rect 4398 2008 4402 2012
rect 4702 2008 4706 2012
rect 330 2003 334 2007
rect 338 2003 341 2007
rect 341 2003 342 2007
rect 1354 2003 1358 2007
rect 1362 2003 1365 2007
rect 1365 2003 1366 2007
rect 1254 1998 1258 2002
rect 2386 2003 2390 2007
rect 2394 2003 2397 2007
rect 2397 2003 2398 2007
rect 3402 2003 3406 2007
rect 3410 2003 3413 2007
rect 3413 2003 3414 2007
rect 4426 2003 4430 2007
rect 4434 2003 4437 2007
rect 4437 2003 4438 2007
rect 2686 1998 2690 2002
rect 3230 1998 3234 2002
rect 3254 1998 3258 2002
rect 3326 1998 3330 2002
rect 4078 1998 4082 2002
rect 4366 1998 4370 2002
rect 4718 1998 4722 2002
rect 4726 1998 4730 2002
rect 1462 1988 1466 1992
rect 1470 1988 1474 1992
rect 1830 1988 1834 1992
rect 1846 1988 1850 1992
rect 2094 1988 2098 1992
rect 2182 1988 2186 1992
rect 3526 1988 3530 1992
rect 4110 1988 4114 1992
rect 1190 1978 1194 1982
rect 1758 1978 1762 1982
rect 1998 1978 2002 1982
rect 3374 1978 3378 1982
rect 3478 1978 3482 1982
rect 3622 1978 3626 1982
rect 3686 1978 3690 1982
rect 4854 1978 4858 1982
rect 4870 1978 4874 1982
rect 4982 1978 4986 1982
rect 694 1968 698 1972
rect 1430 1968 1434 1972
rect 1438 1968 1442 1972
rect 1582 1968 1586 1972
rect 1606 1968 1610 1972
rect 1742 1968 1746 1972
rect 1750 1968 1754 1972
rect 1782 1968 1786 1972
rect 1814 1968 1818 1972
rect 2238 1968 2242 1972
rect 2414 1968 2418 1972
rect 2478 1968 2482 1972
rect 2542 1968 2546 1972
rect 2574 1968 2578 1972
rect 2766 1968 2770 1972
rect 2918 1968 2922 1972
rect 3030 1968 3034 1972
rect 3238 1968 3242 1972
rect 3422 1968 3426 1972
rect 3454 1968 3458 1972
rect 4414 1968 4418 1972
rect 4862 1968 4866 1972
rect 5022 1968 5026 1972
rect 406 1958 410 1962
rect 614 1958 618 1962
rect 894 1958 898 1962
rect 1206 1958 1210 1962
rect 1414 1958 1418 1962
rect 2006 1958 2010 1962
rect 2062 1958 2066 1962
rect 2078 1958 2082 1962
rect 2406 1958 2410 1962
rect 2678 1958 2682 1962
rect 3278 1958 3282 1962
rect 3422 1958 3426 1962
rect 3670 1958 3674 1962
rect 4318 1958 4322 1962
rect 4366 1958 4370 1962
rect 4710 1958 4714 1962
rect 318 1948 322 1952
rect 654 1948 658 1952
rect 1614 1948 1618 1952
rect 1622 1948 1626 1952
rect 1750 1948 1754 1952
rect 2126 1948 2130 1952
rect 2262 1948 2266 1952
rect 2502 1948 2506 1952
rect 2582 1948 2586 1952
rect 2774 1948 2778 1952
rect 3078 1948 3082 1952
rect 3406 1948 3410 1952
rect 3414 1948 3418 1952
rect 3606 1948 3610 1952
rect 582 1938 586 1942
rect 1318 1938 1322 1942
rect 1342 1938 1346 1942
rect 1502 1938 1506 1942
rect 1702 1938 1706 1942
rect 1718 1938 1722 1942
rect 1774 1938 1778 1942
rect 1854 1938 1858 1942
rect 1878 1938 1882 1942
rect 1910 1938 1914 1942
rect 1926 1938 1930 1942
rect 1966 1938 1970 1942
rect 2006 1938 2010 1942
rect 2086 1938 2090 1942
rect 2110 1938 2114 1942
rect 2574 1938 2578 1942
rect 2670 1938 2674 1942
rect 2702 1938 2706 1942
rect 2742 1938 2746 1942
rect 4550 1948 4554 1952
rect 5278 1948 5282 1952
rect 2910 1938 2914 1942
rect 3262 1938 3266 1942
rect 3550 1938 3554 1942
rect 4062 1938 4066 1942
rect 4078 1938 4082 1942
rect 4918 1938 4922 1942
rect 662 1928 666 1932
rect 1030 1928 1034 1932
rect 1142 1928 1146 1932
rect 1406 1928 1410 1932
rect 1582 1928 1586 1932
rect 1590 1928 1594 1932
rect 1694 1928 1698 1932
rect 1718 1928 1722 1932
rect 1742 1928 1746 1932
rect 1918 1928 1922 1932
rect 1942 1928 1946 1932
rect 2062 1928 2066 1932
rect 2254 1928 2258 1932
rect 2630 1928 2634 1932
rect 2790 1928 2794 1932
rect 3318 1928 3322 1932
rect 3678 1928 3682 1932
rect 3862 1928 3866 1932
rect 4094 1928 4098 1932
rect 4374 1928 4378 1932
rect 5006 1928 5010 1932
rect 5294 1928 5298 1932
rect 222 1918 226 1922
rect 1126 1918 1130 1922
rect 1190 1918 1194 1922
rect 2438 1918 2442 1922
rect 2862 1918 2866 1922
rect 2870 1918 2874 1922
rect 3894 1918 3898 1922
rect 4390 1918 4394 1922
rect 5094 1918 5098 1922
rect 5142 1918 5146 1922
rect 1862 1908 1866 1912
rect 2326 1908 2330 1912
rect 2718 1908 2722 1912
rect 4150 1908 4154 1912
rect 5070 1908 5074 1912
rect 850 1903 854 1907
rect 858 1903 861 1907
rect 861 1903 862 1907
rect 1874 1903 1878 1907
rect 1882 1903 1885 1907
rect 1885 1903 1886 1907
rect 1030 1898 1034 1902
rect 1118 1898 1122 1902
rect 1374 1898 1378 1902
rect 1422 1898 1426 1902
rect 1830 1898 1834 1902
rect 1934 1898 1938 1902
rect 2890 1903 2894 1907
rect 2898 1903 2901 1907
rect 2901 1903 2902 1907
rect 3922 1903 3926 1907
rect 3930 1903 3933 1907
rect 3933 1903 3934 1907
rect 4938 1903 4942 1907
rect 4946 1903 4949 1907
rect 4949 1903 4950 1907
rect 2214 1898 2218 1902
rect 2278 1898 2282 1902
rect 2486 1898 2490 1902
rect 3190 1898 3194 1902
rect 3278 1898 3282 1902
rect 3382 1898 3386 1902
rect 3598 1898 3602 1902
rect 3662 1898 3666 1902
rect 3942 1898 3946 1902
rect 3974 1898 3978 1902
rect 3990 1898 3994 1902
rect 4190 1898 4194 1902
rect 4846 1898 4850 1902
rect 710 1888 714 1892
rect 1086 1888 1090 1892
rect 1446 1888 1450 1892
rect 1862 1888 1866 1892
rect 2054 1888 2058 1892
rect 2070 1888 2074 1892
rect 2166 1888 2170 1892
rect 2286 1888 2290 1892
rect 2326 1888 2330 1892
rect 2470 1888 2474 1892
rect 2486 1888 2490 1892
rect 2582 1888 2586 1892
rect 4270 1888 4274 1892
rect 4310 1888 4314 1892
rect 270 1878 274 1882
rect 310 1878 314 1882
rect 366 1878 370 1882
rect 790 1878 794 1882
rect 1198 1878 1202 1882
rect 1206 1878 1210 1882
rect 1310 1878 1314 1882
rect 1454 1878 1458 1882
rect 2558 1878 2562 1882
rect 2766 1878 2770 1882
rect 3294 1878 3298 1882
rect 3574 1878 3578 1882
rect 3614 1878 3618 1882
rect 3782 1878 3786 1882
rect 3998 1878 4002 1882
rect 4014 1878 4018 1882
rect 4854 1888 4858 1892
rect 5118 1888 5122 1892
rect 5166 1888 5170 1892
rect 4534 1878 4538 1882
rect 4590 1878 4594 1882
rect 4822 1878 4826 1882
rect 686 1868 690 1872
rect 838 1868 842 1872
rect 1086 1868 1090 1872
rect 1318 1868 1322 1872
rect 1510 1868 1514 1872
rect 1862 1868 1866 1872
rect 1966 1868 1970 1872
rect 2190 1868 2194 1872
rect 2230 1868 2234 1872
rect 3046 1868 3050 1872
rect 3550 1868 3554 1872
rect 3638 1868 3642 1872
rect 3958 1868 3962 1872
rect 3974 1868 3978 1872
rect 4054 1868 4058 1872
rect 4158 1868 4162 1872
rect 4222 1868 4226 1872
rect 5254 1868 5258 1872
rect 214 1858 218 1862
rect 606 1858 610 1862
rect 678 1858 682 1862
rect 694 1858 698 1862
rect 718 1858 722 1862
rect 774 1858 778 1862
rect 926 1858 930 1862
rect 1294 1858 1298 1862
rect 1374 1858 1378 1862
rect 1758 1858 1762 1862
rect 2070 1858 2074 1862
rect 2326 1858 2330 1862
rect 2582 1858 2586 1862
rect 2790 1858 2794 1862
rect 3494 1858 3498 1862
rect 3654 1858 3658 1862
rect 3974 1858 3978 1862
rect 4246 1858 4250 1862
rect 4854 1858 4858 1862
rect 5038 1858 5042 1862
rect 5102 1858 5106 1862
rect 206 1848 210 1852
rect 358 1848 362 1852
rect 382 1848 386 1852
rect 646 1848 650 1852
rect 710 1848 714 1852
rect 766 1848 770 1852
rect 998 1848 1002 1852
rect 1566 1848 1570 1852
rect 1622 1848 1626 1852
rect 1630 1848 1634 1852
rect 1894 1848 1898 1852
rect 2502 1848 2506 1852
rect 2550 1848 2554 1852
rect 2662 1848 2666 1852
rect 2886 1848 2890 1852
rect 3142 1848 3146 1852
rect 3150 1848 3154 1852
rect 3222 1848 3226 1852
rect 3510 1848 3514 1852
rect 4014 1848 4018 1852
rect 4022 1848 4026 1852
rect 4670 1848 4674 1852
rect 4710 1848 4714 1852
rect 4790 1848 4794 1852
rect 4982 1848 4986 1852
rect 5038 1848 5042 1852
rect 230 1838 234 1842
rect 558 1838 562 1842
rect 1126 1838 1130 1842
rect 1686 1838 1690 1842
rect 2358 1838 2362 1842
rect 2518 1838 2522 1842
rect 2910 1838 2914 1842
rect 3710 1838 3714 1842
rect 4534 1838 4538 1842
rect 590 1828 594 1832
rect 1422 1828 1426 1832
rect 1646 1828 1650 1832
rect 1790 1828 1794 1832
rect 2150 1828 2154 1832
rect 2174 1828 2178 1832
rect 2686 1828 2690 1832
rect 2942 1828 2946 1832
rect 3046 1828 3050 1832
rect 3142 1828 3146 1832
rect 3406 1828 3410 1832
rect 3590 1828 3594 1832
rect 3862 1828 3866 1832
rect 3870 1828 3874 1832
rect 4214 1828 4218 1832
rect 4294 1828 4298 1832
rect 4318 1828 4322 1832
rect 4574 1828 4578 1832
rect 4854 1828 4858 1832
rect 2254 1818 2258 1822
rect 2286 1818 2290 1822
rect 3022 1818 3026 1822
rect 3030 1818 3034 1822
rect 3078 1818 3082 1822
rect 3358 1818 3362 1822
rect 3766 1818 3770 1822
rect 4166 1818 4170 1822
rect 4406 1818 4410 1822
rect 318 1808 322 1812
rect 774 1808 778 1812
rect 1006 1808 1010 1812
rect 1766 1808 1770 1812
rect 2038 1808 2042 1812
rect 2118 1808 2122 1812
rect 2318 1808 2322 1812
rect 2662 1808 2666 1812
rect 2710 1808 2714 1812
rect 2718 1808 2722 1812
rect 3382 1808 3386 1812
rect 330 1803 334 1807
rect 338 1803 341 1807
rect 341 1803 342 1807
rect 1354 1803 1358 1807
rect 1362 1803 1365 1807
rect 1365 1803 1366 1807
rect 2386 1803 2390 1807
rect 2394 1803 2397 1807
rect 2397 1803 2398 1807
rect 3402 1803 3406 1807
rect 3410 1803 3413 1807
rect 3413 1803 3414 1807
rect 4426 1803 4430 1807
rect 4434 1803 4437 1807
rect 4437 1803 4438 1807
rect 518 1798 522 1802
rect 1134 1798 1138 1802
rect 1558 1798 1562 1802
rect 2150 1798 2154 1802
rect 2446 1798 2450 1802
rect 2950 1798 2954 1802
rect 3030 1798 3034 1802
rect 3070 1798 3074 1802
rect 3582 1798 3586 1802
rect 4182 1798 4186 1802
rect 4710 1798 4714 1802
rect 166 1788 170 1792
rect 782 1788 786 1792
rect 2542 1788 2546 1792
rect 2630 1788 2634 1792
rect 3726 1788 3730 1792
rect 4662 1788 4666 1792
rect 726 1778 730 1782
rect 838 1778 842 1782
rect 1494 1778 1498 1782
rect 2046 1778 2050 1782
rect 2750 1778 2754 1782
rect 3110 1778 3114 1782
rect 3966 1778 3970 1782
rect 4350 1778 4354 1782
rect 4726 1778 4730 1782
rect 566 1768 570 1772
rect 726 1768 730 1772
rect 1198 1768 1202 1772
rect 1566 1768 1570 1772
rect 1814 1768 1818 1772
rect 2174 1768 2178 1772
rect 2198 1768 2202 1772
rect 2606 1768 2610 1772
rect 2846 1768 2850 1772
rect 2862 1768 2866 1772
rect 3182 1768 3186 1772
rect 4086 1768 4090 1772
rect 4350 1768 4354 1772
rect 374 1758 378 1762
rect 414 1758 418 1762
rect 1654 1758 1658 1762
rect 1718 1758 1722 1762
rect 1742 1758 1746 1762
rect 1990 1758 1994 1762
rect 2246 1758 2250 1762
rect 2486 1758 2490 1762
rect 2510 1758 2514 1762
rect 2934 1758 2938 1762
rect 3038 1758 3042 1762
rect 4142 1758 4146 1762
rect 4174 1758 4178 1762
rect 4222 1758 4226 1762
rect 4270 1758 4274 1762
rect 4454 1758 4458 1762
rect 4710 1758 4714 1762
rect 5094 1758 5098 1762
rect 582 1748 586 1752
rect 598 1748 602 1752
rect 742 1748 746 1752
rect 982 1748 986 1752
rect 1382 1748 1386 1752
rect 1406 1748 1410 1752
rect 1422 1748 1426 1752
rect 1566 1748 1570 1752
rect 2030 1748 2034 1752
rect 2134 1748 2138 1752
rect 2534 1748 2538 1752
rect 2886 1748 2890 1752
rect 3118 1748 3122 1752
rect 3262 1748 3266 1752
rect 3302 1748 3306 1752
rect 3550 1748 3554 1752
rect 3982 1748 3986 1752
rect 4190 1748 4194 1752
rect 4614 1748 4618 1752
rect 5062 1748 5066 1752
rect 726 1738 730 1742
rect 1150 1738 1154 1742
rect 1326 1738 1330 1742
rect 1574 1738 1578 1742
rect 1942 1738 1946 1742
rect 2174 1738 2178 1742
rect 2574 1738 2578 1742
rect 2582 1738 2586 1742
rect 3142 1738 3146 1742
rect 3942 1738 3946 1742
rect 4270 1738 4274 1742
rect 4502 1738 4506 1742
rect 4606 1738 4610 1742
rect 4894 1738 4898 1742
rect 5094 1738 5098 1742
rect 1670 1728 1674 1732
rect 1782 1728 1786 1732
rect 2102 1728 2106 1732
rect 3246 1728 3250 1732
rect 3502 1728 3506 1732
rect 3638 1728 3642 1732
rect 3854 1728 3858 1732
rect 1430 1718 1434 1722
rect 1822 1718 1826 1722
rect 2510 1718 2514 1722
rect 2542 1718 2546 1722
rect 2614 1718 2618 1722
rect 4166 1718 4170 1722
rect 4238 1718 4242 1722
rect 4310 1718 4314 1722
rect 4342 1718 4346 1722
rect 5126 1718 5130 1722
rect 1622 1708 1626 1712
rect 1958 1708 1962 1712
rect 2518 1708 2522 1712
rect 2670 1708 2674 1712
rect 3022 1708 3026 1712
rect 3382 1708 3386 1712
rect 850 1703 854 1707
rect 858 1703 861 1707
rect 861 1703 862 1707
rect 1874 1703 1878 1707
rect 1882 1703 1885 1707
rect 1885 1703 1886 1707
rect 2890 1703 2894 1707
rect 2898 1703 2901 1707
rect 2901 1703 2902 1707
rect 3922 1703 3926 1707
rect 3930 1703 3933 1707
rect 3933 1703 3934 1707
rect 4938 1703 4942 1707
rect 4946 1703 4949 1707
rect 4949 1703 4950 1707
rect 1118 1698 1122 1702
rect 2038 1698 2042 1702
rect 2566 1698 2570 1702
rect 2870 1698 2874 1702
rect 3014 1698 3018 1702
rect 3102 1698 3106 1702
rect 3150 1698 3154 1702
rect 3654 1698 3658 1702
rect 3902 1698 3906 1702
rect 4598 1698 4602 1702
rect 1990 1688 1994 1692
rect 2054 1688 2058 1692
rect 2606 1688 2610 1692
rect 2758 1688 2762 1692
rect 2910 1688 2914 1692
rect 3166 1688 3170 1692
rect 3238 1688 3242 1692
rect 3550 1688 3554 1692
rect 4022 1688 4026 1692
rect 4070 1688 4074 1692
rect 5206 1688 5210 1692
rect 5238 1688 5242 1692
rect 126 1678 130 1682
rect 566 1678 570 1682
rect 1198 1678 1202 1682
rect 1310 1678 1314 1682
rect 1566 1678 1570 1682
rect 1726 1678 1730 1682
rect 1782 1678 1786 1682
rect 2486 1678 2490 1682
rect 2846 1678 2850 1682
rect 2998 1678 3002 1682
rect 4174 1678 4178 1682
rect 4926 1678 4930 1682
rect 4974 1678 4978 1682
rect 5006 1678 5010 1682
rect 5238 1678 5242 1682
rect 454 1668 458 1672
rect 902 1668 906 1672
rect 918 1668 922 1672
rect 1206 1668 1210 1672
rect 1502 1668 1506 1672
rect 1582 1668 1586 1672
rect 1646 1668 1650 1672
rect 1686 1668 1690 1672
rect 2534 1668 2538 1672
rect 3078 1668 3082 1672
rect 3222 1668 3226 1672
rect 3238 1668 3242 1672
rect 3654 1668 3658 1672
rect 5166 1668 5170 1672
rect 286 1658 290 1662
rect 566 1658 570 1662
rect 1142 1658 1146 1662
rect 1422 1658 1426 1662
rect 2182 1658 2186 1662
rect 2486 1658 2490 1662
rect 2622 1658 2626 1662
rect 2646 1658 2650 1662
rect 2678 1658 2682 1662
rect 2718 1658 2722 1662
rect 3006 1658 3010 1662
rect 3150 1658 3154 1662
rect 3214 1658 3218 1662
rect 3406 1658 3410 1662
rect 3446 1658 3450 1662
rect 3654 1658 3658 1662
rect 4150 1658 4154 1662
rect 4198 1658 4202 1662
rect 4454 1658 4458 1662
rect 4494 1658 4498 1662
rect 4686 1658 4690 1662
rect 4718 1658 4722 1662
rect 4878 1658 4882 1662
rect 5174 1658 5178 1662
rect 5262 1658 5266 1662
rect 310 1648 314 1652
rect 806 1648 810 1652
rect 1326 1648 1330 1652
rect 1534 1648 1538 1652
rect 1670 1648 1674 1652
rect 1750 1648 1754 1652
rect 1814 1648 1818 1652
rect 2014 1648 2018 1652
rect 2126 1648 2130 1652
rect 2758 1648 2762 1652
rect 3110 1648 3114 1652
rect 3326 1648 3330 1652
rect 3374 1648 3378 1652
rect 3390 1648 3394 1652
rect 3646 1648 3650 1652
rect 4094 1648 4098 1652
rect 4646 1648 4650 1652
rect 4862 1648 4866 1652
rect 182 1638 186 1642
rect 446 1638 450 1642
rect 566 1638 570 1642
rect 582 1638 586 1642
rect 2070 1638 2074 1642
rect 2086 1638 2090 1642
rect 2958 1638 2962 1642
rect 3150 1638 3154 1642
rect 4238 1638 4242 1642
rect 1630 1628 1634 1632
rect 1854 1628 1858 1632
rect 3094 1628 3098 1632
rect 4630 1628 4634 1632
rect 4654 1628 4658 1632
rect 390 1618 394 1622
rect 406 1618 410 1622
rect 686 1618 690 1622
rect 2142 1618 2146 1622
rect 2438 1618 2442 1622
rect 2878 1618 2882 1622
rect 3310 1618 3314 1622
rect 4062 1618 4066 1622
rect 4406 1618 4410 1622
rect 1398 1608 1402 1612
rect 2374 1608 2378 1612
rect 2654 1608 2658 1612
rect 2854 1608 2858 1612
rect 3142 1608 3146 1612
rect 4142 1608 4146 1612
rect 4566 1608 4570 1612
rect 330 1603 334 1607
rect 338 1603 341 1607
rect 341 1603 342 1607
rect 1354 1603 1358 1607
rect 1362 1603 1365 1607
rect 1365 1603 1366 1607
rect 694 1598 698 1602
rect 1126 1598 1130 1602
rect 2386 1603 2390 1607
rect 2394 1603 2397 1607
rect 2397 1603 2398 1607
rect 3402 1603 3406 1607
rect 3410 1603 3413 1607
rect 3413 1603 3414 1607
rect 4426 1603 4430 1607
rect 4434 1603 4437 1607
rect 4437 1603 4438 1607
rect 1790 1598 1794 1602
rect 1950 1598 1954 1602
rect 2270 1598 2274 1602
rect 2926 1598 2930 1602
rect 4022 1598 4026 1602
rect 1022 1588 1026 1592
rect 2470 1588 2474 1592
rect 2790 1588 2794 1592
rect 3030 1588 3034 1592
rect 3774 1588 3778 1592
rect 3846 1588 3850 1592
rect 4278 1588 4282 1592
rect 1566 1578 1570 1582
rect 1718 1578 1722 1582
rect 1814 1578 1818 1582
rect 4614 1578 4618 1582
rect 4670 1578 4674 1582
rect 670 1568 674 1572
rect 1054 1568 1058 1572
rect 1454 1568 1458 1572
rect 1462 1568 1466 1572
rect 1830 1568 1834 1572
rect 3022 1568 3026 1572
rect 3366 1568 3370 1572
rect 3422 1568 3426 1572
rect 3838 1568 3842 1572
rect 3902 1568 3906 1572
rect 4102 1568 4106 1572
rect 4238 1568 4242 1572
rect 4334 1568 4338 1572
rect 4566 1568 4570 1572
rect 4598 1568 4602 1572
rect 4654 1568 4658 1572
rect 4702 1568 4706 1572
rect 4766 1568 4770 1572
rect 4926 1568 4930 1572
rect 5262 1568 5266 1572
rect 678 1558 682 1562
rect 1118 1558 1122 1562
rect 1422 1558 1426 1562
rect 1486 1558 1490 1562
rect 1502 1558 1506 1562
rect 1718 1558 1722 1562
rect 1742 1558 1746 1562
rect 1862 1558 1866 1562
rect 1990 1558 1994 1562
rect 2054 1558 2058 1562
rect 2110 1558 2114 1562
rect 2358 1558 2362 1562
rect 3542 1558 3546 1562
rect 4158 1558 4162 1562
rect 4470 1558 4474 1562
rect 4582 1558 4586 1562
rect 4694 1558 4698 1562
rect 150 1548 154 1552
rect 406 1548 410 1552
rect 470 1548 474 1552
rect 622 1548 626 1552
rect 654 1548 658 1552
rect 734 1548 738 1552
rect 758 1548 762 1552
rect 806 1548 810 1552
rect 1014 1548 1018 1552
rect 1166 1548 1170 1552
rect 1638 1548 1642 1552
rect 1974 1548 1978 1552
rect 1998 1548 2002 1552
rect 2918 1548 2922 1552
rect 2950 1548 2954 1552
rect 3270 1548 3274 1552
rect 3350 1548 3354 1552
rect 3814 1548 3818 1552
rect 3846 1548 3850 1552
rect 3886 1548 3890 1552
rect 3902 1548 3906 1552
rect 4302 1548 4306 1552
rect 4318 1548 4322 1552
rect 4598 1548 4602 1552
rect 4622 1548 4626 1552
rect 4862 1548 4866 1552
rect 5030 1548 5034 1552
rect 5062 1548 5066 1552
rect 142 1538 146 1542
rect 526 1538 530 1542
rect 582 1538 586 1542
rect 646 1538 650 1542
rect 662 1538 666 1542
rect 750 1538 754 1542
rect 1126 1538 1130 1542
rect 1470 1538 1474 1542
rect 1526 1538 1530 1542
rect 1542 1538 1546 1542
rect 1742 1538 1746 1542
rect 1934 1538 1938 1542
rect 1990 1538 1994 1542
rect 2486 1538 2490 1542
rect 2798 1538 2802 1542
rect 2814 1538 2818 1542
rect 3078 1538 3082 1542
rect 3086 1538 3090 1542
rect 3102 1538 3106 1542
rect 3118 1538 3122 1542
rect 3262 1538 3266 1542
rect 3494 1538 3498 1542
rect 3630 1538 3634 1542
rect 3694 1538 3698 1542
rect 4110 1538 4114 1542
rect 4150 1538 4154 1542
rect 4190 1538 4194 1542
rect 4246 1538 4250 1542
rect 4374 1538 4378 1542
rect 4398 1538 4402 1542
rect 4494 1538 4498 1542
rect 214 1528 218 1532
rect 558 1528 562 1532
rect 1430 1528 1434 1532
rect 1766 1528 1770 1532
rect 1894 1528 1898 1532
rect 2006 1528 2010 1532
rect 2118 1528 2122 1532
rect 2518 1528 2522 1532
rect 4638 1528 4642 1532
rect 5006 1528 5010 1532
rect 5046 1528 5050 1532
rect 5238 1528 5242 1532
rect 598 1518 602 1522
rect 1726 1518 1730 1522
rect 2078 1518 2082 1522
rect 3014 1518 3018 1522
rect 4110 1518 4114 1522
rect 4718 1518 4722 1522
rect 366 1508 370 1512
rect 1902 1508 1906 1512
rect 2574 1508 2578 1512
rect 2814 1508 2818 1512
rect 2910 1508 2914 1512
rect 3006 1508 3010 1512
rect 3062 1508 3066 1512
rect 4102 1508 4106 1512
rect 4222 1508 4226 1512
rect 4270 1508 4274 1512
rect 4358 1508 4362 1512
rect 4406 1508 4410 1512
rect 4502 1508 4506 1512
rect 4694 1508 4698 1512
rect 850 1503 854 1507
rect 858 1503 861 1507
rect 861 1503 862 1507
rect 1874 1503 1878 1507
rect 1882 1503 1885 1507
rect 1885 1503 1886 1507
rect 2890 1503 2894 1507
rect 2898 1503 2901 1507
rect 2901 1503 2902 1507
rect 3922 1503 3926 1507
rect 3930 1503 3933 1507
rect 3933 1503 3934 1507
rect 4938 1503 4942 1507
rect 4946 1503 4949 1507
rect 4949 1503 4950 1507
rect 214 1498 218 1502
rect 710 1498 714 1502
rect 1494 1498 1498 1502
rect 1758 1498 1762 1502
rect 1926 1498 1930 1502
rect 1958 1498 1962 1502
rect 2046 1498 2050 1502
rect 2062 1498 2066 1502
rect 2198 1498 2202 1502
rect 3022 1498 3026 1502
rect 3038 1498 3042 1502
rect 3286 1498 3290 1502
rect 4566 1498 4570 1502
rect 4622 1498 4626 1502
rect 990 1488 994 1492
rect 1334 1488 1338 1492
rect 1566 1488 1570 1492
rect 1678 1488 1682 1492
rect 1702 1488 1706 1492
rect 2102 1488 2106 1492
rect 2446 1488 2450 1492
rect 4350 1488 4354 1492
rect 4382 1488 4386 1492
rect 4734 1488 4738 1492
rect 5062 1488 5066 1492
rect 454 1478 458 1482
rect 1822 1478 1826 1482
rect 2134 1478 2138 1482
rect 2454 1478 2458 1482
rect 2590 1478 2594 1482
rect 3262 1478 3266 1482
rect 3286 1478 3290 1482
rect 3302 1478 3306 1482
rect 3870 1478 3874 1482
rect 4054 1478 4058 1482
rect 4246 1478 4250 1482
rect 4526 1478 4530 1482
rect 5182 1478 5186 1482
rect 230 1468 234 1472
rect 302 1468 306 1472
rect 614 1468 618 1472
rect 798 1468 802 1472
rect 926 1468 930 1472
rect 1270 1468 1274 1472
rect 1374 1468 1378 1472
rect 1566 1468 1570 1472
rect 1638 1468 1642 1472
rect 1678 1468 1682 1472
rect 1726 1468 1730 1472
rect 1742 1468 1746 1472
rect 1758 1468 1762 1472
rect 1782 1468 1786 1472
rect 1926 1468 1930 1472
rect 2078 1468 2082 1472
rect 3390 1468 3394 1472
rect 3654 1468 3658 1472
rect 4166 1468 4170 1472
rect 4182 1468 4186 1472
rect 4310 1468 4314 1472
rect 4494 1468 4498 1472
rect 4558 1468 4562 1472
rect 4782 1468 4786 1472
rect 4934 1468 4938 1472
rect 5190 1468 5194 1472
rect 390 1458 394 1462
rect 510 1458 514 1462
rect 622 1458 626 1462
rect 870 1458 874 1462
rect 1110 1458 1114 1462
rect 1166 1458 1170 1462
rect 1254 1458 1258 1462
rect 1278 1458 1282 1462
rect 1390 1458 1394 1462
rect 1446 1458 1450 1462
rect 1486 1458 1490 1462
rect 1502 1458 1506 1462
rect 1846 1458 1850 1462
rect 1886 1458 1890 1462
rect 1910 1458 1914 1462
rect 1942 1458 1946 1462
rect 2454 1458 2458 1462
rect 2542 1458 2546 1462
rect 2758 1458 2762 1462
rect 2966 1458 2970 1462
rect 3110 1458 3114 1462
rect 3646 1458 3650 1462
rect 3966 1458 3970 1462
rect 4270 1458 4274 1462
rect 4470 1458 4474 1462
rect 4806 1458 4810 1462
rect 5166 1458 5170 1462
rect 5182 1458 5186 1462
rect 406 1448 410 1452
rect 414 1448 418 1452
rect 582 1448 586 1452
rect 1262 1448 1266 1452
rect 1278 1448 1282 1452
rect 1654 1448 1658 1452
rect 1702 1448 1706 1452
rect 1718 1448 1722 1452
rect 1942 1448 1946 1452
rect 2222 1448 2226 1452
rect 2462 1448 2466 1452
rect 2862 1448 2866 1452
rect 3390 1448 3394 1452
rect 3614 1448 3618 1452
rect 3854 1448 3858 1452
rect 4398 1448 4402 1452
rect 174 1438 178 1442
rect 334 1438 338 1442
rect 694 1438 698 1442
rect 1734 1438 1738 1442
rect 1790 1438 1794 1442
rect 1902 1438 1906 1442
rect 1966 1438 1970 1442
rect 2006 1438 2010 1442
rect 2134 1438 2138 1442
rect 2990 1438 2994 1442
rect 3102 1438 3106 1442
rect 3110 1438 3114 1442
rect 5110 1438 5114 1442
rect 5198 1438 5202 1442
rect 582 1428 586 1432
rect 774 1428 778 1432
rect 1374 1428 1378 1432
rect 1390 1428 1394 1432
rect 1574 1428 1578 1432
rect 1590 1428 1594 1432
rect 1830 1428 1834 1432
rect 2070 1428 2074 1432
rect 2582 1428 2586 1432
rect 3358 1428 3362 1432
rect 4054 1428 4058 1432
rect 5030 1428 5034 1432
rect 1022 1418 1026 1422
rect 1182 1418 1186 1422
rect 2126 1418 2130 1422
rect 2766 1418 2770 1422
rect 3854 1418 3858 1422
rect 4558 1418 4562 1422
rect 4750 1418 4754 1422
rect 4774 1418 4778 1422
rect 4814 1418 4818 1422
rect 5158 1418 5162 1422
rect 1030 1408 1034 1412
rect 1222 1408 1226 1412
rect 1318 1408 1322 1412
rect 2270 1408 2274 1412
rect 2974 1408 2978 1412
rect 3518 1408 3522 1412
rect 4454 1408 4458 1412
rect 330 1403 334 1407
rect 338 1403 341 1407
rect 341 1403 342 1407
rect 1354 1403 1358 1407
rect 1362 1403 1365 1407
rect 1365 1403 1366 1407
rect 2386 1403 2390 1407
rect 2394 1403 2397 1407
rect 2397 1403 2398 1407
rect 3402 1403 3406 1407
rect 3410 1403 3413 1407
rect 3413 1403 3414 1407
rect 4426 1403 4430 1407
rect 4434 1403 4437 1407
rect 4437 1403 4438 1407
rect 2286 1398 2290 1402
rect 2470 1398 2474 1402
rect 2542 1398 2546 1402
rect 3214 1398 3218 1402
rect 3526 1398 3530 1402
rect 3942 1398 3946 1402
rect 4382 1398 4386 1402
rect 4542 1398 4546 1402
rect 5046 1398 5050 1402
rect 654 1388 658 1392
rect 1166 1388 1170 1392
rect 3086 1388 3090 1392
rect 3742 1388 3746 1392
rect 4718 1388 4722 1392
rect 4750 1388 4754 1392
rect 990 1378 994 1382
rect 1342 1378 1346 1382
rect 2214 1378 2218 1382
rect 2870 1378 2874 1382
rect 3078 1378 3082 1382
rect 3542 1378 3546 1382
rect 3598 1378 3602 1382
rect 3750 1378 3754 1382
rect 3966 1378 3970 1382
rect 4510 1378 4514 1382
rect 4966 1378 4970 1382
rect 2238 1368 2242 1372
rect 2342 1368 2346 1372
rect 2950 1368 2954 1372
rect 3294 1368 3298 1372
rect 3390 1368 3394 1372
rect 3790 1368 3794 1372
rect 1014 1358 1018 1362
rect 1462 1358 1466 1362
rect 1982 1358 1986 1362
rect 2046 1358 2050 1362
rect 2518 1358 2522 1362
rect 2534 1358 2538 1362
rect 2798 1358 2802 1362
rect 3054 1358 3058 1362
rect 3350 1358 3354 1362
rect 3678 1358 3682 1362
rect 4222 1358 4226 1362
rect 4414 1358 4418 1362
rect 4470 1358 4474 1362
rect 4510 1358 4514 1362
rect 4574 1358 4578 1362
rect 4606 1358 4610 1362
rect 4622 1358 4626 1362
rect 4766 1358 4770 1362
rect 4814 1358 4818 1362
rect 5126 1358 5130 1362
rect 262 1348 266 1352
rect 390 1348 394 1352
rect 518 1348 522 1352
rect 1054 1348 1058 1352
rect 1214 1348 1218 1352
rect 1582 1348 1586 1352
rect 1694 1348 1698 1352
rect 1718 1348 1722 1352
rect 1790 1348 1794 1352
rect 2030 1348 2034 1352
rect 2094 1348 2098 1352
rect 2558 1348 2562 1352
rect 2582 1348 2586 1352
rect 2702 1348 2706 1352
rect 2966 1348 2970 1352
rect 2998 1348 3002 1352
rect 3158 1348 3162 1352
rect 4014 1348 4018 1352
rect 4222 1348 4226 1352
rect 4382 1348 4386 1352
rect 4614 1348 4618 1352
rect 4718 1348 4722 1352
rect 4758 1348 4762 1352
rect 5070 1348 5074 1352
rect 5094 1348 5098 1352
rect 5166 1348 5170 1352
rect 246 1338 250 1342
rect 422 1338 426 1342
rect 1014 1338 1018 1342
rect 1062 1338 1066 1342
rect 1606 1338 1610 1342
rect 1782 1338 1786 1342
rect 1854 1338 1858 1342
rect 1966 1338 1970 1342
rect 1982 1338 1986 1342
rect 1998 1338 2002 1342
rect 2222 1338 2226 1342
rect 2414 1338 2418 1342
rect 3358 1338 3362 1342
rect 3902 1338 3906 1342
rect 4054 1338 4058 1342
rect 4310 1338 4314 1342
rect 4406 1338 4410 1342
rect 4606 1338 4610 1342
rect 4646 1338 4650 1342
rect 4774 1338 4778 1342
rect 4918 1338 4922 1342
rect 5102 1338 5106 1342
rect 5182 1338 5186 1342
rect 526 1328 530 1332
rect 774 1328 778 1332
rect 1246 1328 1250 1332
rect 1526 1328 1530 1332
rect 1654 1328 1658 1332
rect 1942 1328 1946 1332
rect 1958 1328 1962 1332
rect 2022 1328 2026 1332
rect 2262 1328 2266 1332
rect 2310 1328 2314 1332
rect 2334 1328 2338 1332
rect 2406 1328 2410 1332
rect 3558 1328 3562 1332
rect 3582 1328 3586 1332
rect 4278 1328 4282 1332
rect 790 1318 794 1322
rect 1742 1318 1746 1322
rect 2326 1318 2330 1322
rect 2446 1318 2450 1322
rect 3238 1318 3242 1322
rect 3302 1318 3306 1322
rect 3590 1318 3594 1322
rect 3854 1318 3858 1322
rect 4270 1318 4274 1322
rect 4742 1318 4746 1322
rect 5030 1318 5034 1322
rect 5118 1318 5122 1322
rect 126 1308 130 1312
rect 974 1308 978 1312
rect 1070 1308 1074 1312
rect 1558 1308 1562 1312
rect 1838 1308 1842 1312
rect 2502 1308 2506 1312
rect 3158 1308 3162 1312
rect 3766 1308 3770 1312
rect 3814 1308 3818 1312
rect 4326 1308 4330 1312
rect 4390 1308 4394 1312
rect 5126 1308 5130 1312
rect 5198 1308 5202 1312
rect 850 1303 854 1307
rect 858 1303 861 1307
rect 861 1303 862 1307
rect 238 1298 242 1302
rect 1062 1298 1066 1302
rect 1874 1303 1878 1307
rect 1882 1303 1885 1307
rect 1885 1303 1886 1307
rect 2890 1303 2894 1307
rect 2898 1303 2901 1307
rect 2901 1303 2902 1307
rect 3922 1303 3926 1307
rect 3930 1303 3933 1307
rect 3933 1303 3934 1307
rect 4938 1303 4942 1307
rect 4946 1303 4949 1307
rect 4949 1303 4950 1307
rect 1614 1298 1618 1302
rect 1862 1298 1866 1302
rect 2070 1298 2074 1302
rect 3126 1298 3130 1302
rect 3134 1298 3138 1302
rect 3430 1298 3434 1302
rect 3830 1298 3834 1302
rect 3910 1298 3914 1302
rect 3990 1298 3994 1302
rect 4446 1298 4450 1302
rect 1166 1288 1170 1292
rect 1382 1288 1386 1292
rect 1814 1288 1818 1292
rect 1870 1288 1874 1292
rect 2046 1288 2050 1292
rect 2502 1288 2506 1292
rect 2774 1288 2778 1292
rect 2790 1288 2794 1292
rect 2862 1288 2866 1292
rect 3342 1288 3346 1292
rect 3782 1288 3786 1292
rect 230 1278 234 1282
rect 462 1278 466 1282
rect 870 1278 874 1282
rect 950 1278 954 1282
rect 1430 1278 1434 1282
rect 1926 1278 1930 1282
rect 2062 1278 2066 1282
rect 2406 1278 2410 1282
rect 2774 1278 2778 1282
rect 3358 1278 3362 1282
rect 3510 1278 3514 1282
rect 3870 1278 3874 1282
rect 3886 1278 3890 1282
rect 3990 1278 3994 1282
rect 4262 1278 4266 1282
rect 4286 1278 4290 1282
rect 4566 1278 4570 1282
rect 4814 1278 4818 1282
rect 5102 1278 5106 1282
rect 126 1268 130 1272
rect 286 1268 290 1272
rect 446 1268 450 1272
rect 838 1268 842 1272
rect 862 1268 866 1272
rect 958 1268 962 1272
rect 974 1268 978 1272
rect 1006 1268 1010 1272
rect 1302 1268 1306 1272
rect 1646 1268 1650 1272
rect 1910 1268 1914 1272
rect 2486 1268 2490 1272
rect 2814 1268 2818 1272
rect 3278 1268 3282 1272
rect 4030 1268 4034 1272
rect 4334 1268 4338 1272
rect 230 1258 234 1262
rect 406 1258 410 1262
rect 430 1258 434 1262
rect 814 1258 818 1262
rect 1006 1258 1010 1262
rect 1454 1258 1458 1262
rect 1678 1258 1682 1262
rect 2406 1258 2410 1262
rect 2454 1258 2458 1262
rect 2478 1258 2482 1262
rect 2518 1258 2522 1262
rect 2542 1258 2546 1262
rect 2782 1258 2786 1262
rect 2950 1258 2954 1262
rect 2998 1258 3002 1262
rect 3222 1258 3226 1262
rect 3246 1258 3250 1262
rect 3294 1258 3298 1262
rect 3342 1258 3346 1262
rect 3758 1258 3762 1262
rect 4078 1258 4082 1262
rect 4110 1258 4114 1262
rect 4326 1258 4330 1262
rect 4446 1258 4450 1262
rect 4534 1258 4538 1262
rect 4686 1258 4690 1262
rect 5182 1258 5186 1262
rect 1190 1248 1194 1252
rect 1374 1248 1378 1252
rect 1478 1248 1482 1252
rect 1566 1248 1570 1252
rect 1838 1248 1842 1252
rect 1918 1248 1922 1252
rect 1958 1248 1962 1252
rect 2022 1248 2026 1252
rect 2302 1248 2306 1252
rect 2686 1248 2690 1252
rect 2718 1248 2722 1252
rect 3942 1248 3946 1252
rect 4174 1248 4178 1252
rect 4342 1248 4346 1252
rect 4390 1248 4394 1252
rect 4398 1248 4402 1252
rect 4910 1248 4914 1252
rect 4918 1248 4922 1252
rect 4934 1248 4938 1252
rect 310 1238 314 1242
rect 1446 1238 1450 1242
rect 2774 1238 2778 1242
rect 3270 1238 3274 1242
rect 3726 1238 3730 1242
rect 3742 1238 3746 1242
rect 3094 1228 3098 1232
rect 3974 1228 3978 1232
rect 5086 1228 5090 1232
rect 158 1218 162 1222
rect 742 1218 746 1222
rect 902 1218 906 1222
rect 958 1218 962 1222
rect 1990 1218 1994 1222
rect 2550 1218 2554 1222
rect 2622 1218 2626 1222
rect 3150 1218 3154 1222
rect 3494 1218 3498 1222
rect 3990 1218 3994 1222
rect 4894 1218 4898 1222
rect 1174 1208 1178 1212
rect 1406 1208 1410 1212
rect 1894 1208 1898 1212
rect 2838 1208 2842 1212
rect 2878 1208 2882 1212
rect 2958 1208 2962 1212
rect 3030 1208 3034 1212
rect 3070 1208 3074 1212
rect 3326 1208 3330 1212
rect 5102 1208 5106 1212
rect 330 1203 334 1207
rect 338 1203 341 1207
rect 341 1203 342 1207
rect 1354 1203 1358 1207
rect 1362 1203 1365 1207
rect 1365 1203 1366 1207
rect 2386 1203 2390 1207
rect 2394 1203 2397 1207
rect 2397 1203 2398 1207
rect 3402 1203 3406 1207
rect 3410 1203 3413 1207
rect 3413 1203 3414 1207
rect 4426 1203 4430 1207
rect 4434 1203 4437 1207
rect 4437 1203 4438 1207
rect 1310 1198 1314 1202
rect 1398 1198 1402 1202
rect 1862 1198 1866 1202
rect 2478 1198 2482 1202
rect 2670 1198 2674 1202
rect 3182 1198 3186 1202
rect 3238 1198 3242 1202
rect 4302 1198 4306 1202
rect 4454 1198 4458 1202
rect 5086 1198 5090 1202
rect 886 1188 890 1192
rect 1414 1188 1418 1192
rect 2046 1188 2050 1192
rect 2078 1188 2082 1192
rect 4326 1188 4330 1192
rect 5230 1188 5234 1192
rect 222 1178 226 1182
rect 606 1178 610 1182
rect 1158 1178 1162 1182
rect 1854 1178 1858 1182
rect 2582 1178 2586 1182
rect 2598 1178 2602 1182
rect 2838 1178 2842 1182
rect 3230 1178 3234 1182
rect 3558 1178 3562 1182
rect 3630 1178 3634 1182
rect 4550 1178 4554 1182
rect 958 1168 962 1172
rect 2270 1168 2274 1172
rect 2574 1168 2578 1172
rect 3030 1168 3034 1172
rect 3814 1168 3818 1172
rect 5166 1168 5170 1172
rect 5198 1168 5202 1172
rect 270 1158 274 1162
rect 414 1158 418 1162
rect 718 1158 722 1162
rect 894 1158 898 1162
rect 1214 1158 1218 1162
rect 1334 1158 1338 1162
rect 2094 1158 2098 1162
rect 2318 1158 2322 1162
rect 2478 1158 2482 1162
rect 2942 1158 2946 1162
rect 3022 1158 3026 1162
rect 3110 1158 3114 1162
rect 3318 1158 3322 1162
rect 3550 1158 3554 1162
rect 3574 1158 3578 1162
rect 3630 1158 3634 1162
rect 3806 1158 3810 1162
rect 4006 1158 4010 1162
rect 4022 1158 4026 1162
rect 5190 1158 5194 1162
rect 406 1148 410 1152
rect 718 1148 722 1152
rect 814 1148 818 1152
rect 822 1148 826 1152
rect 838 1148 842 1152
rect 934 1148 938 1152
rect 1022 1148 1026 1152
rect 1374 1148 1378 1152
rect 1526 1148 1530 1152
rect 1614 1148 1618 1152
rect 2222 1148 2226 1152
rect 2254 1148 2258 1152
rect 2366 1148 2370 1152
rect 2566 1148 2570 1152
rect 2598 1148 2602 1152
rect 2734 1148 2738 1152
rect 3262 1148 3266 1152
rect 3334 1148 3338 1152
rect 3350 1148 3354 1152
rect 3358 1148 3362 1152
rect 3774 1148 3778 1152
rect 3782 1148 3786 1152
rect 4134 1148 4138 1152
rect 4166 1148 4170 1152
rect 4294 1148 4298 1152
rect 4542 1148 4546 1152
rect 4670 1148 4674 1152
rect 4734 1148 4738 1152
rect 4910 1148 4914 1152
rect 5118 1148 5122 1152
rect 5166 1148 5170 1152
rect 5286 1148 5290 1152
rect 126 1138 130 1142
rect 150 1138 154 1142
rect 2142 1138 2146 1142
rect 2446 1138 2450 1142
rect 2918 1138 2922 1142
rect 3022 1138 3026 1142
rect 3134 1138 3138 1142
rect 3182 1138 3186 1142
rect 3502 1138 3506 1142
rect 3510 1138 3514 1142
rect 3598 1138 3602 1142
rect 4638 1138 4642 1142
rect 4646 1138 4650 1142
rect 4894 1138 4898 1142
rect 4990 1138 4994 1142
rect 5054 1138 5058 1142
rect 5134 1138 5138 1142
rect 5150 1138 5154 1142
rect 406 1128 410 1132
rect 790 1128 794 1132
rect 950 1128 954 1132
rect 1166 1128 1170 1132
rect 1662 1128 1666 1132
rect 1814 1128 1818 1132
rect 2166 1128 2170 1132
rect 2174 1128 2178 1132
rect 2718 1128 2722 1132
rect 2814 1128 2818 1132
rect 3238 1128 3242 1132
rect 3262 1128 3266 1132
rect 3326 1128 3330 1132
rect 3334 1128 3338 1132
rect 3358 1128 3362 1132
rect 3958 1128 3962 1132
rect 4358 1128 4362 1132
rect 4590 1128 4594 1132
rect 4654 1128 4658 1132
rect 4750 1128 4754 1132
rect 574 1118 578 1122
rect 702 1118 706 1122
rect 1438 1118 1442 1122
rect 2118 1118 2122 1122
rect 2614 1118 2618 1122
rect 2982 1118 2986 1122
rect 3030 1118 3034 1122
rect 3150 1118 3154 1122
rect 3606 1118 3610 1122
rect 3726 1118 3730 1122
rect 3934 1118 3938 1122
rect 4366 1118 4370 1122
rect 4454 1118 4458 1122
rect 4934 1118 4938 1122
rect 4966 1118 4970 1122
rect 302 1108 306 1112
rect 830 1108 834 1112
rect 1294 1108 1298 1112
rect 1766 1108 1770 1112
rect 1838 1108 1842 1112
rect 2334 1108 2338 1112
rect 2870 1108 2874 1112
rect 2950 1108 2954 1112
rect 4766 1108 4770 1112
rect 5094 1108 5098 1112
rect 850 1103 854 1107
rect 858 1103 861 1107
rect 861 1103 862 1107
rect 1874 1103 1878 1107
rect 1882 1103 1885 1107
rect 1885 1103 1886 1107
rect 2890 1103 2894 1107
rect 2898 1103 2901 1107
rect 2901 1103 2902 1107
rect 3922 1103 3926 1107
rect 3930 1103 3933 1107
rect 3933 1103 3934 1107
rect 4938 1103 4942 1107
rect 4946 1103 4949 1107
rect 4949 1103 4950 1107
rect 182 1098 186 1102
rect 302 1098 306 1102
rect 766 1098 770 1102
rect 1214 1098 1218 1102
rect 2918 1098 2922 1102
rect 3374 1098 3378 1102
rect 4086 1098 4090 1102
rect 1638 1088 1642 1092
rect 2686 1088 2690 1092
rect 3958 1088 3962 1092
rect 4206 1088 4210 1092
rect 4774 1088 4778 1092
rect 5166 1088 5170 1092
rect 142 1078 146 1082
rect 750 1078 754 1082
rect 998 1078 1002 1082
rect 1070 1078 1074 1082
rect 1302 1078 1306 1082
rect 1798 1078 1802 1082
rect 2422 1078 2426 1082
rect 3070 1078 3074 1082
rect 3774 1078 3778 1082
rect 4678 1078 4682 1082
rect 4926 1078 4930 1082
rect 5158 1078 5162 1082
rect 686 1068 690 1072
rect 1854 1068 1858 1072
rect 2662 1068 2666 1072
rect 2686 1068 2690 1072
rect 2718 1068 2722 1072
rect 2726 1068 2730 1072
rect 3214 1068 3218 1072
rect 3302 1068 3306 1072
rect 3534 1068 3538 1072
rect 3750 1068 3754 1072
rect 4046 1068 4050 1072
rect 4182 1068 4186 1072
rect 4262 1068 4266 1072
rect 222 1058 226 1062
rect 910 1058 914 1062
rect 1022 1058 1026 1062
rect 1254 1058 1258 1062
rect 2574 1058 2578 1062
rect 2726 1058 2730 1062
rect 3350 1058 3354 1062
rect 3766 1058 3770 1062
rect 3998 1058 4002 1062
rect 4374 1068 4378 1072
rect 4534 1068 4538 1072
rect 4910 1068 4914 1072
rect 4230 1058 4234 1062
rect 4630 1058 4634 1062
rect 5062 1058 5066 1062
rect 838 1048 842 1052
rect 1190 1048 1194 1052
rect 1926 1048 1930 1052
rect 3542 1048 3546 1052
rect 3646 1048 3650 1052
rect 4134 1048 4138 1052
rect 4182 1048 4186 1052
rect 4398 1048 4402 1052
rect 4534 1048 4538 1052
rect 5118 1048 5122 1052
rect 358 1038 362 1042
rect 1238 1038 1242 1042
rect 2142 1038 2146 1042
rect 3214 1038 3218 1042
rect 3494 1038 3498 1042
rect 4150 1038 4154 1042
rect 4782 1038 4786 1042
rect 5110 1038 5114 1042
rect 550 1028 554 1032
rect 950 1028 954 1032
rect 1206 1028 1210 1032
rect 1278 1028 1282 1032
rect 2734 1028 2738 1032
rect 3510 1028 3514 1032
rect 4310 1028 4314 1032
rect 4486 1028 4490 1032
rect 846 1018 850 1022
rect 1054 1018 1058 1022
rect 2966 1018 2970 1022
rect 3886 1018 3890 1022
rect 4246 1018 4250 1022
rect 4262 1018 4266 1022
rect 5270 1018 5274 1022
rect 1294 1008 1298 1012
rect 1902 1008 1906 1012
rect 3174 1008 3178 1012
rect 3438 1008 3442 1012
rect 4758 1008 4762 1012
rect 5110 1008 5114 1012
rect 330 1003 334 1007
rect 338 1003 341 1007
rect 341 1003 342 1007
rect 1354 1003 1358 1007
rect 1362 1003 1365 1007
rect 1365 1003 1366 1007
rect 2386 1003 2390 1007
rect 2394 1003 2397 1007
rect 2397 1003 2398 1007
rect 3402 1003 3406 1007
rect 3410 1003 3413 1007
rect 3413 1003 3414 1007
rect 4426 1003 4430 1007
rect 4434 1003 4437 1007
rect 4437 1003 4438 1007
rect 222 998 226 1002
rect 470 998 474 1002
rect 1046 998 1050 1002
rect 1438 998 1442 1002
rect 1654 998 1658 1002
rect 2766 998 2770 1002
rect 4414 998 4418 1002
rect 4590 998 4594 1002
rect 5270 998 5274 1002
rect 942 988 946 992
rect 1030 988 1034 992
rect 1318 988 1322 992
rect 1462 988 1466 992
rect 2126 988 2130 992
rect 2582 988 2586 992
rect 3958 988 3962 992
rect 4238 988 4242 992
rect 4446 988 4450 992
rect 830 978 834 982
rect 1918 978 1922 982
rect 2558 978 2562 982
rect 2710 978 2714 982
rect 3046 978 3050 982
rect 3750 978 3754 982
rect 4126 978 4130 982
rect 942 968 946 972
rect 998 968 1002 972
rect 1518 968 1522 972
rect 3494 968 3498 972
rect 3734 968 3738 972
rect 3790 968 3794 972
rect 4710 968 4714 972
rect 5278 968 5282 972
rect 182 958 186 962
rect 318 958 322 962
rect 702 958 706 962
rect 846 958 850 962
rect 982 958 986 962
rect 1022 958 1026 962
rect 1286 958 1290 962
rect 2134 958 2138 962
rect 2334 958 2338 962
rect 2646 958 2650 962
rect 2702 958 2706 962
rect 2758 958 2762 962
rect 2790 958 2794 962
rect 3166 958 3170 962
rect 3446 958 3450 962
rect 3470 958 3474 962
rect 4206 958 4210 962
rect 4758 958 4762 962
rect 4926 958 4930 962
rect 5150 958 5154 962
rect 5214 958 5218 962
rect 270 948 274 952
rect 478 948 482 952
rect 670 948 674 952
rect 814 948 818 952
rect 910 948 914 952
rect 998 948 1002 952
rect 1118 948 1122 952
rect 1134 948 1138 952
rect 1166 948 1170 952
rect 1174 948 1178 952
rect 1302 948 1306 952
rect 1414 948 1418 952
rect 1662 948 1666 952
rect 1670 948 1674 952
rect 1678 948 1682 952
rect 2134 948 2138 952
rect 2262 948 2266 952
rect 2302 948 2306 952
rect 2806 948 2810 952
rect 2958 948 2962 952
rect 3118 948 3122 952
rect 3438 948 3442 952
rect 3798 948 3802 952
rect 3974 948 3978 952
rect 4078 948 4082 952
rect 4470 948 4474 952
rect 4510 948 4514 952
rect 4622 948 4626 952
rect 4934 948 4938 952
rect 5214 948 5218 952
rect 118 938 122 942
rect 686 938 690 942
rect 1214 938 1218 942
rect 2022 938 2026 942
rect 2070 938 2074 942
rect 2422 938 2426 942
rect 2710 938 2714 942
rect 2774 938 2778 942
rect 3710 938 3714 942
rect 3726 938 3730 942
rect 4398 938 4402 942
rect 4478 938 4482 942
rect 4486 938 4490 942
rect 4894 938 4898 942
rect 478 928 482 932
rect 1086 928 1090 932
rect 1110 928 1114 932
rect 1966 928 1970 932
rect 2070 928 2074 932
rect 2406 928 2410 932
rect 2998 928 3002 932
rect 3142 928 3146 932
rect 4614 928 4618 932
rect 4982 928 4986 932
rect 182 918 186 922
rect 1334 918 1338 922
rect 1950 918 1954 922
rect 2022 918 2026 922
rect 2054 918 2058 922
rect 2318 918 2322 922
rect 2854 918 2858 922
rect 3190 918 3194 922
rect 3910 918 3914 922
rect 4318 918 4322 922
rect 4742 918 4746 922
rect 4878 918 4882 922
rect 5182 918 5186 922
rect 5254 918 5258 922
rect 894 908 898 912
rect 1118 908 1122 912
rect 1702 908 1706 912
rect 1830 908 1834 912
rect 2126 908 2130 912
rect 2174 908 2178 912
rect 3958 908 3962 912
rect 4198 908 4202 912
rect 4342 908 4346 912
rect 4814 908 4818 912
rect 5254 908 5258 912
rect 850 903 854 907
rect 858 903 861 907
rect 861 903 862 907
rect 1874 903 1878 907
rect 1882 903 1885 907
rect 1885 903 1886 907
rect 158 898 162 902
rect 830 898 834 902
rect 934 898 938 902
rect 1014 898 1018 902
rect 1390 898 1394 902
rect 1534 898 1538 902
rect 2890 903 2894 907
rect 2898 903 2901 907
rect 2901 903 2902 907
rect 3922 903 3926 907
rect 3930 903 3933 907
rect 3933 903 3934 907
rect 4938 903 4942 907
rect 4946 903 4949 907
rect 4949 903 4950 907
rect 2326 898 2330 902
rect 3766 898 3770 902
rect 4094 898 4098 902
rect 4534 898 4538 902
rect 5238 898 5242 902
rect 494 888 498 892
rect 1910 888 1914 892
rect 2174 888 2178 892
rect 2254 888 2258 892
rect 3070 888 3074 892
rect 3822 888 3826 892
rect 3902 888 3906 892
rect 4102 888 4106 892
rect 166 878 170 882
rect 1054 878 1058 882
rect 1702 878 1706 882
rect 2150 878 2154 882
rect 2214 878 2218 882
rect 2494 878 2498 882
rect 2518 878 2522 882
rect 3038 878 3042 882
rect 3094 878 3098 882
rect 3182 878 3186 882
rect 3358 878 3362 882
rect 4254 878 4258 882
rect 4598 878 4602 882
rect 4678 878 4682 882
rect 166 868 170 872
rect 886 868 890 872
rect 942 868 946 872
rect 1470 868 1474 872
rect 1686 868 1690 872
rect 1694 868 1698 872
rect 1718 868 1722 872
rect 2246 868 2250 872
rect 2646 868 2650 872
rect 3078 868 3082 872
rect 3366 868 3370 872
rect 3422 868 3426 872
rect 3494 868 3498 872
rect 3670 868 3674 872
rect 3798 868 3802 872
rect 3806 868 3810 872
rect 4054 868 4058 872
rect 4494 868 4498 872
rect 4982 868 4986 872
rect 5182 868 5186 872
rect 462 858 466 862
rect 486 858 490 862
rect 502 858 506 862
rect 574 858 578 862
rect 614 858 618 862
rect 2158 858 2162 862
rect 2374 858 2378 862
rect 2414 858 2418 862
rect 2606 858 2610 862
rect 2974 858 2978 862
rect 2990 858 2994 862
rect 3062 858 3066 862
rect 3086 858 3090 862
rect 3654 858 3658 862
rect 3718 858 3722 862
rect 3734 858 3738 862
rect 3870 858 3874 862
rect 3966 858 3970 862
rect 3990 858 3994 862
rect 4238 858 4242 862
rect 4390 858 4394 862
rect 4990 858 4994 862
rect 174 848 178 852
rect 382 848 386 852
rect 686 848 690 852
rect 806 848 810 852
rect 918 848 922 852
rect 1230 848 1234 852
rect 1710 848 1714 852
rect 1846 848 1850 852
rect 2462 848 2466 852
rect 2638 848 2642 852
rect 2822 848 2826 852
rect 3950 848 3954 852
rect 4094 848 4098 852
rect 4270 848 4274 852
rect 4590 848 4594 852
rect 5094 848 5098 852
rect 1102 838 1106 842
rect 1742 838 1746 842
rect 2486 838 2490 842
rect 2926 838 2930 842
rect 2990 838 2994 842
rect 3046 838 3050 842
rect 4510 838 4514 842
rect 4894 838 4898 842
rect 5030 838 5034 842
rect 718 828 722 832
rect 1310 828 1314 832
rect 1718 828 1722 832
rect 2710 828 2714 832
rect 4446 828 4450 832
rect 4470 828 4474 832
rect 246 818 250 822
rect 2758 818 2762 822
rect 3078 818 3082 822
rect 4462 818 4466 822
rect 4894 818 4898 822
rect 5038 818 5042 822
rect 5262 818 5266 822
rect 358 808 362 812
rect 1182 808 1186 812
rect 1246 808 1250 812
rect 1614 808 1618 812
rect 2062 808 2066 812
rect 2422 808 2426 812
rect 3030 808 3034 812
rect 3550 808 3554 812
rect 3886 808 3890 812
rect 4174 808 4178 812
rect 4726 808 4730 812
rect 5086 808 5090 812
rect 330 803 334 807
rect 338 803 341 807
rect 341 803 342 807
rect 1354 803 1358 807
rect 1362 803 1365 807
rect 1365 803 1366 807
rect 2386 803 2390 807
rect 2394 803 2397 807
rect 2397 803 2398 807
rect 3402 803 3406 807
rect 3410 803 3413 807
rect 3413 803 3414 807
rect 4426 803 4430 807
rect 4434 803 4437 807
rect 4437 803 4438 807
rect 774 798 778 802
rect 1062 798 1066 802
rect 1590 798 1594 802
rect 2030 798 2034 802
rect 2926 798 2930 802
rect 2998 798 3002 802
rect 4150 798 4154 802
rect 4166 798 4170 802
rect 4494 798 4498 802
rect 4502 798 4506 802
rect 5102 798 5106 802
rect 126 788 130 792
rect 1206 788 1210 792
rect 1374 788 1378 792
rect 1646 788 1650 792
rect 1742 788 1746 792
rect 2086 788 2090 792
rect 3302 788 3306 792
rect 3566 788 3570 792
rect 4350 788 4354 792
rect 5126 788 5130 792
rect 174 778 178 782
rect 822 778 826 782
rect 2454 778 2458 782
rect 4070 768 4074 772
rect 4150 768 4154 772
rect 5086 768 5090 772
rect 5262 768 5266 772
rect 310 758 314 762
rect 430 758 434 762
rect 718 758 722 762
rect 1118 758 1122 762
rect 2238 758 2242 762
rect 2310 758 2314 762
rect 2318 758 2322 762
rect 2350 758 2354 762
rect 2918 758 2922 762
rect 3022 758 3026 762
rect 3134 758 3138 762
rect 3502 758 3506 762
rect 4030 758 4034 762
rect 4150 758 4154 762
rect 4814 758 4818 762
rect 5006 758 5010 762
rect 5118 758 5122 762
rect 30 748 34 752
rect 254 748 258 752
rect 766 748 770 752
rect 830 748 834 752
rect 998 748 1002 752
rect 14 738 18 742
rect 1190 748 1194 752
rect 1222 748 1226 752
rect 2990 748 2994 752
rect 3038 748 3042 752
rect 3566 748 3570 752
rect 3718 748 3722 752
rect 3814 748 3818 752
rect 3982 748 3986 752
rect 4014 748 4018 752
rect 4606 748 4610 752
rect 4766 748 4770 752
rect 4870 748 4874 752
rect 4966 748 4970 752
rect 5054 748 5058 752
rect 5102 748 5106 752
rect 414 738 418 742
rect 470 738 474 742
rect 574 738 578 742
rect 774 738 778 742
rect 982 738 986 742
rect 1006 738 1010 742
rect 1782 738 1786 742
rect 1862 738 1866 742
rect 2070 738 2074 742
rect 2150 738 2154 742
rect 2286 738 2290 742
rect 2486 738 2490 742
rect 2622 738 2626 742
rect 3054 738 3058 742
rect 3238 738 3242 742
rect 3910 738 3914 742
rect 4734 738 4738 742
rect 4974 738 4978 742
rect 4990 738 4994 742
rect 5014 738 5018 742
rect 5070 738 5074 742
rect 118 728 122 732
rect 302 728 306 732
rect 942 728 946 732
rect 1214 728 1218 732
rect 1894 728 1898 732
rect 2830 728 2834 732
rect 2862 728 2866 732
rect 2990 728 2994 732
rect 3806 728 3810 732
rect 4086 728 4090 732
rect 4222 728 4226 732
rect 4446 728 4450 732
rect 5046 728 5050 732
rect 5182 728 5186 732
rect 5270 728 5274 732
rect 718 718 722 722
rect 1534 718 1538 722
rect 2718 718 2722 722
rect 2974 718 2978 722
rect 3014 718 3018 722
rect 3038 718 3042 722
rect 3814 718 3818 722
rect 4326 718 4330 722
rect 4414 718 4418 722
rect 4454 718 4458 722
rect 318 708 322 712
rect 350 708 354 712
rect 702 708 706 712
rect 1526 708 1530 712
rect 1782 708 1786 712
rect 1798 708 1802 712
rect 1862 708 1866 712
rect 2246 708 2250 712
rect 3774 708 3778 712
rect 850 703 854 707
rect 858 703 861 707
rect 861 703 862 707
rect 1874 703 1878 707
rect 1882 703 1885 707
rect 1885 703 1886 707
rect 2890 703 2894 707
rect 2898 703 2901 707
rect 2901 703 2902 707
rect 3922 703 3926 707
rect 3930 703 3933 707
rect 3933 703 3934 707
rect 446 698 450 702
rect 1270 698 1274 702
rect 1966 698 1970 702
rect 2182 698 2186 702
rect 2862 698 2866 702
rect 3102 698 3106 702
rect 3318 698 3322 702
rect 3326 698 3330 702
rect 3638 698 3642 702
rect 4174 698 4178 702
rect 4398 698 4402 702
rect 4938 703 4942 707
rect 4946 703 4949 707
rect 4949 703 4950 707
rect 438 688 442 692
rect 470 688 474 692
rect 2982 688 2986 692
rect 3294 688 3298 692
rect 3710 688 3714 692
rect 4054 688 4058 692
rect 4614 688 4618 692
rect 4726 688 4730 692
rect 4886 688 4890 692
rect 5006 688 5010 692
rect 358 678 362 682
rect 1198 678 1202 682
rect 1206 678 1210 682
rect 1318 678 1322 682
rect 1374 678 1378 682
rect 2094 678 2098 682
rect 2710 678 2714 682
rect 3046 678 3050 682
rect 3166 678 3170 682
rect 3454 678 3458 682
rect 3494 678 3498 682
rect 3838 678 3842 682
rect 4062 678 4066 682
rect 4190 678 4194 682
rect 4526 678 4530 682
rect 4574 678 4578 682
rect 4606 678 4610 682
rect 4678 678 4682 682
rect 4934 678 4938 682
rect 5046 678 5050 682
rect 214 668 218 672
rect 870 668 874 672
rect 998 668 1002 672
rect 1110 668 1114 672
rect 1798 668 1802 672
rect 2246 668 2250 672
rect 2334 668 2338 672
rect 2406 668 2410 672
rect 2694 668 2698 672
rect 2750 668 2754 672
rect 3094 668 3098 672
rect 3126 668 3130 672
rect 3430 668 3434 672
rect 3814 668 3818 672
rect 3982 668 3986 672
rect 4014 668 4018 672
rect 4126 668 4130 672
rect 4310 668 4314 672
rect 4910 668 4914 672
rect 5062 668 5066 672
rect 5070 668 5074 672
rect 54 658 58 662
rect 118 658 122 662
rect 302 658 306 662
rect 406 658 410 662
rect 422 658 426 662
rect 702 658 706 662
rect 1006 658 1010 662
rect 1190 658 1194 662
rect 1382 658 1386 662
rect 1446 658 1450 662
rect 1494 658 1498 662
rect 1814 658 1818 662
rect 2070 658 2074 662
rect 2214 658 2218 662
rect 2246 658 2250 662
rect 2702 658 2706 662
rect 2726 658 2730 662
rect 3526 658 3530 662
rect 3542 658 3546 662
rect 3998 658 4002 662
rect 4038 658 4042 662
rect 4206 658 4210 662
rect 4302 658 4306 662
rect 4654 658 4658 662
rect 4710 658 4714 662
rect 4894 658 4898 662
rect 5046 658 5050 662
rect 350 648 354 652
rect 750 648 754 652
rect 1246 648 1250 652
rect 1806 648 1810 652
rect 2334 648 2338 652
rect 2750 648 2754 652
rect 2870 648 2874 652
rect 3438 648 3442 652
rect 4078 648 4082 652
rect 5030 648 5034 652
rect 478 638 482 642
rect 758 638 762 642
rect 1278 638 1282 642
rect 2014 638 2018 642
rect 3166 638 3170 642
rect 4606 638 4610 642
rect 174 628 178 632
rect 990 628 994 632
rect 1678 628 1682 632
rect 2358 628 2362 632
rect 2742 628 2746 632
rect 3630 628 3634 632
rect 3942 628 3946 632
rect 4446 628 4450 632
rect 4974 628 4978 632
rect 670 618 674 622
rect 2654 618 2658 622
rect 2910 618 2914 622
rect 3542 618 3546 622
rect 4494 618 4498 622
rect 4710 618 4714 622
rect 5078 618 5082 622
rect 190 608 194 612
rect 758 608 762 612
rect 1334 608 1338 612
rect 2030 608 2034 612
rect 3422 608 3426 612
rect 4870 608 4874 612
rect 330 603 334 607
rect 338 603 341 607
rect 341 603 342 607
rect 1354 603 1358 607
rect 1362 603 1365 607
rect 1365 603 1366 607
rect 2386 603 2390 607
rect 2394 603 2397 607
rect 2397 603 2398 607
rect 3402 603 3406 607
rect 3410 603 3413 607
rect 3413 603 3414 607
rect 4426 603 4430 607
rect 4434 603 4437 607
rect 4437 603 4438 607
rect 318 598 322 602
rect 1766 598 1770 602
rect 2918 598 2922 602
rect 3686 598 3690 602
rect 3558 588 3562 592
rect 3806 588 3810 592
rect 4134 588 4138 592
rect 2198 578 2202 582
rect 3206 578 3210 582
rect 3702 578 3706 582
rect 3942 578 3946 582
rect 3974 578 3978 582
rect 4662 578 4666 582
rect 4766 578 4770 582
rect 1014 568 1018 572
rect 1238 568 1242 572
rect 1342 568 1346 572
rect 2486 568 2490 572
rect 3910 568 3914 572
rect 4918 568 4922 572
rect 5134 568 5138 572
rect 534 558 538 562
rect 678 558 682 562
rect 1022 558 1026 562
rect 1382 558 1386 562
rect 1614 558 1618 562
rect 2038 558 2042 562
rect 2230 558 2234 562
rect 2478 558 2482 562
rect 2574 558 2578 562
rect 2662 558 2666 562
rect 3038 558 3042 562
rect 3126 558 3130 562
rect 3798 558 3802 562
rect 3902 558 3906 562
rect 4894 558 4898 562
rect 342 548 346 552
rect 350 548 354 552
rect 494 548 498 552
rect 782 548 786 552
rect 1278 548 1282 552
rect 1294 548 1298 552
rect 1422 548 1426 552
rect 1678 548 1682 552
rect 1790 548 1794 552
rect 1974 548 1978 552
rect 2374 548 2378 552
rect 318 538 322 542
rect 814 538 818 542
rect 950 538 954 542
rect 1262 538 1266 542
rect 1286 538 1290 542
rect 2886 548 2890 552
rect 3198 548 3202 552
rect 3502 548 3506 552
rect 3638 548 3642 552
rect 3694 548 3698 552
rect 3774 548 3778 552
rect 4014 548 4018 552
rect 4150 548 4154 552
rect 4214 548 4218 552
rect 4574 548 4578 552
rect 4590 548 4594 552
rect 4734 548 4738 552
rect 1798 538 1802 542
rect 2054 538 2058 542
rect 2158 538 2162 542
rect 2174 538 2178 542
rect 3742 538 3746 542
rect 4342 538 4346 542
rect 1702 528 1706 532
rect 3086 528 3090 532
rect 3222 528 3226 532
rect 3894 528 3898 532
rect 4030 528 4034 532
rect 5174 528 5178 532
rect 5294 528 5298 532
rect 2118 518 2122 522
rect 2166 518 2170 522
rect 2646 518 2650 522
rect 3830 518 3834 522
rect 4550 518 4554 522
rect 302 508 306 512
rect 1910 508 1914 512
rect 2022 508 2026 512
rect 2630 508 2634 512
rect 3070 508 3074 512
rect 4094 508 4098 512
rect 4406 508 4410 512
rect 4758 508 4762 512
rect 5110 508 5114 512
rect 850 503 854 507
rect 858 503 861 507
rect 861 503 862 507
rect 1874 503 1878 507
rect 1882 503 1885 507
rect 1885 503 1886 507
rect 2890 503 2894 507
rect 2898 503 2901 507
rect 2901 503 2902 507
rect 3922 503 3926 507
rect 3930 503 3933 507
rect 3933 503 3934 507
rect 4938 503 4942 507
rect 4946 503 4949 507
rect 4949 503 4950 507
rect 782 498 786 502
rect 1326 498 1330 502
rect 1934 498 1938 502
rect 2446 498 2450 502
rect 2726 498 2730 502
rect 2734 498 2738 502
rect 3574 498 3578 502
rect 4166 498 4170 502
rect 4542 498 4546 502
rect 5094 498 5098 502
rect 1438 488 1442 492
rect 1566 488 1570 492
rect 1726 488 1730 492
rect 1774 488 1778 492
rect 2926 488 2930 492
rect 3030 488 3034 492
rect 3294 488 3298 492
rect 3390 488 3394 492
rect 4134 488 4138 492
rect 4150 488 4154 492
rect 4526 488 4530 492
rect 5038 488 5042 492
rect 5102 488 5106 492
rect 5182 488 5186 492
rect 486 478 490 482
rect 806 478 810 482
rect 822 478 826 482
rect 1766 478 1770 482
rect 1902 478 1906 482
rect 2678 478 2682 482
rect 3734 478 3738 482
rect 4046 478 4050 482
rect 4534 478 4538 482
rect 4894 478 4898 482
rect 4934 478 4938 482
rect 5206 478 5210 482
rect 5270 478 5274 482
rect 166 468 170 472
rect 550 468 554 472
rect 670 468 674 472
rect 1270 468 1274 472
rect 2062 468 2066 472
rect 2334 468 2338 472
rect 3078 468 3082 472
rect 294 458 298 462
rect 486 458 490 462
rect 774 458 778 462
rect 1302 458 1306 462
rect 1694 458 1698 462
rect 2782 458 2786 462
rect 2926 458 2930 462
rect 3006 458 3010 462
rect 3550 468 3554 472
rect 3702 468 3706 472
rect 3710 468 3714 472
rect 3902 468 3906 472
rect 3910 468 3914 472
rect 3982 468 3986 472
rect 4206 468 4210 472
rect 4406 468 4410 472
rect 4990 468 4994 472
rect 3478 458 3482 462
rect 3542 458 3546 462
rect 3566 458 3570 462
rect 3822 458 3826 462
rect 4118 458 4122 462
rect 4390 458 4394 462
rect 4838 458 4842 462
rect 5014 458 5018 462
rect 5038 458 5042 462
rect 5054 458 5058 462
rect 5182 458 5186 462
rect 5230 458 5234 462
rect 182 448 186 452
rect 806 448 810 452
rect 1670 448 1674 452
rect 1774 448 1778 452
rect 14 438 18 442
rect 390 438 394 442
rect 1302 438 1306 442
rect 1854 438 1858 442
rect 2526 448 2530 452
rect 2870 448 2874 452
rect 3182 448 3186 452
rect 3526 448 3530 452
rect 3542 448 3546 452
rect 3686 448 3690 452
rect 3782 448 3786 452
rect 4774 448 4778 452
rect 4966 448 4970 452
rect 3014 438 3018 442
rect 3110 438 3114 442
rect 4166 438 4170 442
rect 174 428 178 432
rect 1534 428 1538 432
rect 1942 428 1946 432
rect 2518 428 2522 432
rect 766 418 770 422
rect 982 418 986 422
rect 1782 418 1786 422
rect 3278 418 3282 422
rect 4030 418 4034 422
rect 4598 418 4602 422
rect 4686 418 4690 422
rect 4710 418 4714 422
rect 1214 408 1218 412
rect 1806 408 1810 412
rect 2110 408 2114 412
rect 3526 408 3530 412
rect 3774 408 3778 412
rect 4102 408 4106 412
rect 330 403 334 407
rect 338 403 341 407
rect 341 403 342 407
rect 1354 403 1358 407
rect 1362 403 1365 407
rect 1365 403 1366 407
rect 2386 403 2390 407
rect 2394 403 2397 407
rect 2397 403 2398 407
rect 3402 403 3406 407
rect 3410 403 3413 407
rect 3413 403 3414 407
rect 4426 403 4430 407
rect 4434 403 4437 407
rect 4437 403 4438 407
rect 686 398 690 402
rect 1246 398 1250 402
rect 2718 398 2722 402
rect 3438 398 3442 402
rect 4038 398 4042 402
rect 4598 398 4602 402
rect 5286 398 5290 402
rect 550 388 554 392
rect 1382 388 1386 392
rect 1918 388 1922 392
rect 2702 388 2706 392
rect 3262 388 3266 392
rect 3606 388 3610 392
rect 5166 388 5170 392
rect 1374 378 1378 382
rect 1782 378 1786 382
rect 2094 378 2098 382
rect 2150 378 2154 382
rect 2654 378 2658 382
rect 3046 378 3050 382
rect 3342 378 3346 382
rect 4574 378 4578 382
rect 5198 378 5202 382
rect 758 368 762 372
rect 1278 368 1282 372
rect 2126 368 2130 372
rect 2702 368 2706 372
rect 3494 368 3498 372
rect 5254 368 5258 372
rect 206 358 210 362
rect 254 358 258 362
rect 1014 358 1018 362
rect 1542 358 1546 362
rect 2014 358 2018 362
rect 2246 358 2250 362
rect 2414 358 2418 362
rect 3158 358 3162 362
rect 3510 358 3514 362
rect 3702 358 3706 362
rect 3806 358 3810 362
rect 4126 358 4130 362
rect 4582 358 4586 362
rect 4910 358 4914 362
rect 5190 358 5194 362
rect 14 348 18 352
rect 326 348 330 352
rect 1118 348 1122 352
rect 1254 348 1258 352
rect 1590 348 1594 352
rect 1982 348 1986 352
rect 2038 348 2042 352
rect 2094 348 2098 352
rect 2590 348 2594 352
rect 3190 348 3194 352
rect 3550 348 3554 352
rect 3622 348 3626 352
rect 3838 348 3842 352
rect 4030 348 4034 352
rect 4198 348 4202 352
rect 4686 348 4690 352
rect 4710 348 4714 352
rect 5150 348 5154 352
rect 1310 338 1314 342
rect 1766 338 1770 342
rect 1798 338 1802 342
rect 2062 338 2066 342
rect 2134 338 2138 342
rect 2398 338 2402 342
rect 3654 338 3658 342
rect 4174 338 4178 342
rect 4222 338 4226 342
rect 4694 338 4698 342
rect 4974 338 4978 342
rect 5006 338 5010 342
rect 5262 338 5266 342
rect 310 328 314 332
rect 1014 328 1018 332
rect 1566 328 1570 332
rect 2286 328 2290 332
rect 2654 328 2658 332
rect 4486 328 4490 332
rect 5158 328 5162 332
rect 262 318 266 322
rect 1334 318 1338 322
rect 1582 318 1586 322
rect 4926 318 4930 322
rect 4958 318 4962 322
rect 5278 318 5282 322
rect 1742 308 1746 312
rect 2358 308 2362 312
rect 5214 308 5218 312
rect 5238 308 5242 312
rect 850 303 854 307
rect 858 303 861 307
rect 861 303 862 307
rect 1874 303 1878 307
rect 1882 303 1885 307
rect 1885 303 1886 307
rect 2890 303 2894 307
rect 2898 303 2901 307
rect 2901 303 2902 307
rect 3922 303 3926 307
rect 3930 303 3933 307
rect 3933 303 3934 307
rect 4938 303 4942 307
rect 4946 303 4949 307
rect 4949 303 4950 307
rect 286 298 290 302
rect 798 298 802 302
rect 198 288 202 292
rect 958 288 962 292
rect 1526 288 1530 292
rect 2246 288 2250 292
rect 2934 288 2938 292
rect 4998 288 5002 292
rect 5094 288 5098 292
rect 5206 288 5210 292
rect 5246 288 5250 292
rect 350 278 354 282
rect 638 278 642 282
rect 806 278 810 282
rect 878 278 882 282
rect 1958 268 1962 272
rect 3486 278 3490 282
rect 3662 278 3666 282
rect 3710 278 3714 282
rect 4534 278 4538 282
rect 4926 278 4930 282
rect 5214 278 5218 282
rect 5286 278 5290 282
rect 2678 268 2682 272
rect 2734 268 2738 272
rect 2918 268 2922 272
rect 3526 268 3530 272
rect 3566 268 3570 272
rect 3998 268 4002 272
rect 4214 268 4218 272
rect 4582 268 4586 272
rect 4902 268 4906 272
rect 5302 268 5306 272
rect 142 258 146 262
rect 254 258 258 262
rect 686 258 690 262
rect 2150 258 2154 262
rect 2630 258 2634 262
rect 2718 258 2722 262
rect 2726 258 2730 262
rect 3182 258 3186 262
rect 3742 258 3746 262
rect 4198 258 4202 262
rect 4998 258 5002 262
rect 5022 258 5026 262
rect 5062 258 5066 262
rect 5222 258 5226 262
rect 422 248 426 252
rect 1286 248 1290 252
rect 1782 248 1786 252
rect 2334 248 2338 252
rect 1670 238 1674 242
rect 2062 238 2066 242
rect 3022 238 3026 242
rect 3574 248 3578 252
rect 4774 248 4778 252
rect 3382 238 3386 242
rect 2126 228 2130 232
rect 4526 228 4530 232
rect 4550 228 4554 232
rect 5062 228 5066 232
rect 1038 218 1042 222
rect 1566 218 1570 222
rect 1678 218 1682 222
rect 3646 218 3650 222
rect 4414 218 4418 222
rect 4830 218 4834 222
rect 3654 208 3658 212
rect 3894 208 3898 212
rect 330 203 334 207
rect 338 203 341 207
rect 341 203 342 207
rect 1354 203 1358 207
rect 1362 203 1365 207
rect 1365 203 1366 207
rect 2386 203 2390 207
rect 2394 203 2397 207
rect 2397 203 2398 207
rect 3402 203 3406 207
rect 3410 203 3413 207
rect 3413 203 3414 207
rect 4426 203 4430 207
rect 4434 203 4437 207
rect 4437 203 4438 207
rect 2630 198 2634 202
rect 4406 198 4410 202
rect 2662 188 2666 192
rect 3166 188 3170 192
rect 3494 188 3498 192
rect 5078 188 5082 192
rect 1582 178 1586 182
rect 1774 178 1778 182
rect 2358 178 2362 182
rect 4686 178 4690 182
rect 4574 168 4578 172
rect 4702 168 4706 172
rect 5230 168 5234 172
rect 2038 158 2042 162
rect 4102 158 4106 162
rect 4118 158 4122 162
rect 4982 158 4986 162
rect 14 148 18 152
rect 302 148 306 152
rect 1238 148 1242 152
rect 1774 148 1778 152
rect 1846 148 1850 152
rect 2150 148 2154 152
rect 2622 148 2626 152
rect 2662 148 2666 152
rect 2982 148 2986 152
rect 3086 148 3090 152
rect 3094 148 3098 152
rect 3110 148 3114 152
rect 3494 148 3498 152
rect 4214 148 4218 152
rect 4750 148 4754 152
rect 5246 148 5250 152
rect 5270 148 5274 152
rect 390 138 394 142
rect 2934 138 2938 142
rect 3462 138 3466 142
rect 3646 138 3650 142
rect 3982 138 3986 142
rect 4070 138 4074 142
rect 4310 138 4314 142
rect 2086 128 2090 132
rect 2694 128 2698 132
rect 3534 128 3538 132
rect 3638 128 3642 132
rect 4870 128 4874 132
rect 4886 128 4890 132
rect 5262 128 5266 132
rect 838 118 842 122
rect 3574 118 3578 122
rect 1894 108 1898 112
rect 3462 108 3466 112
rect 3942 108 3946 112
rect 4246 108 4250 112
rect 4430 108 4434 112
rect 4438 108 4442 112
rect 4798 108 4802 112
rect 850 103 854 107
rect 858 103 861 107
rect 861 103 862 107
rect 1874 103 1878 107
rect 1882 103 1885 107
rect 1885 103 1886 107
rect 2890 103 2894 107
rect 2898 103 2901 107
rect 2901 103 2902 107
rect 3922 103 3926 107
rect 3930 103 3933 107
rect 3933 103 3934 107
rect 4938 103 4942 107
rect 4946 103 4949 107
rect 4949 103 4950 107
rect 2086 98 2090 102
rect 2646 98 2650 102
rect 2910 98 2914 102
rect 446 88 450 92
rect 1798 88 1802 92
rect 1894 88 1898 92
rect 1918 88 1922 92
rect 3382 88 3386 92
rect 3390 88 3394 92
rect 3470 88 3474 92
rect 3494 88 3498 92
rect 3574 88 3578 92
rect 3710 88 3714 92
rect 3942 88 3946 92
rect 4126 88 4130 92
rect 4374 88 4378 92
rect 4830 88 4834 92
rect 4878 88 4882 92
rect 1374 78 1378 82
rect 1702 78 1706 82
rect 3430 78 3434 82
rect 3502 78 3506 82
rect 4438 78 4442 82
rect 4446 78 4450 82
rect 4526 78 4530 82
rect 4822 78 4826 82
rect 4918 78 4922 82
rect 5030 78 5034 82
rect 2030 68 2034 72
rect 3438 68 3442 72
rect 3734 68 3738 72
rect 3918 68 3922 72
rect 4406 68 4410 72
rect 5142 68 5146 72
rect 5230 68 5234 72
rect 638 58 642 62
rect 1918 58 1922 62
rect 2542 58 2546 62
rect 2726 58 2730 62
rect 2822 58 2826 62
rect 2934 58 2938 62
rect 2958 58 2962 62
rect 3534 58 3538 62
rect 3566 58 3570 62
rect 3606 58 3610 62
rect 4150 58 4154 62
rect 4254 58 4258 62
rect 4726 58 4730 62
rect 4958 58 4962 62
rect 5126 58 5130 62
rect 5166 58 5170 62
rect 4766 48 4770 52
rect 5182 48 5186 52
rect 4982 38 4986 42
rect 2222 8 2226 12
rect 4534 8 4538 12
rect 330 3 334 7
rect 338 3 341 7
rect 341 3 342 7
rect 1354 3 1358 7
rect 1362 3 1365 7
rect 1365 3 1366 7
rect 2386 3 2390 7
rect 2394 3 2397 7
rect 2397 3 2398 7
rect 3402 3 3406 7
rect 3410 3 3413 7
rect 3413 3 3414 7
rect 4426 3 4430 7
rect 4434 3 4437 7
rect 4437 3 4438 7
<< metal4 >>
rect 848 5103 850 5107
rect 854 5103 857 5107
rect 862 5103 864 5107
rect 1872 5103 1874 5107
rect 1878 5103 1881 5107
rect 1886 5103 1888 5107
rect 2888 5103 2890 5107
rect 2894 5103 2897 5107
rect 2902 5103 2904 5107
rect 3920 5103 3922 5107
rect 3926 5103 3929 5107
rect 3934 5103 3936 5107
rect 4936 5103 4938 5107
rect 4942 5103 4945 5107
rect 4950 5103 4952 5107
rect 310 5098 318 5101
rect 1658 5098 1665 5101
rect 310 5072 313 5098
rect 170 5058 174 5061
rect 202 5058 206 5061
rect 328 5003 330 5007
rect 334 5003 337 5007
rect 342 5003 344 5007
rect 186 4948 190 4951
rect 182 4892 185 4948
rect 202 4928 206 4931
rect 118 4868 126 4871
rect 38 4712 41 4858
rect 46 4542 49 4748
rect 46 4382 49 4538
rect 86 4442 89 4758
rect 118 4722 121 4868
rect 170 4848 177 4851
rect 126 4672 129 4688
rect 94 4341 97 4598
rect 90 4338 97 4341
rect 22 4171 25 4298
rect 102 4261 105 4348
rect 98 4258 105 4261
rect 18 4168 25 4171
rect 110 4042 113 4458
rect 134 4352 137 4578
rect 142 4482 145 4738
rect 174 4542 177 4848
rect 214 4842 217 4948
rect 246 4852 249 4948
rect 246 4822 249 4848
rect 286 4762 289 4968
rect 366 4942 369 5028
rect 374 4922 377 4958
rect 328 4803 330 4807
rect 334 4803 337 4807
rect 342 4803 344 4807
rect 414 4752 417 4808
rect 422 4752 425 4958
rect 430 4762 433 4778
rect 438 4772 441 4968
rect 462 4912 465 5058
rect 474 4958 478 4961
rect 486 4932 489 4958
rect 546 4878 550 4881
rect 566 4842 569 5058
rect 486 4778 494 4781
rect 214 4642 217 4738
rect 142 4442 145 4478
rect 38 3771 41 3968
rect 38 3768 46 3771
rect 78 3752 81 3978
rect 122 3878 129 3881
rect 106 3838 110 3841
rect 86 3752 89 3768
rect 94 3752 97 3838
rect 50 3748 54 3751
rect 102 3742 105 3818
rect 30 1822 33 3458
rect 102 3282 105 3738
rect 118 3672 121 3858
rect 126 3832 129 3878
rect 126 3812 129 3828
rect 134 3772 137 4348
rect 214 4282 217 4618
rect 202 4278 206 4281
rect 222 4262 225 4648
rect 278 4392 281 4658
rect 326 4652 329 4678
rect 342 4652 345 4668
rect 328 4603 330 4607
rect 334 4603 337 4607
rect 342 4603 344 4607
rect 328 4403 330 4407
rect 334 4403 337 4407
rect 342 4403 344 4407
rect 254 4272 257 4318
rect 142 3992 145 4188
rect 158 4052 161 4108
rect 254 4102 257 4268
rect 142 3962 145 3988
rect 198 3932 201 4088
rect 278 4052 281 4388
rect 198 3912 201 3928
rect 214 3848 222 3851
rect 214 3842 217 3848
rect 310 3822 313 3958
rect 318 3812 321 4328
rect 358 4252 361 4618
rect 414 4572 417 4638
rect 370 4538 374 4541
rect 390 4351 393 4478
rect 402 4428 409 4431
rect 386 4348 393 4351
rect 328 4203 330 4207
rect 334 4203 337 4207
rect 342 4203 344 4207
rect 350 4192 353 4228
rect 358 4082 361 4248
rect 366 4122 369 4288
rect 398 4242 401 4368
rect 406 4252 409 4428
rect 414 4302 417 4568
rect 450 4558 454 4561
rect 442 4538 446 4541
rect 454 4352 457 4558
rect 462 4342 465 4768
rect 486 4642 489 4778
rect 470 4522 473 4558
rect 494 4471 497 4548
rect 494 4468 502 4471
rect 486 4332 489 4338
rect 328 4003 330 4007
rect 334 4003 337 4007
rect 342 4003 344 4007
rect 350 3972 353 3998
rect 382 3942 385 4178
rect 414 4162 417 4298
rect 470 4222 473 4278
rect 530 4178 534 4181
rect 414 3992 417 4058
rect 382 3862 385 3938
rect 328 3803 330 3807
rect 334 3803 337 3807
rect 342 3803 344 3807
rect 134 3342 137 3728
rect 206 3682 209 3758
rect 150 3562 153 3568
rect 42 2858 46 2861
rect 86 2662 89 2668
rect 110 2662 113 2868
rect 122 2668 126 2671
rect 110 2132 113 2548
rect 142 2442 145 2858
rect 158 2152 161 3058
rect 198 2862 201 3058
rect 206 2882 209 3578
rect 294 3152 297 3618
rect 328 3603 330 3607
rect 334 3603 337 3607
rect 342 3603 344 3607
rect 390 3502 393 3948
rect 446 3842 449 3958
rect 466 3838 470 3841
rect 478 3822 481 4128
rect 494 4012 497 4048
rect 502 3952 505 4138
rect 510 4032 513 4158
rect 534 4122 537 4158
rect 542 4132 545 4518
rect 550 4412 553 4818
rect 606 4792 609 4918
rect 706 4878 710 4881
rect 638 4762 641 4778
rect 634 4728 638 4731
rect 582 4612 585 4618
rect 590 4612 593 4648
rect 558 4382 561 4468
rect 574 4452 577 4568
rect 598 4562 601 4618
rect 582 4432 585 4558
rect 598 4542 601 4558
rect 638 4372 641 4548
rect 662 4532 665 4768
rect 726 4702 729 4968
rect 742 4962 745 4968
rect 758 4932 761 4948
rect 774 4942 777 4948
rect 806 4942 809 5038
rect 794 4858 798 4861
rect 738 4848 742 4851
rect 734 4762 737 4768
rect 742 4732 745 4788
rect 670 4602 673 4668
rect 742 4662 745 4728
rect 694 4612 697 4618
rect 670 4491 673 4598
rect 694 4572 697 4608
rect 670 4488 678 4491
rect 694 4342 697 4568
rect 702 4342 705 4348
rect 566 4332 569 4338
rect 542 3912 545 4098
rect 550 4082 553 4118
rect 566 4092 569 4118
rect 510 3742 513 3898
rect 550 3892 553 4078
rect 558 3952 561 4078
rect 582 4072 585 4268
rect 614 4262 617 4278
rect 594 4258 598 4261
rect 622 4112 625 4258
rect 638 4252 641 4268
rect 650 4248 654 4251
rect 630 4082 633 4188
rect 678 4171 681 4328
rect 678 4168 686 4171
rect 694 4162 697 4338
rect 638 4112 641 4128
rect 566 4032 569 4058
rect 582 3982 585 4068
rect 638 4042 641 4108
rect 594 3978 598 3981
rect 574 3972 577 3978
rect 702 3852 705 4328
rect 710 4172 713 4468
rect 718 4452 721 4458
rect 718 4222 721 4448
rect 726 4412 729 4588
rect 726 4202 729 4378
rect 742 4352 745 4658
rect 774 4442 777 4648
rect 774 4292 777 4438
rect 790 4422 793 4698
rect 806 4512 809 4938
rect 838 4662 841 5058
rect 848 4903 850 4907
rect 854 4903 857 4907
rect 862 4903 864 4907
rect 870 4902 873 4928
rect 874 4858 878 4861
rect 854 4732 857 4748
rect 914 4728 918 4731
rect 848 4703 850 4707
rect 854 4703 857 4707
rect 862 4703 864 4707
rect 926 4701 929 5008
rect 934 4712 937 4918
rect 950 4872 953 5028
rect 922 4698 929 4701
rect 822 4432 825 4618
rect 848 4503 850 4507
rect 854 4503 857 4507
rect 862 4503 864 4507
rect 886 4452 889 4468
rect 798 4372 801 4398
rect 802 4348 806 4351
rect 848 4303 850 4307
rect 854 4303 857 4307
rect 862 4303 864 4307
rect 738 4268 742 4271
rect 878 4262 881 4418
rect 926 4412 929 4698
rect 950 4471 953 4698
rect 946 4468 953 4471
rect 974 4482 977 4588
rect 998 4512 1001 4758
rect 1014 4541 1017 4718
rect 1010 4538 1017 4541
rect 770 4258 777 4261
rect 786 4258 790 4261
rect 774 4252 777 4258
rect 814 4232 817 4258
rect 830 4242 833 4248
rect 886 4202 889 4348
rect 974 4262 977 4478
rect 1022 4352 1025 4868
rect 1030 4432 1033 4538
rect 1038 4532 1041 4758
rect 1046 4522 1049 4878
rect 1070 4462 1073 4478
rect 1070 4452 1073 4458
rect 1078 4372 1081 4858
rect 1134 4762 1137 5078
rect 1352 5003 1354 5007
rect 1358 5003 1361 5007
rect 1366 5003 1368 5007
rect 1458 4948 1462 4951
rect 1134 4742 1137 4758
rect 1174 4732 1177 4868
rect 1246 4748 1254 4751
rect 1102 4728 1110 4731
rect 1102 4662 1105 4728
rect 1246 4592 1249 4748
rect 1150 4552 1153 4558
rect 1022 4282 1025 4348
rect 726 4072 729 4198
rect 848 4103 850 4107
rect 854 4103 857 4107
rect 862 4103 864 4107
rect 510 3652 513 3738
rect 630 3662 633 3668
rect 462 3572 465 3588
rect 398 3452 401 3488
rect 328 3403 330 3407
rect 334 3403 337 3407
rect 342 3403 344 3407
rect 262 2852 265 2858
rect 246 2712 249 2838
rect 258 2748 262 2751
rect 214 2262 217 2698
rect 254 2542 257 2678
rect 214 1862 217 2258
rect 246 2052 249 2228
rect 238 2048 246 2051
rect 30 752 33 1818
rect 126 1312 129 1678
rect 126 1272 129 1308
rect 118 1268 126 1271
rect 118 942 121 1268
rect 14 442 17 738
rect 118 732 121 938
rect 126 792 129 1138
rect 142 1082 145 1538
rect 150 1142 153 1548
rect 158 902 161 1218
rect 166 882 169 1788
rect 174 1638 182 1641
rect 174 1442 177 1638
rect 54 662 57 718
rect 118 662 121 728
rect 166 472 169 868
rect 174 852 177 1438
rect 182 962 185 1098
rect 174 782 177 848
rect 14 352 17 438
rect 174 432 177 628
rect 182 452 185 918
rect 194 608 201 611
rect 14 152 17 348
rect 198 292 201 608
rect 206 542 209 1848
rect 214 1522 217 1528
rect 214 1502 217 1518
rect 222 1491 225 1918
rect 214 1488 225 1491
rect 230 1842 233 2008
rect 214 672 217 1488
rect 230 1472 233 1838
rect 230 1282 233 1468
rect 238 1302 241 2048
rect 262 1352 265 2588
rect 270 2552 273 2868
rect 286 2461 289 2988
rect 294 2592 297 3148
rect 282 2458 289 2461
rect 278 2262 281 2398
rect 290 2268 294 2271
rect 302 2162 305 3318
rect 406 3222 409 3558
rect 466 3528 470 3531
rect 502 3372 505 3578
rect 510 3482 513 3648
rect 562 3528 566 3531
rect 510 3422 513 3458
rect 562 3358 566 3361
rect 430 3342 433 3358
rect 590 3332 593 3528
rect 582 3328 590 3331
rect 446 3282 449 3328
rect 582 3322 585 3328
rect 470 3232 473 3258
rect 328 3203 330 3207
rect 334 3203 337 3207
rect 342 3203 344 3207
rect 328 3003 330 3007
rect 334 3003 337 3007
rect 342 3003 344 3007
rect 310 2742 313 2978
rect 328 2803 330 2807
rect 334 2803 337 2807
rect 342 2803 344 2807
rect 310 2702 313 2738
rect 328 2603 330 2607
rect 334 2603 337 2607
rect 342 2603 344 2607
rect 328 2403 330 2407
rect 334 2403 337 2407
rect 342 2403 344 2407
rect 234 1258 238 1261
rect 222 1062 225 1178
rect 222 1002 225 1058
rect 246 822 249 1338
rect 270 1162 273 1878
rect 286 1662 289 2128
rect 302 1472 305 2098
rect 310 1882 313 2278
rect 318 2251 321 2258
rect 318 2248 326 2251
rect 328 2203 330 2207
rect 334 2203 337 2207
rect 342 2203 344 2207
rect 328 2003 330 2007
rect 334 2003 337 2007
rect 342 2003 344 2007
rect 318 1822 321 1948
rect 358 1852 361 2818
rect 366 2282 369 3098
rect 394 2838 401 2841
rect 398 2672 401 2838
rect 374 2272 377 2558
rect 270 952 273 1158
rect 206 362 209 538
rect 254 362 257 748
rect 254 262 257 358
rect 262 262 265 318
rect 286 302 289 1268
rect 302 1112 305 1468
rect 310 1242 313 1648
rect 302 732 305 1098
rect 318 962 321 1808
rect 328 1803 330 1807
rect 334 1803 337 1807
rect 342 1803 344 1807
rect 328 1603 330 1607
rect 334 1603 337 1607
rect 342 1603 344 1607
rect 366 1512 369 1878
rect 374 1762 377 2028
rect 406 1962 409 3218
rect 582 3122 585 3318
rect 590 3272 593 3308
rect 594 3128 598 3131
rect 454 2892 457 2908
rect 470 2562 473 2798
rect 490 2688 494 2691
rect 338 1438 342 1441
rect 328 1403 330 1407
rect 334 1403 337 1407
rect 342 1403 344 1407
rect 328 1203 330 1207
rect 334 1203 337 1207
rect 342 1203 344 1207
rect 328 1003 330 1007
rect 334 1003 337 1007
rect 342 1003 344 1007
rect 302 662 305 728
rect 302 461 305 508
rect 298 458 305 461
rect 146 258 150 261
rect 302 152 305 458
rect 310 332 313 758
rect 318 712 321 938
rect 358 812 361 1038
rect 382 852 385 1848
rect 406 1622 409 1958
rect 390 1462 393 1618
rect 414 1562 417 1758
rect 406 1542 409 1548
rect 406 1452 409 1458
rect 394 1348 398 1351
rect 406 1262 409 1268
rect 414 1162 417 1448
rect 422 1342 425 1348
rect 430 1262 433 2428
rect 502 2351 505 2918
rect 518 2852 521 2968
rect 510 2842 513 2848
rect 526 2682 529 2868
rect 558 2862 561 3058
rect 606 2952 609 3078
rect 614 2882 617 3108
rect 598 2832 601 2878
rect 534 2672 537 2818
rect 590 2712 593 2748
rect 498 2348 505 2351
rect 518 2362 521 2668
rect 550 2652 553 2668
rect 590 2662 593 2708
rect 582 2492 585 2658
rect 530 2368 534 2371
rect 518 2342 521 2358
rect 458 2338 462 2341
rect 526 2262 529 2348
rect 446 1642 449 2108
rect 542 2082 545 2088
rect 506 2048 510 2051
rect 454 1582 457 1668
rect 454 1482 457 1578
rect 438 1268 446 1271
rect 406 1132 409 1148
rect 328 803 330 807
rect 334 803 337 807
rect 342 803 344 807
rect 350 652 353 708
rect 358 682 361 808
rect 406 662 409 1128
rect 430 762 433 1258
rect 438 1252 441 1268
rect 414 732 417 738
rect 438 692 441 1248
rect 462 862 465 1278
rect 470 1062 473 1548
rect 502 1458 510 1461
rect 470 742 473 998
rect 478 952 481 988
rect 328 603 330 607
rect 334 603 337 607
rect 342 603 344 607
rect 318 542 321 598
rect 342 552 345 558
rect 350 552 353 648
rect 328 403 330 407
rect 334 403 337 407
rect 342 403 344 407
rect 330 348 334 351
rect 350 282 353 548
rect 328 203 330 207
rect 334 203 337 207
rect 342 203 344 207
rect 390 142 393 438
rect 422 252 425 658
rect 446 92 449 698
rect 470 692 473 738
rect 478 642 481 928
rect 486 482 489 858
rect 494 622 497 888
rect 502 862 505 1458
rect 518 1352 521 1798
rect 526 1332 529 1538
rect 550 1032 553 2348
rect 558 2042 561 2228
rect 558 1532 561 1838
rect 566 1772 569 2138
rect 566 1662 569 1678
rect 566 1172 569 1638
rect 574 1122 577 2398
rect 586 1938 590 1941
rect 582 1642 585 1748
rect 582 1452 585 1538
rect 582 1432 585 1448
rect 590 982 593 1828
rect 598 1752 601 2828
rect 610 2748 614 2751
rect 614 2462 617 2618
rect 622 2612 625 3548
rect 630 3342 633 3648
rect 646 3612 649 3768
rect 714 3658 718 3661
rect 734 3582 737 3948
rect 838 3912 841 4078
rect 848 3903 850 3907
rect 854 3903 857 3907
rect 862 3903 864 3907
rect 870 3902 873 3918
rect 934 3862 937 3918
rect 966 3862 969 3878
rect 922 3728 926 3731
rect 848 3703 850 3707
rect 854 3703 857 3707
rect 862 3703 864 3707
rect 750 3652 753 3658
rect 638 3512 641 3548
rect 782 3542 785 3558
rect 634 3328 641 3331
rect 638 3162 641 3328
rect 646 3322 649 3468
rect 654 3432 657 3518
rect 822 3482 825 3558
rect 830 3462 833 3548
rect 846 3542 849 3668
rect 862 3532 865 3538
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 862 3503 864 3507
rect 654 3152 657 3428
rect 674 3238 681 3241
rect 678 3112 681 3238
rect 710 3152 713 3448
rect 734 3312 737 3318
rect 730 3258 734 3261
rect 638 2922 641 2978
rect 634 2688 638 2691
rect 614 2352 617 2458
rect 646 2452 649 2848
rect 662 2552 665 2948
rect 654 2532 657 2548
rect 662 2362 665 2368
rect 654 2292 657 2348
rect 662 2142 665 2188
rect 670 2122 673 3068
rect 678 2942 681 2948
rect 686 2822 689 3148
rect 718 2952 721 3208
rect 726 3152 729 3228
rect 686 2512 689 2808
rect 694 2742 697 2928
rect 718 2872 721 2948
rect 702 2792 705 2838
rect 718 2752 721 2758
rect 694 2632 697 2738
rect 710 2672 713 2678
rect 702 2462 705 2468
rect 698 2348 702 2351
rect 626 2048 630 2051
rect 686 2022 689 2168
rect 606 1762 609 1858
rect 598 1522 601 1528
rect 606 1182 609 1758
rect 614 1472 617 1958
rect 654 1942 657 1948
rect 662 1932 665 1938
rect 646 1852 649 1878
rect 686 1872 689 2018
rect 694 1972 697 2048
rect 626 1548 630 1551
rect 642 1538 646 1541
rect 618 1458 622 1461
rect 654 1392 657 1548
rect 662 1542 665 1548
rect 670 952 673 1568
rect 678 1562 681 1858
rect 686 1622 689 1868
rect 694 1862 697 1968
rect 710 1892 713 2428
rect 718 2342 721 2578
rect 718 2262 721 2338
rect 718 1862 721 2158
rect 710 1852 713 1858
rect 694 1602 697 1828
rect 726 1782 729 3138
rect 734 3122 737 3138
rect 742 3122 745 3318
rect 766 3282 769 3358
rect 754 3268 758 3271
rect 734 2822 737 2848
rect 734 2752 737 2758
rect 734 2572 737 2738
rect 742 2352 745 2368
rect 742 2312 745 2348
rect 734 2172 737 2188
rect 742 2162 745 2308
rect 750 2202 753 2868
rect 782 2802 785 3418
rect 798 3341 801 3348
rect 798 3338 806 3341
rect 806 3312 809 3328
rect 798 3132 801 3148
rect 806 2948 814 2951
rect 758 2652 761 2658
rect 758 2602 761 2648
rect 758 2261 761 2268
rect 758 2258 766 2261
rect 678 1292 681 1558
rect 690 1438 694 1441
rect 702 1122 705 1528
rect 710 1502 713 1768
rect 726 1742 729 1768
rect 734 1552 737 2128
rect 718 1162 721 1548
rect 742 1222 745 1748
rect 750 1542 753 2118
rect 758 1762 761 2258
rect 766 1861 769 2118
rect 778 2058 782 2061
rect 790 1882 793 2948
rect 806 2872 809 2948
rect 814 2892 817 2898
rect 822 2832 825 3128
rect 814 2332 817 2658
rect 822 2492 825 2788
rect 830 2782 833 3338
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 862 3303 864 3307
rect 842 3128 846 3131
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 862 3103 864 3107
rect 830 2662 833 2778
rect 838 2572 841 3098
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 862 2903 864 2907
rect 870 2871 873 3578
rect 878 3362 881 3728
rect 918 3592 921 3728
rect 974 3602 977 4028
rect 998 3822 1001 3858
rect 894 3462 897 3468
rect 878 3282 881 3338
rect 886 3332 889 3348
rect 870 2868 878 2871
rect 882 2738 886 2741
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 862 2703 864 2707
rect 846 2602 849 2658
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 862 2503 864 2507
rect 858 2468 862 2471
rect 798 2272 801 2278
rect 766 1858 774 1861
rect 614 862 617 868
rect 578 858 582 861
rect 574 722 577 738
rect 670 622 673 948
rect 686 942 689 1068
rect 702 962 705 1118
rect 686 852 689 938
rect 702 712 705 948
rect 718 832 721 1148
rect 718 722 721 758
rect 702 662 705 708
rect 750 652 753 1078
rect 758 642 761 1548
rect 766 1102 769 1848
rect 774 1432 777 1808
rect 782 1792 785 1818
rect 806 1652 809 2188
rect 806 1552 809 1648
rect 794 1468 798 1471
rect 774 802 777 1328
rect 790 1132 793 1318
rect 494 552 497 618
rect 534 562 537 588
rect 486 462 489 478
rect 670 472 673 548
rect 550 392 553 468
rect 678 382 681 558
rect 638 62 641 278
rect 686 262 689 398
rect 758 372 761 608
rect 766 422 769 748
rect 774 742 777 798
rect 774 462 777 738
rect 782 502 785 548
rect 798 352 801 1288
rect 814 1262 817 2288
rect 838 2242 841 2318
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 862 2303 864 2307
rect 822 1152 825 1948
rect 838 1872 841 2108
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 862 2103 864 2107
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 862 1903 864 1907
rect 842 1868 846 1871
rect 838 1272 841 1778
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 862 1703 864 1707
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 862 1503 864 1507
rect 870 1462 873 2568
rect 894 2512 897 3198
rect 910 3092 913 3458
rect 902 2802 905 2838
rect 878 2452 881 2458
rect 894 2422 897 2448
rect 894 1962 897 2418
rect 902 2412 905 2428
rect 902 2062 905 2068
rect 902 1672 905 2048
rect 870 1332 873 1458
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 862 1303 864 1307
rect 858 1268 862 1271
rect 838 1152 841 1158
rect 806 1148 814 1151
rect 806 852 809 1148
rect 830 982 833 1108
rect 838 1052 841 1148
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 862 1103 864 1107
rect 838 1018 846 1021
rect 814 952 817 958
rect 806 472 809 478
rect 798 302 801 348
rect 806 282 809 448
rect 814 372 817 538
rect 822 482 825 778
rect 830 752 833 898
rect 838 122 841 1018
rect 846 962 849 978
rect 848 903 850 907
rect 854 903 857 907
rect 862 903 864 907
rect 848 703 850 707
rect 854 703 857 707
rect 862 703 864 707
rect 870 692 873 1278
rect 886 872 889 1188
rect 894 912 897 1158
rect 870 672 873 688
rect 848 503 850 507
rect 854 503 857 507
rect 862 503 864 507
rect 848 303 850 307
rect 854 303 857 307
rect 862 303 864 307
rect 878 282 881 698
rect 902 482 905 1218
rect 910 1062 913 2948
rect 918 2352 921 3258
rect 966 3222 969 3478
rect 982 3472 985 3678
rect 926 3162 929 3208
rect 942 3142 945 3198
rect 990 3072 993 3248
rect 926 2692 929 2848
rect 966 2762 969 2918
rect 946 2758 950 2761
rect 974 2752 977 2918
rect 978 2748 985 2751
rect 926 2352 929 2568
rect 934 2432 937 2508
rect 926 1862 929 2348
rect 934 2342 937 2358
rect 934 2332 937 2338
rect 966 2232 969 2668
rect 974 2432 977 2458
rect 974 2292 977 2308
rect 974 2262 977 2268
rect 922 1668 926 1671
rect 918 1468 926 1471
rect 918 1192 921 1468
rect 910 942 913 948
rect 934 902 937 1148
rect 942 992 945 2188
rect 950 2062 953 2148
rect 950 2002 953 2058
rect 982 1752 985 2748
rect 990 2262 993 2758
rect 998 1852 1001 3818
rect 1014 3582 1017 3798
rect 1018 3538 1025 3541
rect 1022 3532 1025 3538
rect 1014 2442 1017 3328
rect 1030 2952 1033 3838
rect 1038 3592 1041 4248
rect 1062 3862 1065 3898
rect 1086 3862 1089 3868
rect 1062 3712 1065 3858
rect 1094 3642 1097 3858
rect 1110 3702 1113 3958
rect 1118 3662 1121 3668
rect 1054 3552 1057 3638
rect 1126 3632 1129 4528
rect 1158 4462 1161 4578
rect 1174 4162 1177 4498
rect 1194 4448 1198 4451
rect 1190 4282 1193 4358
rect 1206 3902 1209 4138
rect 1214 3911 1217 4378
rect 1262 4352 1265 4668
rect 1310 4462 1313 4748
rect 1318 4662 1321 4898
rect 1352 4803 1354 4807
rect 1358 4803 1361 4807
rect 1366 4803 1368 4807
rect 1342 4682 1345 4768
rect 1450 4748 1454 4751
rect 1342 4482 1345 4678
rect 1352 4603 1354 4607
rect 1358 4603 1361 4607
rect 1366 4603 1368 4607
rect 1462 4562 1465 4858
rect 1534 4672 1537 5068
rect 1662 5002 1665 5098
rect 1782 5052 1785 5058
rect 2384 5003 2386 5007
rect 2390 5003 2393 5007
rect 2398 5003 2400 5007
rect 1730 4948 1734 4951
rect 1872 4903 1874 4907
rect 1878 4903 1881 4907
rect 1886 4903 1888 4907
rect 1358 4552 1361 4558
rect 1262 4332 1265 4348
rect 1278 4122 1281 4138
rect 1286 3952 1289 4148
rect 1294 4122 1297 4128
rect 1274 3928 1281 3931
rect 1214 3908 1222 3911
rect 1162 3878 1166 3881
rect 1178 3878 1185 3881
rect 1182 3872 1185 3878
rect 1038 2891 1041 2948
rect 1038 2888 1046 2891
rect 1038 2792 1041 2888
rect 1054 2862 1057 3148
rect 1006 2272 1009 2438
rect 1014 2282 1017 2438
rect 1022 2302 1025 2468
rect 1046 2412 1049 2768
rect 1006 2082 1009 2128
rect 1022 2092 1025 2298
rect 1054 2252 1057 2538
rect 1062 2412 1065 2978
rect 1078 2891 1081 3018
rect 1086 2982 1089 3438
rect 1094 2942 1097 3018
rect 1074 2888 1081 2891
rect 1086 2852 1089 2908
rect 1102 2852 1105 3618
rect 1150 3362 1153 3758
rect 1174 3632 1177 3648
rect 1174 3562 1177 3628
rect 1174 3528 1182 3531
rect 1174 3492 1177 3528
rect 1142 3312 1145 3338
rect 1150 3332 1153 3338
rect 1130 3128 1134 3131
rect 1094 2848 1102 2851
rect 1070 2652 1073 2738
rect 1086 2662 1089 2788
rect 1070 2612 1073 2648
rect 1094 2582 1097 2848
rect 1102 2742 1105 2798
rect 1102 2662 1105 2678
rect 1110 2632 1113 2728
rect 1118 2722 1121 2848
rect 1134 2832 1137 2948
rect 1158 2842 1161 3258
rect 1166 3162 1169 3428
rect 1174 3282 1177 3488
rect 1206 3472 1209 3898
rect 1222 3882 1225 3888
rect 1234 3878 1238 3881
rect 1250 3738 1254 3741
rect 1214 3672 1217 3678
rect 1198 3442 1201 3448
rect 1178 3148 1182 3151
rect 1178 3138 1185 3141
rect 1170 2948 1174 2951
rect 1126 2682 1129 2758
rect 974 1312 977 1568
rect 994 1488 998 1491
rect 950 1221 953 1278
rect 970 1268 974 1271
rect 958 1262 961 1268
rect 950 1218 958 1221
rect 950 1032 953 1128
rect 946 968 950 971
rect 934 872 937 898
rect 942 872 945 878
rect 918 822 921 848
rect 938 728 942 731
rect 950 532 953 538
rect 958 292 961 1168
rect 982 992 985 1388
rect 982 962 985 988
rect 982 422 985 738
rect 990 632 993 1378
rect 1006 1272 1009 1808
rect 1014 1552 1017 2078
rect 1030 1932 1033 2118
rect 1022 1898 1030 1901
rect 1022 1592 1025 1898
rect 1014 1342 1017 1358
rect 998 1082 1001 1088
rect 998 952 1001 968
rect 998 752 1001 758
rect 998 672 1001 748
rect 1006 742 1009 1258
rect 1014 1061 1017 1168
rect 1022 1152 1025 1418
rect 1014 1058 1022 1061
rect 1030 992 1033 1408
rect 1022 942 1025 958
rect 1006 662 1009 738
rect 990 342 993 628
rect 1014 572 1017 898
rect 1022 862 1025 938
rect 1014 362 1017 568
rect 1022 562 1025 568
rect 1014 332 1017 358
rect 1038 222 1041 2118
rect 1054 1572 1057 2248
rect 1062 1582 1065 2408
rect 1102 2032 1105 2308
rect 1086 1872 1089 1888
rect 1054 1022 1057 1348
rect 1062 1302 1065 1338
rect 1070 1082 1073 1308
rect 1046 881 1049 998
rect 1094 952 1097 2018
rect 1102 1902 1105 2028
rect 1090 928 1094 931
rect 1046 878 1054 881
rect 1102 842 1105 1728
rect 1110 1542 1113 2608
rect 1118 2572 1121 2668
rect 1142 2572 1145 2798
rect 1158 2722 1161 2758
rect 1150 2692 1153 2718
rect 1166 2692 1169 2888
rect 1174 2712 1177 2728
rect 1182 2722 1185 3138
rect 1130 2338 1134 2341
rect 1142 2042 1145 2558
rect 1118 1902 1121 1908
rect 1126 1892 1129 1918
rect 1142 1872 1145 1928
rect 1118 1562 1121 1698
rect 1126 1602 1129 1838
rect 1118 1538 1126 1541
rect 1110 1462 1113 1538
rect 1118 1532 1121 1538
rect 1134 1082 1137 1798
rect 1142 1741 1145 1868
rect 1158 1842 1161 2438
rect 1166 2152 1169 2348
rect 1190 2312 1193 3158
rect 1198 3062 1201 3438
rect 1206 3138 1214 3141
rect 1206 3092 1209 3138
rect 1206 2992 1209 3088
rect 1222 3062 1225 3068
rect 1142 1738 1150 1741
rect 1142 1662 1145 1668
rect 1158 1182 1161 1838
rect 1166 1552 1169 2148
rect 1174 2072 1177 2078
rect 1182 2052 1185 2258
rect 1166 1452 1169 1458
rect 1166 1292 1169 1388
rect 1174 1212 1177 2018
rect 1182 1422 1185 2048
rect 1190 1982 1193 2108
rect 1198 2082 1201 2458
rect 1206 2272 1209 2828
rect 1214 2342 1217 2798
rect 1222 2182 1225 2568
rect 1230 2442 1233 3738
rect 1278 3732 1281 3928
rect 1286 3922 1289 3948
rect 1242 3668 1246 3671
rect 1242 3648 1249 3651
rect 1246 3372 1249 3648
rect 1270 3472 1273 3588
rect 1278 3542 1281 3728
rect 1270 3452 1273 3458
rect 1238 2552 1241 3108
rect 1230 2392 1233 2428
rect 1238 2142 1241 2278
rect 1246 2262 1249 3368
rect 1254 2882 1257 2948
rect 1262 2942 1265 3188
rect 1262 2582 1265 2898
rect 1270 2322 1273 2988
rect 1278 2902 1281 3458
rect 1294 3382 1297 4028
rect 1302 3872 1305 4268
rect 1310 3862 1313 4458
rect 1342 4422 1345 4448
rect 1322 3868 1326 3871
rect 1302 3752 1305 3858
rect 1302 3492 1305 3748
rect 1310 3648 1318 3651
rect 1286 3001 1289 3258
rect 1310 3082 1313 3648
rect 1334 3612 1337 3628
rect 1322 3338 1326 3341
rect 1334 3272 1337 3488
rect 1342 3482 1345 4418
rect 1352 4403 1354 4407
rect 1358 4403 1361 4407
rect 1366 4403 1368 4407
rect 1454 4372 1457 4548
rect 1462 4452 1465 4538
rect 1462 4292 1465 4448
rect 1470 4361 1473 4568
rect 1470 4358 1478 4361
rect 1542 4331 1545 4508
rect 1538 4328 1545 4331
rect 1352 4203 1354 4207
rect 1358 4203 1361 4207
rect 1366 4203 1368 4207
rect 1390 4052 1393 4188
rect 1478 4152 1481 4158
rect 1352 4003 1354 4007
rect 1358 4003 1361 4007
rect 1366 4003 1368 4007
rect 1374 3942 1377 4008
rect 1350 3872 1353 3878
rect 1374 3862 1377 3938
rect 1390 3912 1393 4048
rect 1446 4042 1449 4048
rect 1352 3803 1354 3807
rect 1358 3803 1361 3807
rect 1366 3803 1368 3807
rect 1350 3682 1353 3688
rect 1374 3682 1377 3858
rect 1414 3832 1417 3928
rect 1352 3603 1354 3607
rect 1358 3603 1361 3607
rect 1366 3603 1368 3607
rect 1286 2998 1294 3001
rect 1294 2872 1297 2988
rect 1302 2868 1310 2871
rect 1286 2852 1289 2858
rect 1270 2282 1273 2318
rect 1278 2202 1281 2348
rect 1218 2138 1222 2141
rect 1206 1962 1209 2058
rect 1214 2052 1217 2078
rect 1246 2062 1249 2168
rect 1230 1992 1233 2058
rect 1254 2002 1257 2158
rect 1190 1411 1193 1918
rect 1198 1772 1201 1878
rect 1182 1408 1193 1411
rect 1166 1022 1169 1128
rect 1118 952 1121 958
rect 1166 952 1169 1018
rect 1174 952 1177 958
rect 1130 948 1134 951
rect 1062 792 1065 798
rect 1110 672 1113 928
rect 1118 912 1121 948
rect 1118 762 1121 908
rect 1182 812 1185 1408
rect 1190 1232 1193 1248
rect 1190 752 1193 1048
rect 1118 352 1121 668
rect 1190 662 1193 748
rect 1198 682 1201 1678
rect 1206 1672 1209 1878
rect 1206 1032 1209 1628
rect 1222 1412 1225 1738
rect 1230 1552 1233 1988
rect 1214 1352 1217 1358
rect 1222 1161 1225 1328
rect 1218 1158 1225 1161
rect 1214 942 1217 1098
rect 1230 852 1233 1528
rect 1238 1042 1241 1588
rect 1254 1462 1257 1998
rect 1246 862 1249 1328
rect 1254 1062 1257 1458
rect 1262 1452 1265 1518
rect 1270 1462 1273 1468
rect 1278 1462 1281 1468
rect 1278 1272 1281 1448
rect 1246 812 1249 818
rect 1206 682 1209 788
rect 1222 752 1225 758
rect 1214 412 1217 728
rect 1238 152 1241 568
rect 1246 402 1249 648
rect 1254 352 1257 1038
rect 1262 542 1265 558
rect 1270 472 1273 698
rect 1278 642 1281 1028
rect 1286 962 1289 2268
rect 1294 1862 1297 2868
rect 1302 2852 1305 2868
rect 1314 2848 1318 2851
rect 1326 2642 1329 3068
rect 1334 3062 1337 3068
rect 1334 2812 1337 2888
rect 1326 2552 1329 2588
rect 1334 2532 1337 2668
rect 1342 2632 1345 3448
rect 1352 3403 1354 3407
rect 1358 3403 1361 3407
rect 1366 3403 1368 3407
rect 1352 3203 1354 3207
rect 1358 3203 1361 3207
rect 1366 3203 1368 3207
rect 1402 3168 1406 3171
rect 1374 3082 1377 3168
rect 1402 3128 1406 3131
rect 1382 3052 1385 3088
rect 1352 3003 1354 3007
rect 1358 3003 1361 3007
rect 1366 3003 1368 3007
rect 1374 2922 1377 3048
rect 1352 2803 1354 2807
rect 1358 2803 1361 2807
rect 1366 2803 1368 2807
rect 1352 2603 1354 2607
rect 1358 2603 1361 2607
rect 1366 2603 1368 2607
rect 1398 2602 1401 2778
rect 1414 2691 1417 3828
rect 1446 3792 1449 4038
rect 1454 4002 1457 4138
rect 1566 4102 1569 4748
rect 1606 4732 1609 4768
rect 1714 4748 1718 4751
rect 1614 4732 1617 4748
rect 1606 4622 1609 4728
rect 1646 4102 1649 4548
rect 1654 4272 1657 4698
rect 1662 4482 1665 4528
rect 1682 4268 1686 4271
rect 1654 4062 1657 4258
rect 1670 4252 1673 4258
rect 1422 3742 1425 3768
rect 1478 3552 1481 3738
rect 1486 3672 1489 3878
rect 1494 3642 1497 3828
rect 1502 3782 1505 4058
rect 1502 3748 1510 3751
rect 1446 3512 1449 3538
rect 1430 3508 1438 3511
rect 1422 2722 1425 3488
rect 1430 3272 1433 3508
rect 1430 3262 1433 3268
rect 1438 3112 1441 3478
rect 1454 3442 1457 3458
rect 1486 3362 1489 3548
rect 1494 3372 1497 3448
rect 1502 3351 1505 3748
rect 1534 3732 1537 3798
rect 1514 3438 1518 3441
rect 1502 3348 1513 3351
rect 1478 3328 1486 3331
rect 1478 3252 1481 3328
rect 1458 3248 1462 3251
rect 1426 2708 1430 2711
rect 1414 2688 1425 2691
rect 1406 2658 1414 2661
rect 1302 2262 1305 2438
rect 1342 2412 1345 2428
rect 1406 2412 1409 2658
rect 1422 2552 1425 2688
rect 1352 2403 1354 2407
rect 1358 2403 1361 2407
rect 1366 2403 1368 2407
rect 1386 2398 1390 2401
rect 1302 2252 1305 2258
rect 1302 1681 1305 2158
rect 1310 1882 1313 2358
rect 1370 2348 1377 2351
rect 1374 2292 1377 2348
rect 1366 2278 1374 2281
rect 1334 2182 1337 2208
rect 1322 2068 1326 2071
rect 1318 1872 1321 1938
rect 1326 1861 1329 2058
rect 1318 1858 1329 1861
rect 1302 1678 1310 1681
rect 1318 1412 1321 1858
rect 1326 1652 1329 1738
rect 1334 1492 1337 2018
rect 1342 1942 1345 2248
rect 1366 2222 1369 2278
rect 1352 2203 1354 2207
rect 1358 2203 1361 2207
rect 1366 2203 1368 2207
rect 1382 2062 1385 2388
rect 1398 2342 1401 2398
rect 1414 2282 1417 2518
rect 1430 2352 1433 2358
rect 1378 2058 1382 2061
rect 1352 2003 1354 2007
rect 1358 2003 1361 2007
rect 1366 2003 1368 2007
rect 1374 1902 1377 1908
rect 1374 1812 1377 1858
rect 1352 1803 1354 1807
rect 1358 1803 1361 1807
rect 1366 1803 1368 1807
rect 1352 1603 1354 1607
rect 1358 1603 1361 1607
rect 1366 1603 1368 1607
rect 1374 1472 1377 1808
rect 1382 1752 1385 1798
rect 1390 1462 1393 2278
rect 1422 2252 1425 2328
rect 1430 2132 1433 2348
rect 1438 2302 1441 3088
rect 1454 3061 1457 3168
rect 1462 3132 1465 3138
rect 1450 3058 1457 3061
rect 1450 3048 1454 3051
rect 1462 2972 1465 3118
rect 1470 3102 1473 3218
rect 1478 3182 1481 3248
rect 1478 3012 1481 3128
rect 1486 3062 1489 3278
rect 1498 3238 1502 3241
rect 1510 3232 1513 3348
rect 1526 3262 1529 3558
rect 1538 3518 1542 3521
rect 1534 3472 1537 3508
rect 1550 3412 1553 3648
rect 1538 3308 1542 3311
rect 1530 3248 1534 3251
rect 1494 3132 1497 3158
rect 1478 2872 1481 2898
rect 1446 2532 1449 2598
rect 1406 1932 1409 2058
rect 1422 2042 1425 2058
rect 1418 1958 1422 1961
rect 1406 1752 1409 1928
rect 1422 1832 1425 1898
rect 1418 1748 1422 1751
rect 1430 1722 1433 1968
rect 1422 1662 1425 1668
rect 1398 1612 1401 1648
rect 1352 1403 1354 1407
rect 1358 1403 1361 1407
rect 1366 1403 1368 1407
rect 1294 1012 1297 1108
rect 1302 1082 1305 1268
rect 1310 1202 1313 1208
rect 1330 1158 1334 1161
rect 1278 552 1281 558
rect 1278 372 1281 548
rect 1294 542 1297 548
rect 1286 252 1289 538
rect 1302 462 1305 948
rect 1298 438 1302 441
rect 1310 342 1313 828
rect 1318 682 1321 988
rect 1334 612 1337 918
rect 1342 592 1345 1378
rect 1374 1252 1377 1428
rect 1352 1203 1354 1207
rect 1358 1203 1361 1207
rect 1366 1203 1368 1207
rect 1352 1003 1354 1007
rect 1358 1003 1361 1007
rect 1366 1003 1368 1007
rect 1352 803 1354 807
rect 1358 803 1361 807
rect 1366 803 1368 807
rect 1374 792 1377 1148
rect 1382 702 1385 1288
rect 1390 902 1393 1428
rect 1398 1202 1401 1608
rect 1414 1561 1417 1578
rect 1414 1558 1422 1561
rect 1406 1212 1409 1268
rect 1414 1192 1417 1478
rect 1414 952 1417 958
rect 1374 672 1377 678
rect 1352 603 1354 607
rect 1358 603 1361 607
rect 1366 603 1368 607
rect 1342 572 1345 588
rect 1382 562 1385 658
rect 1422 622 1425 1558
rect 1430 1532 1433 1598
rect 1430 1282 1433 1288
rect 1438 1122 1441 1968
rect 1446 1952 1449 2528
rect 1454 2522 1457 2728
rect 1462 2522 1465 2568
rect 1454 2452 1457 2518
rect 1470 2412 1473 2418
rect 1446 1472 1449 1888
rect 1454 1882 1457 2388
rect 1462 2192 1465 2348
rect 1470 2012 1473 2408
rect 1486 2292 1489 2718
rect 1494 2501 1497 3128
rect 1502 2732 1505 2748
rect 1494 2498 1502 2501
rect 1498 2468 1502 2471
rect 1478 2258 1486 2261
rect 1478 2222 1481 2258
rect 1486 2212 1489 2218
rect 1486 2132 1489 2208
rect 1494 2112 1497 2218
rect 1462 1972 1465 1988
rect 1462 1572 1465 1718
rect 1470 1642 1473 1988
rect 1494 1782 1497 2058
rect 1502 2012 1505 2338
rect 1446 1242 1449 1458
rect 1454 1262 1457 1568
rect 1462 1392 1465 1568
rect 1478 1561 1481 1688
rect 1502 1672 1505 1938
rect 1510 1872 1513 2768
rect 1518 2502 1521 3108
rect 1542 3082 1545 3148
rect 1534 2712 1537 2968
rect 1542 2852 1545 3078
rect 1526 2572 1529 2578
rect 1526 2462 1529 2558
rect 1534 2512 1537 2708
rect 1542 2462 1545 2818
rect 1550 2412 1553 3408
rect 1558 2992 1561 3778
rect 1574 3362 1577 3928
rect 1582 3742 1585 3788
rect 1602 3748 1606 3751
rect 1582 3671 1585 3738
rect 1582 3668 1590 3671
rect 1582 3502 1585 3548
rect 1590 3482 1593 3658
rect 1598 3342 1601 3748
rect 1618 3738 1622 3741
rect 1630 3632 1633 3638
rect 1638 3582 1641 3738
rect 1614 3532 1617 3548
rect 1630 3531 1633 3568
rect 1626 3528 1633 3531
rect 1622 3511 1625 3518
rect 1618 3508 1625 3511
rect 1606 3492 1609 3508
rect 1566 3142 1569 3318
rect 1574 3312 1577 3318
rect 1582 3252 1585 3278
rect 1590 3192 1593 3308
rect 1606 3252 1609 3488
rect 1566 3082 1569 3088
rect 1598 3052 1601 3058
rect 1558 2851 1561 2858
rect 1558 2848 1566 2851
rect 1582 2832 1585 3038
rect 1590 2882 1593 2898
rect 1558 2782 1561 2808
rect 1558 2752 1561 2778
rect 1566 2712 1569 2718
rect 1558 2561 1561 2678
rect 1558 2558 1566 2561
rect 1558 2422 1561 2478
rect 1574 2471 1577 2778
rect 1582 2772 1585 2828
rect 1590 2722 1593 2858
rect 1598 2792 1601 3018
rect 1606 2882 1609 3248
rect 1614 3242 1617 3248
rect 1630 3151 1633 3158
rect 1626 3148 1633 3151
rect 1626 3138 1630 3141
rect 1622 3082 1625 3108
rect 1638 3072 1641 3578
rect 1646 3142 1649 3548
rect 1654 3202 1657 4058
rect 1662 3922 1665 4018
rect 1662 3722 1665 3918
rect 1670 3582 1673 3948
rect 1662 3552 1665 3568
rect 1678 3522 1681 4038
rect 1686 3742 1689 4108
rect 1694 4062 1697 4558
rect 1694 3812 1697 3978
rect 1694 3632 1697 3738
rect 1694 3542 1697 3548
rect 1686 3522 1689 3538
rect 1638 3042 1641 3068
rect 1646 3062 1649 3138
rect 1662 3122 1665 3518
rect 1670 3152 1673 3158
rect 1694 3142 1697 3148
rect 1654 3072 1657 3078
rect 1626 2978 1630 2981
rect 1638 2932 1641 2938
rect 1594 2708 1598 2711
rect 1566 2468 1577 2471
rect 1622 2472 1625 2598
rect 1630 2532 1633 2858
rect 1646 2842 1649 2968
rect 1654 2952 1657 2958
rect 1646 2691 1649 2838
rect 1662 2752 1665 3118
rect 1646 2688 1654 2691
rect 1518 2322 1521 2328
rect 1518 2032 1521 2128
rect 1526 2122 1529 2348
rect 1542 2152 1545 2358
rect 1550 2272 1553 2318
rect 1538 2138 1542 2141
rect 1526 1822 1529 2088
rect 1558 2072 1561 2318
rect 1566 2182 1569 2468
rect 1578 2458 1582 2461
rect 1582 2082 1585 2378
rect 1638 2372 1641 2388
rect 1634 2338 1638 2341
rect 1602 2318 1606 2321
rect 1590 2182 1593 2188
rect 1606 2132 1609 2288
rect 1566 2072 1569 2078
rect 1582 2022 1585 2078
rect 1606 2052 1609 2128
rect 1582 1942 1585 1968
rect 1606 1942 1609 1968
rect 1614 1952 1617 2328
rect 1646 2212 1649 2448
rect 1642 2138 1646 2141
rect 1590 1932 1593 1938
rect 1582 1922 1585 1928
rect 1566 1852 1569 1888
rect 1622 1882 1625 1948
rect 1622 1852 1625 1878
rect 1630 1852 1633 1898
rect 1494 1668 1502 1671
rect 1478 1558 1486 1561
rect 1470 1522 1473 1538
rect 1494 1502 1497 1668
rect 1506 1558 1510 1561
rect 1526 1532 1529 1538
rect 1330 498 1337 501
rect 1334 322 1337 498
rect 1352 403 1354 407
rect 1358 403 1361 407
rect 1366 403 1368 407
rect 1382 392 1385 558
rect 1422 552 1425 618
rect 1438 492 1441 998
rect 1462 992 1465 1358
rect 1470 872 1473 1468
rect 1506 1458 1510 1461
rect 1486 1252 1489 1458
rect 1478 1122 1481 1248
rect 1486 852 1489 1248
rect 1494 692 1497 1338
rect 1518 972 1521 1428
rect 1526 1332 1529 1528
rect 1526 1152 1529 1158
rect 1534 902 1537 1648
rect 1542 1492 1545 1538
rect 1558 1312 1561 1798
rect 1566 1752 1569 1768
rect 1574 1742 1577 1848
rect 1566 1582 1569 1678
rect 1574 1522 1577 1738
rect 1566 1472 1569 1488
rect 1570 1468 1574 1471
rect 1566 1428 1574 1431
rect 1566 1252 1569 1428
rect 1582 1352 1585 1668
rect 1590 802 1593 1428
rect 1606 1342 1609 1348
rect 1614 1302 1617 1848
rect 1626 1708 1633 1711
rect 1630 1632 1633 1708
rect 1638 1552 1641 2098
rect 1646 1832 1649 1928
rect 1654 1762 1657 2188
rect 1650 1668 1657 1671
rect 1634 1468 1638 1471
rect 1654 1452 1657 1668
rect 1618 1148 1622 1151
rect 1638 1082 1641 1088
rect 1494 662 1497 688
rect 1450 658 1454 661
rect 1352 203 1354 207
rect 1358 203 1361 207
rect 1366 203 1368 207
rect 848 103 850 107
rect 854 103 857 107
rect 862 103 864 107
rect 1374 82 1377 378
rect 1526 292 1529 708
rect 1534 432 1537 718
rect 1614 562 1617 808
rect 1646 792 1649 1268
rect 1654 1252 1657 1328
rect 1654 1002 1657 1248
rect 1662 1132 1665 2748
rect 1670 2392 1673 3078
rect 1686 3032 1689 3138
rect 1702 3112 1705 4408
rect 1718 4152 1721 4348
rect 1718 4072 1721 4078
rect 1734 4062 1737 4218
rect 1710 3992 1713 4058
rect 1742 4022 1745 4118
rect 1710 3452 1713 3988
rect 1742 3932 1745 3938
rect 1750 3932 1753 4248
rect 1774 4081 1777 4218
rect 1774 4078 1782 4081
rect 1742 3862 1745 3888
rect 1678 2642 1681 2758
rect 1670 2352 1673 2358
rect 1670 2142 1673 2158
rect 1670 1732 1673 1748
rect 1678 1671 1681 2638
rect 1686 2602 1689 2828
rect 1694 2722 1697 2738
rect 1686 2592 1689 2598
rect 1702 2572 1705 2988
rect 1710 2902 1713 3218
rect 1718 3082 1721 3178
rect 1726 3092 1729 3748
rect 1734 3172 1737 3588
rect 1742 3462 1745 3838
rect 1750 3532 1753 3928
rect 1742 3282 1745 3288
rect 1734 2952 1737 2978
rect 1714 2748 1718 2751
rect 1710 2652 1713 2718
rect 1726 2552 1729 2628
rect 1702 2341 1705 2348
rect 1698 2338 1705 2341
rect 1690 2318 1697 2321
rect 1694 2232 1697 2318
rect 1718 2172 1721 2218
rect 1726 2202 1729 2208
rect 1686 2122 1689 2168
rect 1698 2128 1702 2131
rect 1718 2122 1721 2168
rect 1686 1842 1689 2008
rect 1694 1932 1697 2058
rect 1726 1962 1729 1988
rect 1702 1942 1705 1958
rect 1722 1938 1729 1941
rect 1690 1838 1697 1841
rect 1678 1668 1686 1671
rect 1674 1648 1678 1651
rect 1678 1472 1681 1488
rect 1674 1258 1678 1261
rect 1662 952 1665 968
rect 1670 952 1673 958
rect 1678 932 1681 948
rect 1686 872 1689 1668
rect 1694 1352 1697 1838
rect 1718 1762 1721 1928
rect 1726 1922 1729 1938
rect 1718 1582 1721 1758
rect 1706 1488 1710 1491
rect 1702 1452 1705 1458
rect 1718 1452 1721 1558
rect 1726 1522 1729 1678
rect 1726 1472 1729 1518
rect 1734 1442 1737 2948
rect 1742 2812 1745 3008
rect 1750 2882 1753 3398
rect 1758 2842 1761 4078
rect 1790 3902 1793 3938
rect 1778 3878 1782 3881
rect 1798 3852 1801 4728
rect 1846 4402 1849 4468
rect 1794 3648 1798 3651
rect 1790 3628 1798 3631
rect 1790 3562 1793 3628
rect 1798 3562 1801 3588
rect 1766 3382 1769 3548
rect 1774 3362 1777 3508
rect 1782 3442 1785 3558
rect 1790 3542 1793 3548
rect 1806 3502 1809 4168
rect 1814 3872 1817 4118
rect 1822 3932 1825 4258
rect 1830 4162 1833 4358
rect 1846 4062 1849 4398
rect 1854 4142 1857 4768
rect 2102 4761 2105 4898
rect 2158 4792 2161 4918
rect 2098 4758 2105 4761
rect 2182 4732 2185 4858
rect 2222 4801 2225 4958
rect 2218 4798 2225 4801
rect 1872 4703 1874 4707
rect 1878 4703 1881 4707
rect 1886 4703 1888 4707
rect 1872 4503 1874 4507
rect 1878 4503 1881 4507
rect 1886 4503 1888 4507
rect 1872 4303 1874 4307
rect 1878 4303 1881 4307
rect 1886 4303 1888 4307
rect 1878 4122 1881 4138
rect 1872 4103 1874 4107
rect 1878 4103 1881 4107
rect 1886 4103 1888 4107
rect 1838 3872 1841 3998
rect 1822 3862 1825 3868
rect 1830 3848 1838 3851
rect 1830 3582 1833 3848
rect 1838 3682 1841 3688
rect 1822 3512 1825 3548
rect 1790 3462 1793 3468
rect 1778 3338 1782 3341
rect 1782 3132 1785 3138
rect 1766 2912 1769 2978
rect 1782 2872 1785 2988
rect 1758 2772 1761 2838
rect 1758 2742 1761 2748
rect 1758 2582 1761 2738
rect 1766 2561 1769 2858
rect 1782 2632 1785 2718
rect 1790 2642 1793 3268
rect 1798 2902 1801 3468
rect 1810 3458 1814 3461
rect 1806 2952 1809 3378
rect 1814 2942 1817 3268
rect 1822 3012 1825 3498
rect 1818 2938 1822 2941
rect 1830 2932 1833 3578
rect 1838 3152 1841 3588
rect 1846 3552 1849 4048
rect 1854 4002 1857 4038
rect 1894 3952 1897 4608
rect 1950 4372 1953 4528
rect 1918 4192 1921 4368
rect 1926 4272 1929 4368
rect 1906 4138 1910 4141
rect 1926 4092 1929 4108
rect 1918 4082 1921 4088
rect 1872 3903 1874 3907
rect 1878 3903 1881 3907
rect 1886 3903 1888 3907
rect 1918 3872 1921 4058
rect 1926 3862 1929 4088
rect 1934 4072 1937 4088
rect 1942 4062 1945 4078
rect 1894 3852 1897 3858
rect 1934 3772 1937 3938
rect 1942 3792 1945 3938
rect 1934 3752 1937 3768
rect 1906 3738 1910 3741
rect 1934 3722 1937 3728
rect 1942 3711 1945 3788
rect 1950 3742 1953 4118
rect 1950 3722 1953 3738
rect 1942 3708 1953 3711
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1886 3703 1888 3707
rect 1858 3678 1862 3681
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1886 3503 1888 3507
rect 1850 3458 1854 3461
rect 1838 2942 1841 3068
rect 1762 2558 1769 2561
rect 1742 2202 1745 2348
rect 1750 2342 1753 2418
rect 1774 2402 1777 2608
rect 1742 2172 1745 2188
rect 1750 2152 1753 2218
rect 1758 2132 1761 2318
rect 1758 2072 1761 2078
rect 1750 1972 1753 2008
rect 1742 1932 1745 1968
rect 1750 1932 1753 1948
rect 1742 1562 1745 1758
rect 1750 1652 1753 1888
rect 1758 1862 1761 1978
rect 1766 1812 1769 2088
rect 1774 1942 1777 2358
rect 1782 2062 1785 2628
rect 1782 1982 1785 1998
rect 1782 1972 1785 1978
rect 1790 1911 1793 2628
rect 1798 2462 1801 2728
rect 1806 2362 1809 2878
rect 1814 2662 1817 2928
rect 1830 2732 1833 2738
rect 1782 1908 1793 1911
rect 1782 1732 1785 1908
rect 1790 1762 1793 1828
rect 1742 1542 1745 1548
rect 1766 1532 1769 1628
rect 1758 1492 1761 1498
rect 1758 1472 1761 1488
rect 1746 1468 1750 1471
rect 1714 1348 1718 1351
rect 1702 882 1705 908
rect 1678 552 1681 628
rect 1570 488 1574 491
rect 1534 361 1537 368
rect 1534 358 1542 361
rect 1590 352 1593 378
rect 1566 222 1569 328
rect 1582 182 1585 318
rect 1670 242 1673 448
rect 1678 222 1681 548
rect 1694 482 1697 868
rect 1710 852 1713 858
rect 1718 832 1721 868
rect 1694 462 1697 478
rect 1702 82 1705 528
rect 1726 492 1729 1438
rect 1766 1342 1769 1528
rect 1742 842 1745 1318
rect 1742 312 1745 788
rect 1766 602 1769 1108
rect 1774 492 1777 1518
rect 1782 1472 1785 1678
rect 1790 1602 1793 1758
rect 1790 1442 1793 1598
rect 1790 1352 1793 1358
rect 1782 1342 1785 1348
rect 1798 1082 1801 2358
rect 1814 2262 1817 2658
rect 1830 2472 1833 2548
rect 1838 2462 1841 2688
rect 1814 1802 1817 1968
rect 1814 1652 1817 1768
rect 1822 1722 1825 2448
rect 1830 2332 1833 2388
rect 1838 2352 1841 2408
rect 1846 2382 1849 3458
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1886 3303 1888 3307
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1886 3103 1888 3107
rect 1894 3082 1897 3098
rect 1858 3058 1862 3061
rect 1870 3052 1873 3068
rect 1894 3052 1897 3068
rect 1902 3052 1905 3358
rect 1854 3012 1857 3028
rect 1854 2662 1857 2898
rect 1862 2722 1865 3048
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1886 2903 1888 2907
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1886 2703 1888 2707
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1886 2503 1888 2507
rect 1882 2468 1886 2471
rect 1894 2462 1897 3038
rect 1902 2752 1905 3048
rect 1918 3042 1921 3128
rect 1910 2912 1913 3008
rect 1918 2912 1921 2918
rect 1902 2562 1905 2618
rect 1902 2472 1905 2478
rect 1838 2342 1841 2348
rect 1846 2332 1849 2368
rect 1878 2342 1881 2368
rect 1910 2322 1913 2908
rect 1926 2802 1929 3118
rect 1918 2562 1921 2768
rect 1934 2712 1937 3328
rect 1942 3292 1945 3378
rect 1950 3022 1953 3708
rect 1958 3352 1961 4548
rect 1986 4448 1990 4451
rect 1998 4242 2001 4458
rect 1966 4212 1969 4238
rect 1966 4062 1969 4068
rect 1958 2962 1961 2978
rect 1950 2952 1953 2958
rect 1966 2952 1969 3148
rect 1974 2952 1977 3998
rect 1982 3502 1985 3928
rect 1934 2602 1937 2708
rect 1918 2552 1921 2558
rect 1942 2552 1945 2838
rect 1942 2532 1945 2548
rect 1918 2452 1921 2478
rect 1930 2458 1934 2461
rect 1930 2448 1934 2451
rect 1942 2422 1945 2508
rect 1958 2442 1961 2748
rect 1966 2622 1969 2948
rect 1966 2602 1969 2618
rect 1946 2418 1953 2421
rect 1926 2352 1929 2368
rect 1862 2292 1865 2308
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1886 2303 1888 2307
rect 1830 2051 1833 2198
rect 1862 2148 1870 2151
rect 1850 2058 1854 2061
rect 1830 2048 1841 2051
rect 1830 1992 1833 2028
rect 1782 732 1785 738
rect 1782 712 1785 728
rect 1798 672 1801 708
rect 1806 652 1809 1458
rect 1814 1292 1817 1578
rect 1822 1482 1825 1618
rect 1830 1572 1833 1898
rect 1830 1432 1833 1498
rect 1814 662 1817 1128
rect 1830 912 1833 1408
rect 1838 1312 1841 2048
rect 1850 1988 1854 1991
rect 1862 1982 1865 2148
rect 1894 2112 1897 2258
rect 1942 2232 1945 2258
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1886 2103 1888 2107
rect 1926 2082 1929 2228
rect 1934 2142 1937 2148
rect 1882 2068 1886 2071
rect 1918 2052 1921 2068
rect 1910 1942 1913 1948
rect 1926 1942 1929 2078
rect 1934 2062 1937 2078
rect 1934 2042 1937 2048
rect 1942 2032 1945 2188
rect 1882 1938 1886 1941
rect 1846 1562 1849 1758
rect 1854 1632 1857 1938
rect 1918 1932 1921 1938
rect 1950 1931 1953 2418
rect 1966 2352 1969 2448
rect 1958 2302 1961 2348
rect 1974 2312 1977 2938
rect 1982 2852 1985 3078
rect 1990 2762 1993 4198
rect 1998 3871 2001 4238
rect 2006 3952 2009 4718
rect 2018 4448 2022 4451
rect 2014 4062 2017 4318
rect 2014 3922 2017 3938
rect 1998 3868 2006 3871
rect 2006 3842 2009 3858
rect 1998 2742 2001 3218
rect 2006 3162 2009 3838
rect 2014 3642 2017 3918
rect 2022 3782 2025 4268
rect 2046 4052 2049 4298
rect 2054 4282 2057 4648
rect 2074 4458 2078 4461
rect 2058 4258 2062 4261
rect 2070 4232 2073 4408
rect 2086 4262 2089 4438
rect 2094 4352 2097 4448
rect 2038 3952 2041 3958
rect 2034 3938 2038 3941
rect 2038 3852 2041 3858
rect 2014 3232 2017 3438
rect 2022 3372 2025 3428
rect 2022 3232 2025 3238
rect 1990 2732 1993 2738
rect 1958 2292 1961 2298
rect 1946 1928 1953 1931
rect 1958 2158 1966 2161
rect 1862 1892 1865 1908
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1886 1903 1888 1907
rect 1862 1682 1865 1868
rect 1894 1852 1897 1908
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1886 1703 1888 1707
rect 1838 1112 1841 1248
rect 1846 852 1849 1458
rect 1854 1182 1857 1338
rect 1862 1302 1865 1558
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1886 1503 1888 1507
rect 1886 1462 1889 1468
rect 1894 1442 1897 1528
rect 1902 1452 1905 1508
rect 1910 1452 1913 1458
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1886 1303 1888 1307
rect 1870 1262 1873 1288
rect 1894 1212 1897 1358
rect 1790 542 1793 548
rect 1798 542 1801 558
rect 1770 478 1774 481
rect 1762 338 1766 341
rect 1774 182 1777 448
rect 1782 422 1785 538
rect 1806 412 1809 648
rect 1814 632 1817 658
rect 1854 442 1857 1068
rect 1862 742 1865 1198
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1886 1103 1888 1107
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1886 903 1888 907
rect 1862 712 1865 738
rect 1894 732 1897 1208
rect 1902 1012 1905 1438
rect 1910 982 1913 1268
rect 1918 1252 1921 1788
rect 1934 1542 1937 1898
rect 1930 1498 1934 1501
rect 1930 1468 1934 1471
rect 1942 1462 1945 1738
rect 1950 1602 1953 1818
rect 1958 1712 1961 2158
rect 1974 1941 1977 1948
rect 1970 1938 1977 1941
rect 1938 1448 1942 1451
rect 1918 992 1921 1248
rect 1926 1052 1929 1278
rect 1930 1048 1934 1051
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1886 703 1888 707
rect 1910 512 1913 888
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1886 503 1888 507
rect 1898 478 1902 481
rect 1918 392 1921 978
rect 1934 492 1937 498
rect 1942 432 1945 1328
rect 1950 922 1953 1598
rect 1958 1332 1961 1498
rect 1966 1442 1969 1868
rect 1958 1242 1961 1248
rect 1966 1042 1969 1338
rect 1966 932 1969 948
rect 1958 702 1961 728
rect 1962 698 1966 701
rect 1974 552 1977 1548
rect 1982 1362 1985 2578
rect 1990 2312 1993 2488
rect 1990 2022 1993 2298
rect 1998 2272 2001 2638
rect 2006 2292 2009 3148
rect 2014 2442 2017 3228
rect 2030 3152 2033 3398
rect 2038 3262 2041 3528
rect 2022 3062 2025 3118
rect 2022 2492 2025 2748
rect 2022 2462 2025 2468
rect 1998 1982 2001 2068
rect 2006 1962 2009 2228
rect 2022 2222 2025 2278
rect 2014 2032 2017 2048
rect 1990 1692 1993 1758
rect 1994 1558 1998 1561
rect 1990 1532 1993 1538
rect 1982 392 1985 1338
rect 1990 1222 1993 1508
rect 1998 1342 2001 1548
rect 2006 1532 2009 1938
rect 2014 1652 2017 1658
rect 2006 1442 2009 1448
rect 2014 642 2017 1528
rect 2022 1332 2025 2208
rect 2030 2162 2033 2868
rect 2038 2332 2041 3238
rect 2046 3182 2049 4048
rect 2054 3872 2057 4048
rect 2078 4042 2081 4058
rect 2078 3952 2081 4008
rect 2086 3952 2089 4258
rect 2102 3872 2105 4558
rect 2126 4252 2129 4658
rect 2114 4138 2118 4141
rect 2118 4092 2121 4128
rect 2126 4072 2129 4248
rect 2134 4142 2137 4458
rect 2054 3422 2057 3658
rect 2062 3642 2065 3848
rect 2086 3762 2089 3868
rect 2086 3752 2089 3758
rect 2078 3722 2081 3738
rect 2070 3702 2073 3708
rect 2062 3602 2065 3638
rect 2054 3262 2057 3418
rect 2062 3362 2065 3538
rect 2074 3338 2078 3341
rect 2062 3282 2065 3298
rect 2086 3242 2089 3748
rect 2094 3702 2097 3828
rect 2102 3632 2105 3698
rect 2110 3692 2113 3778
rect 2126 3732 2129 4068
rect 2134 3982 2137 4068
rect 2134 3952 2137 3958
rect 2134 3892 2137 3928
rect 2142 3882 2145 4028
rect 2046 2702 2049 2838
rect 2070 2722 2073 3218
rect 2094 2822 2097 3338
rect 2102 3311 2105 3618
rect 2134 3482 2137 3868
rect 2130 3368 2134 3371
rect 2134 3352 2137 3358
rect 2122 3338 2126 3341
rect 2102 3308 2110 3311
rect 2102 3222 2105 3238
rect 2102 2811 2105 3218
rect 2114 3148 2118 3151
rect 2126 3102 2129 3108
rect 2098 2808 2105 2811
rect 2086 2762 2089 2808
rect 2046 2682 2049 2698
rect 2062 2682 2065 2688
rect 2050 2668 2054 2671
rect 2058 2658 2065 2661
rect 2054 2472 2057 2488
rect 2038 2201 2041 2308
rect 2046 2272 2049 2418
rect 2054 2372 2057 2398
rect 2062 2322 2065 2658
rect 2070 2382 2073 2698
rect 2078 2602 2081 2678
rect 2094 2632 2097 2808
rect 2102 2572 2105 2658
rect 2082 2558 2086 2561
rect 2082 2498 2086 2501
rect 2094 2492 2097 2568
rect 2102 2522 2105 2528
rect 2054 2282 2057 2288
rect 2062 2282 2065 2308
rect 2070 2272 2073 2348
rect 2070 2242 2073 2268
rect 2038 2198 2049 2201
rect 2030 1781 2033 2018
rect 2038 1872 2041 2028
rect 2038 1812 2041 1868
rect 2046 1782 2049 2198
rect 2054 2052 2057 2138
rect 2070 2112 2073 2168
rect 2054 1961 2057 2048
rect 2078 1962 2081 2458
rect 2086 2452 2089 2478
rect 2086 2412 2089 2438
rect 2094 2412 2097 2448
rect 2102 2362 2105 2478
rect 2110 2462 2113 2778
rect 2118 2662 2121 2668
rect 2118 2402 2121 2568
rect 2126 2532 2129 3078
rect 2134 3032 2137 3038
rect 2142 2982 2145 3878
rect 2150 3862 2153 4378
rect 2170 4148 2174 4151
rect 2166 3948 2174 3951
rect 2158 3722 2161 3728
rect 2166 3622 2169 3948
rect 2182 3932 2185 4728
rect 2190 4552 2193 4798
rect 2262 4312 2265 4808
rect 2350 4752 2353 4818
rect 2384 4803 2386 4807
rect 2390 4803 2393 4807
rect 2398 4803 2400 4807
rect 2198 4242 2201 4258
rect 2206 4252 2209 4268
rect 2194 4148 2198 4151
rect 2206 4002 2209 4168
rect 2190 3931 2193 3938
rect 2190 3928 2198 3931
rect 2150 3182 2153 3538
rect 2166 3362 2169 3548
rect 2182 3472 2185 3928
rect 2190 3682 2193 3928
rect 2206 3682 2209 3938
rect 2146 2888 2153 2891
rect 2150 2872 2153 2888
rect 2158 2882 2161 3088
rect 2142 2858 2150 2861
rect 2134 2572 2137 2808
rect 2142 2662 2145 2858
rect 2150 2682 2153 2748
rect 2150 2652 2153 2668
rect 2166 2662 2169 3348
rect 2158 2642 2161 2648
rect 2126 2462 2129 2468
rect 2094 2312 2097 2358
rect 2110 2212 2113 2328
rect 2086 2172 2089 2198
rect 2094 2012 2097 2148
rect 2102 2032 2105 2058
rect 2054 1958 2062 1961
rect 2082 1938 2086 1941
rect 2054 1892 2057 1898
rect 2062 1872 2065 1928
rect 2070 1862 2073 1888
rect 2094 1882 2097 1988
rect 2118 1982 2121 2358
rect 2134 2352 2137 2518
rect 2142 2452 2145 2458
rect 2126 2012 2129 2258
rect 2142 2252 2145 2438
rect 2110 1932 2113 1938
rect 2070 1792 2073 1808
rect 2030 1778 2038 1781
rect 2030 1752 2033 1778
rect 2042 1698 2049 1701
rect 2030 1352 2033 1698
rect 2046 1632 2049 1698
rect 2054 1562 2057 1688
rect 2070 1592 2073 1638
rect 2078 1522 2081 1868
rect 2102 1732 2105 1748
rect 2042 1498 2046 1501
rect 2022 942 2025 1248
rect 1782 252 1785 378
rect 1982 352 1985 388
rect 2014 362 2017 638
rect 2022 512 2025 918
rect 2030 802 2033 1348
rect 2046 1292 2049 1358
rect 2046 1192 2049 1288
rect 2062 1282 2065 1498
rect 2070 1342 2073 1428
rect 1778 148 1782 151
rect 1798 92 1801 338
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1886 303 1888 307
rect 1962 268 1966 271
rect 2030 252 2033 608
rect 2042 558 2046 561
rect 2054 542 2057 918
rect 2062 812 2065 1258
rect 2070 942 2073 1298
rect 2078 1192 2081 1468
rect 2086 1162 2089 1638
rect 2102 1492 2105 1588
rect 2110 1562 2113 1878
rect 2118 1812 2121 1978
rect 2118 1532 2121 1778
rect 2126 1652 2129 1948
rect 2134 1482 2137 1748
rect 2142 1622 2145 2248
rect 2150 1832 2153 2628
rect 2174 2612 2177 2948
rect 2182 2762 2185 3268
rect 2190 3202 2193 3668
rect 2182 2702 2185 2718
rect 2182 2672 2185 2678
rect 2174 2562 2177 2598
rect 2182 2562 2185 2588
rect 2158 2482 2161 2498
rect 2174 2492 2177 2498
rect 2158 2382 2161 2418
rect 2158 2222 2161 2268
rect 2162 2068 2166 2071
rect 2094 1282 2097 1348
rect 2094 1162 2097 1248
rect 2118 1122 2121 1148
rect 2070 742 2073 928
rect 2118 911 2121 1118
rect 2126 992 2129 1418
rect 2134 962 2137 1438
rect 2142 1142 2145 1238
rect 2142 1032 2145 1038
rect 2118 908 2126 911
rect 2070 662 2073 738
rect 2086 681 2089 788
rect 2086 678 2094 681
rect 2054 471 2057 538
rect 2110 518 2118 521
rect 2054 468 2062 471
rect 2110 412 2113 518
rect 2094 352 2097 378
rect 2126 372 2129 908
rect 1842 148 1846 151
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1886 103 1888 107
rect 1894 92 1897 108
rect 1918 62 1921 88
rect 2030 72 2033 248
rect 2038 162 2041 348
rect 2062 242 2065 338
rect 2126 232 2129 368
rect 2134 342 2137 948
rect 2150 882 2153 1798
rect 2158 862 2161 1968
rect 2166 1771 2169 1888
rect 2174 1832 2177 2348
rect 2182 2172 2185 2558
rect 2190 2322 2193 3198
rect 2206 3192 2209 3518
rect 2198 2912 2201 3088
rect 2198 2682 2201 2788
rect 2206 2782 2209 3188
rect 2198 2602 2201 2648
rect 2214 2642 2217 4188
rect 2238 4062 2241 4198
rect 2250 4138 2254 4141
rect 2222 3102 2225 3758
rect 2230 3652 2233 3918
rect 2230 2941 2233 3498
rect 2238 3362 2241 4058
rect 2262 3782 2265 4308
rect 2270 3722 2273 4298
rect 2258 3698 2265 3701
rect 2254 3582 2257 3628
rect 2262 3572 2265 3698
rect 2246 3492 2249 3558
rect 2246 3412 2249 3418
rect 2238 3142 2241 3148
rect 2230 2938 2241 2941
rect 2222 2692 2225 2708
rect 2206 2542 2209 2558
rect 2214 2542 2217 2618
rect 2198 2432 2201 2488
rect 2198 2312 2201 2428
rect 2174 1802 2177 1828
rect 2166 1768 2174 1771
rect 2174 1682 2177 1738
rect 2182 1662 2185 1988
rect 2190 1872 2193 2308
rect 2198 1772 2201 2258
rect 2206 2212 2209 2358
rect 2222 2312 2225 2608
rect 2230 2522 2233 2928
rect 2238 2682 2241 2938
rect 2246 2752 2249 3378
rect 2254 3302 2257 3318
rect 2254 2952 2257 3208
rect 2254 2872 2257 2938
rect 2262 2782 2265 3568
rect 2270 3292 2273 3298
rect 2270 3132 2273 3148
rect 2278 3142 2281 3148
rect 2278 2822 2281 3008
rect 2270 2782 2273 2818
rect 2238 2562 2241 2658
rect 2246 2612 2249 2738
rect 2254 2652 2257 2728
rect 2246 2572 2249 2608
rect 2206 2192 2209 2198
rect 2230 2162 2233 2368
rect 2238 2202 2241 2558
rect 2246 2232 2249 2338
rect 2254 2272 2257 2558
rect 2262 2532 2265 2738
rect 2262 2361 2265 2378
rect 2270 2372 2273 2668
rect 2278 2372 2281 2738
rect 2286 2702 2289 3588
rect 2294 2901 2297 3808
rect 2306 3758 2313 3761
rect 2310 3212 2313 3758
rect 2318 3492 2321 4128
rect 2326 4012 2329 4418
rect 2326 3962 2329 4008
rect 2326 3922 2329 3938
rect 2326 3512 2329 3918
rect 2334 3892 2337 4568
rect 2350 4522 2353 4748
rect 2358 4572 2361 4778
rect 2342 3852 2345 4458
rect 2350 4152 2353 4518
rect 2366 4271 2369 4578
rect 2362 4268 2369 4271
rect 2374 4082 2377 4698
rect 2384 4603 2386 4607
rect 2390 4603 2393 4607
rect 2398 4603 2400 4607
rect 2406 4482 2409 4868
rect 2438 4812 2441 5018
rect 2422 4732 2425 4788
rect 2422 4672 2425 4728
rect 2384 4403 2386 4407
rect 2390 4403 2393 4407
rect 2398 4403 2400 4407
rect 2414 4371 2417 4548
rect 2414 4368 2422 4371
rect 2384 4203 2386 4207
rect 2390 4203 2393 4207
rect 2398 4203 2400 4207
rect 2384 4003 2386 4007
rect 2390 4003 2393 4007
rect 2398 4003 2400 4007
rect 2342 3552 2345 3628
rect 2318 3332 2321 3428
rect 2310 3042 2313 3138
rect 2302 2922 2305 2968
rect 2294 2898 2305 2901
rect 2286 2462 2289 2678
rect 2262 2358 2270 2361
rect 2278 2302 2281 2318
rect 2206 1832 2209 2158
rect 2214 2002 2217 2108
rect 2230 2082 2233 2098
rect 2166 1472 2169 1578
rect 2182 1492 2185 1658
rect 2166 1162 2169 1188
rect 2166 1132 2169 1158
rect 2150 382 2153 738
rect 2158 542 2161 548
rect 2166 522 2169 1108
rect 2174 912 2177 1128
rect 2174 542 2177 888
rect 2186 698 2190 701
rect 2198 582 2201 1498
rect 2214 1382 2217 1898
rect 2222 1452 2225 2068
rect 2230 1852 2233 1868
rect 2238 1772 2241 1968
rect 2246 1762 2249 2158
rect 2254 2032 2257 2258
rect 2262 1982 2265 2198
rect 2270 2182 2273 2278
rect 2286 2212 2289 2228
rect 2270 2122 2273 2138
rect 2254 1932 2257 1958
rect 2262 1952 2265 1958
rect 2230 1352 2233 1378
rect 2230 1341 2233 1348
rect 2226 1338 2233 1341
rect 2214 662 2217 878
rect 2150 262 2153 378
rect 2150 152 2153 258
rect 2086 102 2089 128
rect 2222 12 2225 1148
rect 2238 762 2241 1368
rect 2254 1152 2257 1818
rect 2270 1742 2273 2078
rect 2278 1902 2281 2198
rect 2294 2152 2297 2888
rect 2302 2872 2305 2898
rect 2310 2842 2313 2968
rect 2302 2512 2305 2778
rect 2310 2632 2313 2658
rect 2302 2272 2305 2508
rect 2318 2451 2321 3318
rect 2334 3311 2337 3498
rect 2330 3308 2337 3311
rect 2342 3312 2345 3548
rect 2350 3532 2353 3728
rect 2342 2892 2345 3118
rect 2334 2662 2337 2798
rect 2334 2462 2337 2638
rect 2350 2512 2353 3128
rect 2358 3072 2361 3848
rect 2384 3803 2386 3807
rect 2390 3803 2393 3807
rect 2398 3803 2400 3807
rect 2394 3788 2398 3791
rect 2366 3412 2369 3768
rect 2406 3752 2409 3868
rect 2414 3692 2417 4348
rect 2438 4232 2441 4428
rect 2446 4342 2449 4378
rect 2438 3952 2441 4148
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2398 3603 2400 3607
rect 2358 2992 2361 3068
rect 2366 2992 2369 2998
rect 2318 2448 2326 2451
rect 2326 2412 2329 2448
rect 2342 2442 2345 2508
rect 2358 2472 2361 2948
rect 2366 2462 2369 2778
rect 2374 2492 2377 3488
rect 2406 3412 2409 3538
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2398 3403 2400 3407
rect 2406 3382 2409 3408
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2398 3203 2400 3207
rect 2406 3162 2409 3208
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2398 3003 2400 3007
rect 2406 2812 2409 3158
rect 2414 2952 2417 3678
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2398 2803 2400 2807
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2398 2603 2400 2607
rect 2402 2558 2406 2561
rect 2382 2482 2385 2528
rect 2310 2261 2313 2378
rect 2358 2342 2361 2428
rect 2322 2328 2326 2331
rect 2302 2258 2313 2261
rect 2302 2172 2305 2258
rect 2318 2251 2321 2308
rect 2310 2248 2321 2251
rect 2342 2252 2345 2308
rect 2350 2252 2353 2268
rect 2290 2138 2294 2141
rect 2294 2052 2297 2108
rect 2286 1822 2289 1888
rect 2282 1708 2289 1711
rect 2266 1598 2270 1601
rect 2270 1412 2273 1438
rect 2286 1402 2289 1708
rect 2294 1482 2297 2018
rect 2262 1332 2265 1388
rect 2302 1252 2305 2148
rect 2310 1412 2313 2248
rect 2318 2112 2321 2228
rect 2318 1812 2321 2008
rect 2326 1912 2329 2178
rect 2334 2132 2337 2168
rect 2342 2142 2345 2178
rect 2326 1882 2329 1888
rect 2334 1861 2337 1898
rect 2330 1858 2337 1861
rect 2342 1372 2345 2028
rect 2350 1652 2353 2248
rect 2358 2232 2361 2278
rect 2366 2242 2369 2388
rect 2374 2222 2377 2458
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2398 2403 2400 2407
rect 2406 2262 2409 2348
rect 2358 2042 2361 2208
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2398 2203 2400 2207
rect 2374 2192 2377 2198
rect 2370 2128 2374 2131
rect 2358 1842 2361 1938
rect 2278 1171 2281 1188
rect 2274 1168 2281 1171
rect 2262 952 2265 958
rect 2298 948 2302 951
rect 2238 752 2241 758
rect 2246 712 2249 868
rect 2246 672 2249 708
rect 2234 558 2241 561
rect 2238 552 2241 558
rect 2246 362 2249 658
rect 2254 572 2257 888
rect 2310 792 2313 1328
rect 2318 1162 2321 1268
rect 2318 872 2321 918
rect 2326 902 2329 1318
rect 2334 1112 2337 1328
rect 2310 762 2313 788
rect 2318 762 2321 768
rect 2246 292 2249 358
rect 2286 332 2289 738
rect 2334 672 2337 958
rect 2350 762 2353 1648
rect 2358 662 2361 1558
rect 2366 1152 2369 2068
rect 2374 1612 2377 2108
rect 2406 2102 2409 2208
rect 2414 2062 2417 2908
rect 2422 2581 2425 3878
rect 2430 2882 2433 3948
rect 2438 3762 2441 3928
rect 2446 3842 2449 4198
rect 2454 4192 2457 4878
rect 2482 4748 2486 4751
rect 2462 4428 2470 4431
rect 2462 4292 2465 4428
rect 2470 4272 2473 4278
rect 2478 4272 2481 4708
rect 2558 4372 2561 4848
rect 2566 4462 2569 4808
rect 2454 4072 2457 4168
rect 2442 3738 2449 3741
rect 2446 3712 2449 3738
rect 2438 3662 2441 3678
rect 2442 3648 2446 3651
rect 2438 3352 2441 3358
rect 2442 3278 2446 3281
rect 2442 3158 2446 3161
rect 2462 2992 2465 3868
rect 2470 3202 2473 4038
rect 2486 3742 2489 4238
rect 2494 3972 2497 4238
rect 2510 4132 2513 4278
rect 2502 3801 2505 4078
rect 2510 4012 2513 4128
rect 2518 3842 2521 4338
rect 2502 3798 2510 3801
rect 2494 3742 2497 3778
rect 2478 3262 2481 3568
rect 2502 3512 2505 3568
rect 2478 3132 2481 3248
rect 2486 3172 2489 3288
rect 2486 3162 2489 3168
rect 2494 3102 2497 3258
rect 2486 3082 2489 3098
rect 2486 3042 2489 3068
rect 2462 2818 2470 2821
rect 2422 2578 2433 2581
rect 2422 2562 2425 2568
rect 2422 2252 2425 2538
rect 2430 2352 2433 2578
rect 2438 2552 2441 2568
rect 2446 2481 2449 2738
rect 2438 2478 2449 2481
rect 2438 2422 2441 2478
rect 2446 2462 2449 2468
rect 2454 2452 2457 2788
rect 2462 2782 2465 2818
rect 2478 2772 2481 2958
rect 2486 2932 2489 2958
rect 2462 2452 2465 2458
rect 2438 2408 2446 2411
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2398 2003 2400 2007
rect 2406 1962 2409 2048
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2398 1803 2400 1807
rect 2414 1642 2417 1968
rect 2422 1832 2425 2238
rect 2406 1612 2409 1638
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2398 1603 2400 1607
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2398 1403 2400 1407
rect 2406 1341 2409 1438
rect 2414 1362 2417 1638
rect 2430 1602 2433 2098
rect 2438 1931 2441 2408
rect 2478 2392 2481 2698
rect 2486 2282 2489 2928
rect 2494 2752 2497 3098
rect 2502 3052 2505 3378
rect 2510 3062 2513 3538
rect 2502 2952 2505 2978
rect 2502 2812 2505 2948
rect 2494 2372 2497 2448
rect 2502 2372 2505 2798
rect 2510 2702 2513 3058
rect 2518 2962 2521 3348
rect 2526 3072 2529 3758
rect 2518 2682 2521 2708
rect 2510 2462 2513 2608
rect 2518 2462 2521 2678
rect 2526 2372 2529 3048
rect 2534 2942 2537 4258
rect 2542 3272 2545 4038
rect 2550 3272 2553 4018
rect 2550 3212 2553 3268
rect 2542 3052 2545 3198
rect 2534 2592 2537 2808
rect 2542 2742 2545 3048
rect 2474 2268 2478 2271
rect 2450 2258 2454 2261
rect 2462 2242 2465 2258
rect 2438 1928 2449 1931
rect 2438 1622 2441 1918
rect 2446 1802 2449 1928
rect 2454 1872 2457 2238
rect 2478 2122 2481 2158
rect 2466 2078 2470 2081
rect 2478 1972 2481 1978
rect 2486 1902 2489 2178
rect 2462 1888 2470 1891
rect 2462 1882 2465 1888
rect 2486 1862 2489 1888
rect 2486 1682 2489 1758
rect 2486 1662 2489 1668
rect 2406 1338 2414 1341
rect 2406 1282 2409 1328
rect 2446 1322 2449 1488
rect 2454 1482 2457 1548
rect 2454 1462 2457 1468
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2398 1203 2400 1207
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2398 1003 2400 1007
rect 2406 932 2409 1258
rect 2422 1082 2425 1208
rect 2414 882 2417 998
rect 2422 942 2425 958
rect 2414 862 2417 878
rect 2374 842 2377 858
rect 2334 472 2337 648
rect 2358 632 2361 658
rect 2374 552 2377 838
rect 2414 808 2422 811
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2398 803 2400 807
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2398 603 2400 607
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2398 403 2400 407
rect 2406 341 2409 668
rect 2414 362 2417 808
rect 2446 502 2449 1138
rect 2454 782 2457 1258
rect 2462 852 2465 1448
rect 2470 1402 2473 1588
rect 2486 1542 2489 1648
rect 2486 1272 2489 1538
rect 2482 1258 2486 1261
rect 2478 1162 2481 1198
rect 2478 1152 2481 1158
rect 2494 882 2497 2138
rect 2502 2072 2505 2368
rect 2510 2292 2513 2338
rect 2502 1902 2505 1948
rect 2502 1852 2505 1878
rect 2510 1762 2513 2188
rect 2518 2062 2521 2358
rect 2526 2172 2529 2318
rect 2534 2242 2537 2438
rect 2542 2422 2545 2458
rect 2542 2302 2545 2348
rect 2534 2202 2537 2218
rect 2526 2122 2529 2168
rect 2518 1872 2521 2018
rect 2518 1842 2521 1848
rect 2510 1572 2513 1718
rect 2518 1532 2521 1708
rect 2518 1352 2521 1358
rect 2502 1292 2505 1308
rect 2518 1262 2521 1278
rect 2478 572 2481 848
rect 2486 842 2489 858
rect 2494 822 2497 878
rect 2486 572 2489 738
rect 2478 562 2481 568
rect 2518 432 2521 878
rect 2526 482 2529 2038
rect 2534 1752 2537 2188
rect 2542 2142 2545 2298
rect 2550 2192 2553 3148
rect 2558 3122 2561 4368
rect 2574 4332 2577 4398
rect 2566 4222 2569 4258
rect 2574 4102 2577 4288
rect 2582 4162 2585 4888
rect 2630 4842 2633 4958
rect 2598 4472 2601 4728
rect 2566 3292 2569 3618
rect 2574 3562 2577 3568
rect 2574 3151 2577 3558
rect 2582 3301 2585 4108
rect 2590 3712 2593 4288
rect 2606 4062 2609 4748
rect 2638 4282 2641 4518
rect 2614 4142 2617 4148
rect 2614 3892 2617 4098
rect 2606 3612 2609 3618
rect 2590 3542 2593 3548
rect 2598 3312 2601 3448
rect 2582 3298 2593 3301
rect 2566 3148 2577 3151
rect 2558 3012 2561 3068
rect 2558 2562 2561 2938
rect 2566 2632 2569 3148
rect 2574 2902 2577 2948
rect 2582 2942 2585 2978
rect 2582 2862 2585 2888
rect 2590 2731 2593 3298
rect 2598 3062 2601 3108
rect 2606 2932 2609 3588
rect 2638 3372 2641 3388
rect 2618 3338 2622 3341
rect 2586 2728 2593 2731
rect 2566 2572 2569 2628
rect 2574 2612 2577 2728
rect 2590 2722 2593 2728
rect 2582 2612 2585 2708
rect 2558 2482 2561 2538
rect 2558 2462 2561 2478
rect 2558 2402 2561 2408
rect 2566 2271 2569 2548
rect 2574 2292 2577 2388
rect 2566 2268 2574 2271
rect 2558 2232 2561 2248
rect 2542 1851 2545 1968
rect 2550 1952 2553 2168
rect 2542 1848 2550 1851
rect 2542 1722 2545 1788
rect 2534 1662 2537 1668
rect 2558 1512 2561 1878
rect 2566 1822 2569 2258
rect 2574 2242 2577 2258
rect 2574 2032 2577 2188
rect 2590 2172 2593 2698
rect 2598 2632 2601 2928
rect 2606 2862 2609 2898
rect 2614 2732 2617 3318
rect 2622 3142 2625 3158
rect 2606 2692 2609 2718
rect 2614 2702 2617 2708
rect 2622 2622 2625 3098
rect 2630 3072 2633 3138
rect 2646 3112 2649 4128
rect 2654 3712 2657 4758
rect 2662 4512 2665 4718
rect 2654 3692 2657 3698
rect 2662 3682 2665 4448
rect 2686 4442 2689 4458
rect 2670 3872 2673 4108
rect 2686 4012 2689 4428
rect 2682 3868 2686 3871
rect 2670 3822 2673 3868
rect 2654 3152 2657 3198
rect 2630 2862 2633 3068
rect 2646 3022 2649 3108
rect 2654 3062 2657 3128
rect 2646 2831 2649 3018
rect 2654 2912 2657 3008
rect 2662 3002 2665 3638
rect 2670 3582 2673 3818
rect 2686 3662 2689 3678
rect 2682 3638 2686 3641
rect 2670 3372 2673 3498
rect 2670 2962 2673 3348
rect 2678 3232 2681 3548
rect 2686 3242 2689 3468
rect 2694 3402 2697 4608
rect 2726 4352 2729 4868
rect 2750 4672 2753 5088
rect 4498 5078 4502 5081
rect 4486 5072 4489 5078
rect 4578 5058 4582 5061
rect 2888 4903 2890 4907
rect 2894 4903 2897 4907
rect 2902 4903 2904 4907
rect 2878 4752 2881 4898
rect 3262 4851 3265 4858
rect 3258 4848 3265 4851
rect 2930 4838 2937 4841
rect 2858 4728 2862 4731
rect 2846 4642 2849 4718
rect 2870 4662 2873 4738
rect 2882 4728 2886 4731
rect 2888 4703 2890 4707
rect 2894 4703 2897 4707
rect 2902 4703 2904 4707
rect 2902 4672 2905 4678
rect 2934 4662 2937 4838
rect 3058 4748 3065 4751
rect 2734 4542 2737 4588
rect 2726 4272 2729 4338
rect 2718 3912 2721 4128
rect 2734 4042 2737 4528
rect 2742 4122 2745 4628
rect 2790 4552 2793 4558
rect 2710 3732 2713 3738
rect 2710 3702 2713 3708
rect 2726 3562 2729 3698
rect 2742 3612 2745 3868
rect 2710 3482 2713 3538
rect 2726 3492 2729 3558
rect 2678 3142 2681 3178
rect 2670 2942 2673 2958
rect 2654 2882 2657 2908
rect 2658 2858 2662 2861
rect 2638 2828 2649 2831
rect 2574 1942 2577 1968
rect 2582 1952 2585 2098
rect 2566 1782 2569 1818
rect 2574 1742 2577 1938
rect 2582 1892 2585 1948
rect 2586 1858 2590 1861
rect 2546 1458 2550 1461
rect 2550 1401 2553 1418
rect 2546 1398 2553 1401
rect 2538 1358 2542 1361
rect 2538 1258 2542 1261
rect 2550 1222 2553 1338
rect 2558 982 2561 1348
rect 2566 1152 2569 1698
rect 2574 1351 2577 1508
rect 2582 1432 2585 1738
rect 2574 1348 2582 1351
rect 2574 1172 2577 1288
rect 2574 562 2577 1058
rect 2582 992 2585 1178
rect 2526 452 2529 478
rect 2590 352 2593 1478
rect 2598 1182 2601 2588
rect 2618 2358 2622 2361
rect 2610 2168 2614 2171
rect 2606 1772 2609 2168
rect 2598 1132 2601 1148
rect 2606 862 2609 1688
rect 2614 1122 2617 1718
rect 2622 1662 2625 2158
rect 2630 2032 2633 2498
rect 2638 2232 2641 2828
rect 2654 2522 2657 2818
rect 2670 2811 2673 2938
rect 2666 2808 2673 2811
rect 2678 2812 2681 2828
rect 2686 2822 2689 3118
rect 2694 2932 2697 3178
rect 2702 3092 2705 3448
rect 2710 3332 2713 3478
rect 2710 3322 2713 3328
rect 2734 3322 2737 3608
rect 2750 3351 2753 4488
rect 2758 3662 2761 4498
rect 2766 4132 2769 4228
rect 2774 4192 2777 4358
rect 2798 4342 2801 4618
rect 2782 4142 2785 4178
rect 2766 3672 2769 4128
rect 2782 3732 2785 3748
rect 2742 3348 2753 3351
rect 2742 3312 2745 3348
rect 2758 3341 2761 3608
rect 2750 3338 2761 3341
rect 2718 3232 2721 3278
rect 2702 2772 2705 2798
rect 2662 2472 2665 2478
rect 2654 2361 2657 2378
rect 2650 2358 2657 2361
rect 2662 2292 2665 2418
rect 2670 2332 2673 2518
rect 2670 2312 2673 2328
rect 2646 2262 2649 2268
rect 2658 2258 2662 2261
rect 2670 2112 2673 2288
rect 2630 1912 2633 1928
rect 2630 1792 2633 1808
rect 2622 1622 2625 1658
rect 2622 1222 2625 1478
rect 2638 1392 2641 2068
rect 2678 2002 2681 2698
rect 2694 2462 2697 2508
rect 2690 2398 2694 2401
rect 2686 2252 2689 2298
rect 2694 2232 2697 2378
rect 2646 1722 2649 1998
rect 2678 1952 2681 1958
rect 2666 1938 2670 1941
rect 2646 1662 2649 1718
rect 2654 1612 2657 1878
rect 2666 1848 2670 1851
rect 2686 1832 2689 1998
rect 2662 1802 2665 1808
rect 2630 851 2633 1088
rect 2646 962 2649 1458
rect 2670 1202 2673 1708
rect 2678 1662 2681 1668
rect 2686 1252 2689 1828
rect 2694 1632 2697 2078
rect 2702 2062 2705 2768
rect 2710 2692 2713 3218
rect 2718 2542 2721 3018
rect 2718 2472 2721 2528
rect 2726 2522 2729 3278
rect 2734 3272 2737 3298
rect 2742 3262 2745 3268
rect 2734 2732 2737 3068
rect 2750 2942 2753 3338
rect 2758 3242 2761 3328
rect 2750 2902 2753 2918
rect 2758 2832 2761 3238
rect 2766 3232 2769 3498
rect 2774 3242 2777 3608
rect 2782 3282 2785 3698
rect 2790 3412 2793 3748
rect 2766 2852 2769 2948
rect 2726 2462 2729 2508
rect 2710 2292 2713 2458
rect 2726 2401 2729 2408
rect 2722 2398 2729 2401
rect 2718 2302 2721 2318
rect 2726 2252 2729 2258
rect 2714 2248 2718 2251
rect 2710 2052 2713 2058
rect 2734 2022 2737 2728
rect 2766 2622 2769 2848
rect 2782 2602 2785 3188
rect 2790 3052 2793 3398
rect 2798 3202 2801 4338
rect 2814 4262 2817 4548
rect 2826 4538 2830 4541
rect 2862 4522 2865 4528
rect 2838 4302 2841 4348
rect 2826 4278 2830 4281
rect 2814 4222 2817 4258
rect 2822 4112 2825 4138
rect 2806 3402 2809 3778
rect 2822 3732 2825 4018
rect 2830 3902 2833 4248
rect 2838 4192 2841 4298
rect 2854 4192 2857 4238
rect 2862 4232 2865 4268
rect 2814 3481 2817 3698
rect 2814 3478 2822 3481
rect 2830 3462 2833 3898
rect 2846 3861 2849 4088
rect 2854 4042 2857 4188
rect 2870 4032 2873 4658
rect 2954 4548 2958 4551
rect 2888 4503 2890 4507
rect 2894 4503 2897 4507
rect 2902 4503 2904 4507
rect 2854 3972 2857 4028
rect 2878 4012 2881 4328
rect 2888 4303 2890 4307
rect 2894 4303 2897 4307
rect 2902 4303 2904 4307
rect 2890 4278 2894 4281
rect 2888 4103 2890 4107
rect 2894 4103 2897 4107
rect 2902 4103 2904 4107
rect 2918 4042 2921 4238
rect 2926 4152 2929 4248
rect 2854 3951 2857 3968
rect 2854 3948 2862 3951
rect 2854 3932 2857 3938
rect 2846 3858 2854 3861
rect 2870 3842 2873 4008
rect 2838 3681 2841 3768
rect 2838 3678 2846 3681
rect 2838 3312 2841 3578
rect 2834 3288 2841 3291
rect 2838 3272 2841 3288
rect 2834 3248 2838 3251
rect 2794 2748 2798 2751
rect 2790 2642 2793 2738
rect 2806 2672 2809 3248
rect 2822 3162 2825 3168
rect 2838 3152 2841 3158
rect 2798 2652 2801 2658
rect 2822 2612 2825 3138
rect 2838 3082 2841 3108
rect 2830 3062 2833 3068
rect 2846 2832 2849 3638
rect 2854 3632 2857 3638
rect 2862 3532 2865 3728
rect 2854 3252 2857 3298
rect 2870 3162 2873 3838
rect 2878 3832 2881 3948
rect 2888 3903 2890 3907
rect 2894 3903 2897 3907
rect 2902 3903 2904 3907
rect 2878 3382 2881 3788
rect 2888 3703 2890 3707
rect 2894 3703 2897 3707
rect 2902 3703 2904 3707
rect 2910 3542 2913 3878
rect 2888 3503 2890 3507
rect 2894 3503 2897 3507
rect 2902 3503 2904 3507
rect 2910 3382 2913 3508
rect 2888 3303 2890 3307
rect 2894 3303 2897 3307
rect 2902 3303 2904 3307
rect 2898 3238 2905 3241
rect 2902 3232 2905 3238
rect 2910 3182 2913 3338
rect 2854 3122 2857 3128
rect 2758 2561 2761 2568
rect 2758 2558 2766 2561
rect 2742 2528 2750 2531
rect 2742 2432 2745 2528
rect 2754 2468 2758 2471
rect 2766 2462 2769 2558
rect 2782 2522 2785 2548
rect 2742 2252 2745 2428
rect 2766 2342 2769 2458
rect 2774 2232 2777 2518
rect 2790 2502 2793 2548
rect 2802 2508 2806 2511
rect 2782 2462 2785 2488
rect 2798 2411 2801 2488
rect 2794 2408 2801 2411
rect 2814 2372 2817 2428
rect 2790 2282 2793 2368
rect 2822 2352 2825 2548
rect 2838 2412 2841 2448
rect 2846 2342 2849 2458
rect 2806 2332 2809 2338
rect 2742 2228 2750 2231
rect 2742 2212 2745 2228
rect 2742 1962 2745 2208
rect 2754 2118 2758 2121
rect 2702 1352 2705 1938
rect 2718 1812 2721 1908
rect 2710 1782 2713 1808
rect 2714 1658 2718 1661
rect 2686 1172 2689 1248
rect 2686 1072 2689 1088
rect 2666 1068 2670 1071
rect 2702 1022 2705 1218
rect 2718 1132 2721 1248
rect 2726 1072 2729 1168
rect 2702 962 2705 1018
rect 2710 972 2713 978
rect 2646 872 2649 958
rect 2710 942 2713 948
rect 2630 848 2638 851
rect 2402 338 2409 341
rect 2330 248 2334 251
rect 2358 182 2361 308
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2398 203 2400 207
rect 2622 152 2625 738
rect 2710 682 2713 828
rect 2718 722 2721 1068
rect 2630 262 2633 508
rect 2630 202 2633 258
rect 2646 102 2649 518
rect 2654 382 2657 618
rect 2654 332 2657 378
rect 2662 192 2665 558
rect 2678 272 2681 478
rect 2662 152 2665 188
rect 2694 132 2697 668
rect 2726 662 2729 1058
rect 2734 1032 2737 1148
rect 2702 452 2705 658
rect 2742 632 2745 1938
rect 2750 1862 2753 2068
rect 2750 1772 2753 1778
rect 2758 1692 2761 2098
rect 2766 1932 2769 1968
rect 2774 1952 2777 1958
rect 2766 1882 2769 1918
rect 2758 1462 2761 1648
rect 2766 1002 2769 1418
rect 2774 1292 2777 1318
rect 2774 1242 2777 1278
rect 2782 1262 2785 2248
rect 2790 1932 2793 2278
rect 2798 1972 2801 2178
rect 2806 2082 2809 2298
rect 2846 2272 2849 2278
rect 2818 2258 2825 2261
rect 2822 2252 2825 2258
rect 2806 2011 2809 2068
rect 2806 2008 2814 2011
rect 2790 1592 2793 1858
rect 2790 1292 2793 1588
rect 2798 1542 2801 1588
rect 2798 1352 2801 1358
rect 2790 962 2793 988
rect 2758 822 2761 958
rect 2806 952 2809 1978
rect 2822 1892 2825 2188
rect 2814 1512 2817 1538
rect 2814 1132 2817 1268
rect 2778 938 2782 941
rect 2822 852 2825 1858
rect 2830 732 2833 2098
rect 2838 1522 2841 2198
rect 2854 2022 2857 3118
rect 2870 2832 2873 3158
rect 2888 3103 2890 3107
rect 2894 3103 2897 3107
rect 2902 3103 2904 3107
rect 2878 3072 2881 3098
rect 2910 2972 2913 3178
rect 2918 3102 2921 4038
rect 2926 3732 2929 4148
rect 2934 3852 2937 4118
rect 2934 3782 2937 3848
rect 2942 3732 2945 4488
rect 3062 4462 3065 4748
rect 3070 4652 3073 4748
rect 2950 4242 2953 4248
rect 2958 4242 2961 4248
rect 2950 3872 2953 3958
rect 2888 2903 2890 2907
rect 2894 2903 2897 2907
rect 2902 2903 2904 2907
rect 2910 2892 2913 2898
rect 2862 2412 2865 2448
rect 2862 2352 2865 2358
rect 2870 2152 2873 2758
rect 2878 2712 2881 2758
rect 2888 2703 2890 2707
rect 2894 2703 2897 2707
rect 2902 2703 2904 2707
rect 2878 2522 2881 2678
rect 2886 2532 2889 2618
rect 2898 2558 2902 2561
rect 2878 2482 2881 2518
rect 2888 2503 2890 2507
rect 2894 2503 2897 2507
rect 2902 2503 2904 2507
rect 2898 2428 2902 2431
rect 2890 2338 2894 2341
rect 2888 2303 2890 2307
rect 2894 2303 2897 2307
rect 2902 2303 2904 2307
rect 2910 2252 2913 2828
rect 2918 2492 2921 3028
rect 2926 2852 2929 3708
rect 2934 3652 2937 3668
rect 2942 3652 2945 3718
rect 2950 3662 2953 3868
rect 2934 3362 2937 3608
rect 2950 3562 2953 3658
rect 2942 3302 2945 3358
rect 2934 3102 2937 3148
rect 2942 3142 2945 3188
rect 2918 2272 2921 2308
rect 2846 1772 2849 1958
rect 2862 1852 2865 1918
rect 2870 1842 2873 1918
rect 2850 1678 2857 1681
rect 2854 1612 2857 1678
rect 2838 1212 2841 1518
rect 2862 1452 2865 1768
rect 2870 1732 2873 1838
rect 2870 1382 2873 1698
rect 2878 1622 2881 2218
rect 2888 2103 2890 2107
rect 2894 2103 2897 2107
rect 2902 2103 2904 2107
rect 2910 1942 2913 2118
rect 2918 1972 2921 2148
rect 2926 2102 2929 2568
rect 2934 2522 2937 3048
rect 2942 2892 2945 3098
rect 2942 2512 2945 2858
rect 2950 2622 2953 3178
rect 2958 2792 2961 4238
rect 2966 3692 2969 4288
rect 3010 4278 3017 4281
rect 3014 4232 3017 4278
rect 3022 4202 3025 4368
rect 3038 4152 3041 4158
rect 3034 4138 3038 4141
rect 2974 3632 2977 3678
rect 2982 3652 2985 3718
rect 2990 3702 2993 3718
rect 2966 3532 2969 3538
rect 2982 3472 2985 3638
rect 2966 3242 2969 3388
rect 2966 2802 2969 3238
rect 2958 2761 2961 2778
rect 2958 2758 2966 2761
rect 2958 2742 2961 2748
rect 2974 2732 2977 3368
rect 2982 2672 2985 3378
rect 2998 3142 3001 3698
rect 2990 3042 2993 3088
rect 2990 2942 2993 2948
rect 2998 2872 3001 2948
rect 3006 2922 3009 4128
rect 3014 4062 3017 4068
rect 3054 4032 3057 4068
rect 3042 3758 3046 3761
rect 3030 3672 3033 3678
rect 3046 3662 3049 3678
rect 3034 3658 3038 3661
rect 3030 3582 3033 3658
rect 3014 3322 3017 3418
rect 3006 2872 3009 2918
rect 2990 2792 2993 2838
rect 2998 2782 3001 2868
rect 3014 2802 3017 3318
rect 2950 2512 2953 2548
rect 2934 2452 2937 2458
rect 2942 2292 2945 2488
rect 2958 2432 2961 2648
rect 2990 2642 2993 2678
rect 2982 2552 2985 2558
rect 2990 2542 2993 2568
rect 2970 2458 2974 2461
rect 2950 2352 2953 2408
rect 2966 2341 2969 2398
rect 2974 2372 2977 2388
rect 2962 2338 2969 2341
rect 2950 2212 2953 2298
rect 2888 1903 2890 1907
rect 2894 1903 2897 1907
rect 2902 1903 2904 1907
rect 2886 1752 2889 1848
rect 2914 1838 2918 1841
rect 2888 1703 2890 1707
rect 2894 1703 2897 1707
rect 2902 1703 2904 1707
rect 2914 1688 2918 1691
rect 2918 1592 2921 1608
rect 2926 1602 2929 2038
rect 2942 1832 2945 2118
rect 2958 2082 2961 2088
rect 2982 2072 2985 2488
rect 2990 2342 2993 2538
rect 2990 2282 2993 2298
rect 2998 2282 3001 2778
rect 3022 2642 3025 3538
rect 3038 3352 3041 3408
rect 3054 3372 3057 4018
rect 3062 3412 3065 4448
rect 3070 3852 3073 4398
rect 3070 3822 3073 3838
rect 3038 3342 3041 3348
rect 3030 3152 3033 3158
rect 3038 3072 3041 3178
rect 3046 3032 3049 3148
rect 3054 3132 3057 3338
rect 3030 2982 3033 2998
rect 3038 2952 3041 3028
rect 3046 2972 3049 3028
rect 3030 2932 3033 2938
rect 3054 2912 3057 3028
rect 3062 2992 3065 3028
rect 3030 2702 3033 2888
rect 3070 2852 3073 3818
rect 3078 3732 3081 4178
rect 3086 4012 3089 4458
rect 3094 4062 3097 4498
rect 3118 4472 3121 4568
rect 3122 4458 3126 4461
rect 3126 4362 3129 4458
rect 3078 3192 3081 3728
rect 3086 3442 3089 3798
rect 3094 3782 3097 3838
rect 3102 3542 3105 3848
rect 3086 3072 3089 3438
rect 3094 3332 3097 3518
rect 3086 3062 3089 3068
rect 3010 2548 3014 2551
rect 3022 2512 3025 2548
rect 3030 2542 3033 2548
rect 3006 2432 3009 2508
rect 3014 2462 3017 2498
rect 3026 2488 3030 2491
rect 3006 2342 3009 2428
rect 3014 2272 3017 2358
rect 3030 2352 3033 2368
rect 3022 2332 3025 2338
rect 2998 2202 3001 2258
rect 3006 2102 3009 2108
rect 2958 1962 2961 2048
rect 2934 1752 2937 1758
rect 2918 1552 2921 1588
rect 2888 1503 2890 1507
rect 2894 1503 2897 1507
rect 2902 1503 2904 1507
rect 2910 1462 2913 1508
rect 2842 1178 2846 1181
rect 2854 922 2857 1338
rect 2888 1303 2890 1307
rect 2894 1303 2897 1307
rect 2902 1303 2904 1307
rect 2862 732 2865 1288
rect 2862 702 2865 728
rect 2750 652 2753 668
rect 2870 652 2873 1108
rect 2878 992 2881 1208
rect 2942 1162 2945 1828
rect 2950 1752 2953 1798
rect 2958 1652 2961 1958
rect 2950 1372 2953 1548
rect 2958 1302 2961 1638
rect 2966 1462 2969 2018
rect 2954 1258 2958 1261
rect 2910 1138 2918 1141
rect 2888 1103 2890 1107
rect 2894 1103 2897 1107
rect 2902 1103 2904 1107
rect 2888 903 2890 907
rect 2894 903 2897 907
rect 2902 903 2904 907
rect 2888 703 2890 707
rect 2894 703 2897 707
rect 2902 703 2904 707
rect 2910 622 2913 1138
rect 2946 1108 2950 1111
rect 2918 1062 2921 1098
rect 2918 762 2921 1058
rect 2942 1052 2945 1108
rect 2958 952 2961 1208
rect 2966 1022 2969 1348
rect 2926 842 2929 898
rect 2974 862 2977 1408
rect 2982 1342 2985 2068
rect 3022 2042 3025 2048
rect 3030 1972 3033 2278
rect 3038 2051 3041 2638
rect 3054 2602 3057 2728
rect 3062 2602 3065 2818
rect 3070 2782 3073 2808
rect 3086 2612 3089 3018
rect 3094 2602 3097 3328
rect 3102 3182 3105 3508
rect 3110 3442 3113 4138
rect 3118 4088 3126 4091
rect 3118 3872 3121 4088
rect 3150 3792 3153 4728
rect 3174 4272 3177 4278
rect 3118 3572 3121 3768
rect 3134 3732 3137 3778
rect 3146 3758 3153 3761
rect 3150 3752 3153 3758
rect 3110 3402 3113 3438
rect 3102 2812 3105 3178
rect 3110 2802 3113 3138
rect 3118 3052 3121 3568
rect 3126 3082 3129 3568
rect 3134 3272 3137 3668
rect 3150 3542 3153 3578
rect 3142 3442 3145 3458
rect 3150 3452 3153 3468
rect 3142 3212 3145 3438
rect 3158 3372 3161 4048
rect 3166 3651 3169 4268
rect 3182 4082 3185 4768
rect 3182 3952 3185 3978
rect 3174 3872 3177 3888
rect 3190 3762 3193 4708
rect 3230 4632 3233 4638
rect 3214 4472 3217 4558
rect 3206 4292 3209 4348
rect 3206 4272 3209 4288
rect 3198 4052 3201 4108
rect 3206 4012 3209 4268
rect 3210 3828 3214 3831
rect 3206 3712 3209 3758
rect 3214 3752 3217 3758
rect 3214 3652 3217 3658
rect 3166 3648 3174 3651
rect 3166 3542 3169 3618
rect 3166 3312 3169 3538
rect 3174 3472 3177 3478
rect 3102 2632 3105 2738
rect 3046 2472 3049 2498
rect 3046 2352 3049 2368
rect 3038 2048 3049 2051
rect 3022 1742 3025 1818
rect 3030 1812 3033 1818
rect 2998 1652 3001 1678
rect 3006 1512 3009 1658
rect 3014 1522 3017 1698
rect 3022 1572 3025 1708
rect 3030 1701 3033 1798
rect 3038 1762 3041 2038
rect 3046 1872 3049 2048
rect 3030 1698 3041 1701
rect 2998 1441 3001 1448
rect 2994 1438 3001 1441
rect 3006 1372 3009 1388
rect 3002 1348 3009 1351
rect 3006 1322 3009 1348
rect 2994 1258 2998 1261
rect 3014 1172 3017 1518
rect 3022 1502 3025 1518
rect 3022 1162 3025 1338
rect 3030 1212 3033 1588
rect 3038 1502 3041 1698
rect 3030 1162 3033 1168
rect 3038 1162 3041 1228
rect 3018 1138 3022 1141
rect 3030 1122 3033 1128
rect 2886 552 2889 558
rect 2888 503 2890 507
rect 2894 503 2897 507
rect 2902 503 2904 507
rect 2702 392 2705 448
rect 2702 372 2705 388
rect 2718 262 2721 398
rect 2726 262 2729 498
rect 2734 272 2737 498
rect 2782 462 2785 468
rect 2870 452 2873 458
rect 2888 303 2890 307
rect 2894 303 2897 307
rect 2902 303 2904 307
rect 2918 272 2921 598
rect 2926 492 2929 798
rect 2974 722 2977 728
rect 2982 692 2985 1118
rect 2990 872 2993 1068
rect 2990 862 2993 868
rect 2990 842 2993 848
rect 2998 802 3001 928
rect 3030 812 3033 888
rect 3038 882 3041 1158
rect 3046 982 3049 1828
rect 3054 1362 3057 2598
rect 3062 2432 3065 2578
rect 3070 2562 3073 2588
rect 3078 2542 3081 2558
rect 3086 2542 3089 2548
rect 3094 2532 3097 2598
rect 3102 2542 3105 2548
rect 3062 2362 3065 2408
rect 3078 2392 3081 2478
rect 3098 2398 3102 2401
rect 3062 2352 3065 2358
rect 3074 2118 3081 2121
rect 3062 2052 3065 2118
rect 3078 2112 3081 2118
rect 3070 1802 3073 2038
rect 3078 1952 3081 1978
rect 3078 1672 3081 1818
rect 3094 1632 3097 2348
rect 3110 2342 3113 2798
rect 3118 2362 3121 2818
rect 3134 2712 3137 3198
rect 3150 3122 3153 3148
rect 3142 3048 3150 3051
rect 3142 2982 3145 3048
rect 3142 2852 3145 2968
rect 3150 2742 3153 3028
rect 3146 2698 3150 2701
rect 3126 2272 3129 2538
rect 3134 2512 3137 2528
rect 3150 2432 3153 2438
rect 3134 2322 3137 2328
rect 3142 2322 3145 2398
rect 3134 2262 3137 2268
rect 3150 2092 3153 2428
rect 3102 1702 3105 2008
rect 3142 1852 3145 2088
rect 3150 1852 3153 1868
rect 3142 1832 3145 1848
rect 3110 1782 3113 1818
rect 3062 1422 3065 1508
rect 3070 1212 3073 1598
rect 3078 1382 3081 1538
rect 3086 1532 3089 1538
rect 3070 892 3073 1078
rect 3022 762 3025 768
rect 3026 758 3030 761
rect 2990 732 2993 748
rect 3038 722 3041 748
rect 2926 462 2929 488
rect 3006 452 3009 458
rect 3014 442 3017 718
rect 3046 682 3049 838
rect 3054 742 3057 818
rect 3062 652 3065 858
rect 3078 822 3081 868
rect 3086 862 3089 1388
rect 3094 1232 3097 1568
rect 3102 1542 3105 1698
rect 3110 1652 3113 1658
rect 3118 1562 3121 1748
rect 3142 1672 3145 1738
rect 3150 1692 3153 1698
rect 3142 1612 3145 1668
rect 3150 1662 3153 1668
rect 3114 1538 3118 1541
rect 3102 1452 3105 1538
rect 3110 1442 3113 1458
rect 3038 562 3041 628
rect 3086 532 3089 858
rect 3094 672 3097 878
rect 3102 702 3105 1438
rect 3110 1152 3113 1158
rect 3118 952 3121 1448
rect 3126 1282 3129 1298
rect 3134 1272 3137 1298
rect 3134 762 3137 1138
rect 3142 932 3145 1528
rect 3150 1222 3153 1638
rect 3158 1352 3161 3178
rect 3166 2832 3169 3128
rect 3174 3102 3177 3408
rect 3182 3122 3185 3468
rect 3190 3232 3193 3588
rect 3214 3541 3217 3608
rect 3210 3538 3217 3541
rect 3222 3592 3225 4448
rect 3230 3932 3233 4628
rect 3198 3522 3201 3528
rect 3206 3482 3209 3498
rect 3202 3458 3209 3461
rect 3206 3452 3209 3458
rect 3214 3402 3217 3518
rect 3214 3332 3217 3368
rect 3198 3152 3201 3168
rect 3174 2982 3177 3098
rect 3174 2972 3177 2978
rect 3198 2922 3201 3008
rect 3206 2982 3209 2988
rect 3198 2871 3201 2918
rect 3198 2868 3206 2871
rect 3166 2752 3169 2758
rect 3166 2542 3169 2738
rect 3174 2522 3177 2858
rect 3190 2842 3193 2848
rect 3166 2462 3169 2518
rect 3166 2352 3169 2378
rect 3174 2182 3177 2518
rect 3182 2462 3185 2468
rect 3190 2441 3193 2838
rect 3214 2592 3217 3328
rect 3222 2732 3225 3588
rect 3230 3542 3233 3888
rect 3238 3672 3241 4168
rect 3254 4132 3257 4438
rect 3262 4412 3265 4848
rect 3278 4662 3281 5048
rect 3400 5003 3402 5007
rect 3406 5003 3409 5007
rect 3414 5003 3416 5007
rect 3558 5002 3561 5048
rect 3400 4803 3402 4807
rect 3406 4803 3409 4807
rect 3414 4803 3416 4807
rect 3422 4772 3425 4818
rect 3270 4312 3273 4658
rect 3270 4262 3273 4308
rect 3286 4152 3289 4548
rect 3342 4542 3345 4688
rect 3358 4552 3361 4738
rect 3370 4668 3374 4671
rect 3400 4603 3402 4607
rect 3406 4603 3409 4607
rect 3414 4603 3416 4607
rect 3400 4403 3402 4407
rect 3406 4403 3409 4407
rect 3414 4403 3416 4407
rect 3338 4348 3342 4351
rect 3402 4348 3406 4351
rect 3286 4132 3289 4148
rect 3298 3858 3302 3861
rect 3270 3822 3273 3848
rect 3262 3742 3265 3758
rect 3254 3542 3257 3628
rect 3230 3432 3233 3448
rect 3230 2922 3233 3398
rect 3238 3082 3241 3498
rect 3262 3312 3265 3738
rect 3270 3671 3273 3818
rect 3270 3668 3278 3671
rect 3294 3632 3297 3728
rect 3278 3482 3281 3578
rect 3294 3562 3297 3628
rect 3254 2962 3257 2988
rect 3262 2852 3265 3068
rect 3246 2702 3249 2848
rect 3222 2592 3225 2628
rect 3198 2471 3201 2488
rect 3198 2468 3206 2471
rect 3222 2462 3225 2498
rect 3238 2482 3241 2618
rect 3246 2552 3249 2608
rect 3182 2438 3193 2441
rect 3166 1792 3169 2118
rect 3150 1082 3153 1118
rect 3142 922 3145 928
rect 3126 562 3129 668
rect 3158 532 3161 1308
rect 3166 1292 3169 1688
rect 3166 962 3169 1168
rect 3174 1012 3177 2078
rect 3182 1901 3185 2438
rect 3190 2402 3193 2428
rect 3222 2362 3225 2418
rect 3190 2312 3193 2348
rect 3198 2122 3201 2338
rect 3214 2292 3217 2328
rect 3230 2302 3233 2478
rect 3242 2448 3246 2451
rect 3222 2292 3225 2298
rect 3254 2271 3257 2558
rect 3254 2268 3262 2271
rect 3206 2252 3209 2268
rect 3206 2212 3209 2248
rect 3222 2052 3225 2138
rect 3230 2002 3233 2258
rect 3238 2158 3246 2161
rect 3238 2052 3241 2158
rect 3254 2122 3257 2178
rect 3262 2162 3265 2218
rect 3182 1898 3190 1901
rect 3182 1882 3185 1898
rect 3182 1202 3185 1768
rect 3166 682 3169 958
rect 3174 952 3177 1008
rect 3182 882 3185 1138
rect 3190 922 3193 1828
rect 3198 1732 3201 1928
rect 3074 508 3081 511
rect 3022 488 3030 491
rect 2934 142 2937 288
rect 3022 242 3025 488
rect 3078 472 3081 508
rect 3054 381 3057 388
rect 3050 378 3057 381
rect 3110 152 3113 438
rect 3158 362 3161 528
rect 3166 192 3169 638
rect 3198 552 3201 1728
rect 3206 582 3209 1978
rect 3214 1848 3222 1851
rect 3214 1662 3217 1848
rect 3238 1692 3241 1968
rect 3222 1662 3225 1668
rect 3214 1072 3217 1398
rect 3222 1262 3225 1278
rect 3230 1182 3233 1688
rect 3238 1672 3241 1678
rect 3238 1202 3241 1318
rect 3246 1262 3249 1728
rect 3254 1452 3257 1998
rect 3270 1952 3273 2508
rect 3278 2492 3281 3348
rect 3286 3002 3289 3538
rect 3294 3281 3297 3558
rect 3302 3422 3305 3858
rect 3310 3682 3313 4048
rect 3310 3572 3313 3658
rect 3318 3552 3321 4158
rect 3334 3692 3337 4328
rect 3386 4318 3393 4321
rect 3390 4302 3393 4318
rect 3342 3812 3345 4078
rect 3382 3992 3385 4228
rect 3374 3901 3377 3948
rect 3382 3942 3385 3988
rect 3390 3962 3393 4298
rect 3400 4203 3402 4207
rect 3406 4203 3409 4207
rect 3414 4203 3416 4207
rect 3400 4003 3402 4007
rect 3406 4003 3409 4007
rect 3414 4003 3416 4007
rect 3398 3922 3401 3938
rect 3374 3898 3382 3901
rect 3378 3848 3385 3851
rect 3382 3822 3385 3848
rect 3386 3818 3393 3821
rect 3378 3748 3382 3751
rect 3294 3278 3302 3281
rect 3298 3268 3302 3271
rect 3302 3042 3305 3238
rect 3302 3012 3305 3038
rect 3286 2752 3289 2788
rect 3294 2532 3297 2918
rect 3302 2622 3305 2998
rect 3310 2972 3313 3518
rect 3318 2652 3321 3518
rect 3326 2912 3329 3628
rect 3334 3292 3337 3688
rect 3334 3042 3337 3048
rect 3326 2762 3329 2908
rect 3334 2832 3337 3038
rect 3286 2472 3289 2488
rect 3278 1992 3281 2208
rect 3286 2142 3289 2148
rect 3286 2052 3289 2058
rect 3278 1962 3281 1988
rect 3266 1938 3270 1941
rect 3262 1752 3265 1938
rect 3278 1582 3281 1898
rect 3262 1482 3265 1538
rect 3270 1242 3273 1548
rect 3278 1481 3281 1578
rect 3286 1502 3289 2038
rect 3294 1882 3297 2518
rect 3326 2512 3329 2688
rect 3334 2532 3337 2828
rect 3302 2202 3305 2498
rect 3310 2452 3313 2508
rect 3342 2502 3345 3728
rect 3358 3712 3361 3738
rect 3350 3672 3353 3678
rect 3358 3342 3361 3708
rect 3366 3662 3369 3748
rect 3366 3482 3369 3658
rect 3350 3272 3353 3278
rect 3350 2522 3353 2978
rect 3358 2912 3361 3028
rect 3366 2842 3369 3478
rect 3382 3372 3385 3528
rect 3390 3332 3393 3818
rect 3400 3803 3402 3807
rect 3406 3803 3409 3807
rect 3414 3803 3416 3807
rect 3422 3642 3425 4768
rect 3430 4542 3433 4878
rect 3438 4702 3441 4838
rect 3526 4712 3529 4868
rect 3438 4062 3441 4698
rect 3550 4652 3553 4988
rect 3462 4532 3465 4538
rect 3454 4242 3457 4448
rect 3454 4122 3457 4218
rect 3430 3872 3433 3878
rect 3400 3603 3402 3607
rect 3406 3603 3409 3607
rect 3414 3603 3416 3607
rect 3438 3552 3441 3778
rect 3446 3612 3449 3838
rect 3454 3702 3457 4118
rect 3462 3832 3465 4528
rect 3470 4002 3473 4528
rect 3462 3762 3465 3808
rect 3442 3528 3446 3531
rect 3400 3403 3402 3407
rect 3406 3403 3409 3407
rect 3414 3403 3416 3407
rect 3374 3202 3377 3298
rect 3400 3203 3402 3207
rect 3406 3203 3409 3207
rect 3414 3203 3416 3207
rect 3358 2712 3361 2738
rect 3338 2468 3342 2471
rect 3326 2462 3329 2468
rect 3334 2412 3337 2468
rect 3342 2392 3345 2438
rect 3314 2378 3321 2381
rect 3318 2372 3321 2378
rect 3318 2272 3321 2358
rect 3326 2332 3329 2348
rect 3334 2342 3337 2368
rect 3342 2322 3345 2338
rect 3302 2152 3305 2188
rect 3302 1912 3305 2138
rect 3310 2042 3313 2148
rect 3326 2002 3329 2198
rect 3334 2132 3337 2138
rect 3278 1478 3286 1481
rect 3286 1442 3289 1478
rect 3294 1372 3297 1878
rect 3302 1752 3305 1768
rect 3302 1482 3305 1748
rect 3294 1342 3297 1368
rect 3302 1322 3305 1458
rect 3278 1272 3281 1278
rect 3230 1092 3233 1178
rect 3266 1148 3270 1151
rect 3214 1042 3217 1068
rect 3222 962 3225 1048
rect 3222 532 3225 958
rect 3238 742 3241 1128
rect 3182 262 3185 448
rect 3262 392 3265 1128
rect 3294 1102 3297 1258
rect 3310 1241 3313 1618
rect 3302 1238 3313 1241
rect 3302 1072 3305 1238
rect 3318 1212 3321 1928
rect 3326 1212 3329 1648
rect 3334 1562 3337 2128
rect 3314 1158 3318 1161
rect 3334 1152 3337 1558
rect 3342 1552 3345 2188
rect 3350 1882 3353 2498
rect 3358 2242 3361 2708
rect 3366 2512 3369 2618
rect 3366 2272 3369 2438
rect 3374 2322 3377 3198
rect 3382 3042 3385 3188
rect 3386 3018 3390 3021
rect 3400 3003 3402 3007
rect 3406 3003 3409 3007
rect 3414 3003 3416 3007
rect 3382 2262 3385 2948
rect 3390 2942 3393 2948
rect 3422 2932 3425 3358
rect 3430 3122 3433 3508
rect 3446 3342 3449 3408
rect 3462 3222 3465 3558
rect 3470 3512 3473 3758
rect 3478 3731 3481 4588
rect 3518 4542 3521 4568
rect 3530 4548 3534 4551
rect 3510 4328 3518 4331
rect 3490 4218 3494 4221
rect 3494 4101 3497 4158
rect 3490 4098 3497 4101
rect 3510 4062 3513 4328
rect 3526 4262 3529 4458
rect 3554 4258 3558 4261
rect 3526 4251 3529 4258
rect 3522 4248 3529 4251
rect 3510 4022 3513 4058
rect 3490 3948 3494 3951
rect 3478 3728 3489 3731
rect 3486 3672 3489 3728
rect 3486 3492 3489 3668
rect 3494 3552 3497 3868
rect 3502 3541 3505 3948
rect 3518 3892 3521 4108
rect 3494 3538 3505 3541
rect 3450 3158 3454 3161
rect 3430 3092 3433 3118
rect 3430 3032 3433 3068
rect 3400 2803 3402 2807
rect 3406 2803 3409 2807
rect 3414 2803 3416 2807
rect 3422 2622 3425 2918
rect 3400 2603 3402 2607
rect 3406 2603 3409 2607
rect 3414 2603 3416 2607
rect 3390 2522 3393 2598
rect 3410 2558 3414 2561
rect 3400 2403 3402 2407
rect 3406 2403 3409 2407
rect 3414 2403 3416 2407
rect 3394 2328 3398 2331
rect 3414 2322 3417 2338
rect 3406 2312 3409 2318
rect 3390 2252 3393 2308
rect 3374 2242 3377 2248
rect 3400 2203 3402 2207
rect 3406 2203 3409 2207
rect 3414 2203 3416 2207
rect 3362 2148 3366 2151
rect 3422 2092 3425 2618
rect 3430 2082 3433 2928
rect 3446 2382 3449 2928
rect 3462 2922 3465 3218
rect 3462 2722 3465 2818
rect 3454 2642 3457 2648
rect 3446 2351 3449 2358
rect 3442 2348 3449 2351
rect 3438 2272 3441 2288
rect 3410 2068 3414 2071
rect 3350 1552 3353 1878
rect 3342 1292 3345 1548
rect 3358 1432 3361 1818
rect 3366 1572 3369 2048
rect 3374 1982 3377 2068
rect 3374 1652 3377 1978
rect 3382 1812 3385 1898
rect 3382 1712 3385 1798
rect 3390 1652 3393 2018
rect 3400 2003 3402 2007
rect 3406 2003 3409 2007
rect 3414 2003 3416 2007
rect 3426 1968 3430 1971
rect 3414 1952 3417 1958
rect 3406 1832 3409 1948
rect 3400 1803 3402 1807
rect 3406 1803 3409 1807
rect 3414 1803 3416 1807
rect 3402 1658 3406 1661
rect 3390 1472 3393 1648
rect 3400 1603 3402 1607
rect 3406 1603 3409 1607
rect 3414 1603 3416 1607
rect 3422 1572 3425 1958
rect 3390 1372 3393 1448
rect 3400 1403 3402 1407
rect 3406 1403 3409 1407
rect 3414 1403 3416 1407
rect 3350 1362 3353 1368
rect 3358 1282 3361 1338
rect 3430 1302 3433 1548
rect 3438 1432 3441 2178
rect 3454 1972 3457 2228
rect 3462 2222 3465 2718
rect 3470 2652 3473 3108
rect 3486 2672 3489 3458
rect 3494 2752 3497 3538
rect 3502 3292 3505 3498
rect 3510 3422 3513 3668
rect 3518 3502 3521 3888
rect 3526 3852 3529 3988
rect 3574 3972 3577 4948
rect 3590 4912 3593 4948
rect 3582 4832 3585 4848
rect 3590 4482 3593 4908
rect 3686 4792 3689 5018
rect 3598 4242 3601 4258
rect 3526 3802 3529 3848
rect 3534 3712 3537 3738
rect 3542 3708 3550 3711
rect 3542 3702 3545 3708
rect 3518 3322 3521 3388
rect 3526 3262 3529 3548
rect 3534 2981 3537 3638
rect 3542 3392 3545 3698
rect 3558 3622 3561 3658
rect 3526 2978 3537 2981
rect 3494 2682 3497 2688
rect 3470 2472 3473 2518
rect 3470 2292 3473 2298
rect 3470 2262 3473 2268
rect 3334 1132 3337 1138
rect 3294 692 3297 728
rect 3302 491 3305 788
rect 3326 702 3329 1128
rect 3318 662 3321 698
rect 3298 488 3305 491
rect 3278 362 3281 418
rect 3342 382 3345 1258
rect 3358 1152 3361 1198
rect 3350 1062 3353 1148
rect 3358 1142 3361 1148
rect 3358 1122 3361 1128
rect 3366 1098 3374 1101
rect 3358 872 3361 878
rect 3366 872 3369 1098
rect 3390 492 3393 1208
rect 3400 1203 3402 1207
rect 3406 1203 3409 1207
rect 3414 1203 3416 1207
rect 3400 1003 3402 1007
rect 3406 1003 3409 1007
rect 3414 1003 3416 1007
rect 3438 952 3441 1008
rect 3446 962 3449 1658
rect 3454 1612 3457 1968
rect 3454 1592 3457 1608
rect 3462 1392 3465 2098
rect 3470 2012 3473 2208
rect 3478 1982 3481 2568
rect 3486 2412 3489 2528
rect 3486 2342 3489 2368
rect 3486 2322 3489 2328
rect 3486 2222 3489 2268
rect 3494 1862 3497 2608
rect 3502 2532 3505 2688
rect 3518 2452 3521 2468
rect 3506 2368 3510 2371
rect 3502 2272 3505 2348
rect 3518 2312 3521 2318
rect 3526 2282 3529 2978
rect 3542 2832 3545 2858
rect 3538 2658 3542 2661
rect 3534 2612 3537 2638
rect 3534 2282 3537 2608
rect 3550 2572 3553 3588
rect 3558 3242 3561 3618
rect 3566 3562 3569 3938
rect 3574 3502 3577 3898
rect 3566 3482 3569 3488
rect 3574 3472 3577 3488
rect 3574 3352 3577 3358
rect 3562 2968 3566 2971
rect 3558 2772 3561 2848
rect 3558 2592 3561 2598
rect 3522 2268 3526 2271
rect 3502 1732 3505 1948
rect 3470 962 3473 1538
rect 3494 1472 3497 1538
rect 3494 1042 3497 1218
rect 3502 1142 3505 1388
rect 3510 1282 3513 1848
rect 3518 1412 3521 2068
rect 3526 1402 3529 1988
rect 3526 1312 3529 1398
rect 3510 1032 3513 1138
rect 3418 868 3422 871
rect 3400 803 3402 807
rect 3406 803 3409 807
rect 3414 803 3416 807
rect 3422 668 3430 671
rect 3422 612 3425 668
rect 3438 652 3441 948
rect 3494 872 3497 968
rect 3498 758 3502 761
rect 3454 682 3457 688
rect 3400 603 3402 607
rect 3406 603 3409 607
rect 3414 603 3416 607
rect 3470 458 3478 461
rect 3470 452 3473 458
rect 3400 403 3402 407
rect 3406 403 3409 407
rect 3414 403 3416 407
rect 3194 348 3198 351
rect 2986 148 2990 151
rect 3082 148 3086 151
rect 3098 148 3102 151
rect 2888 103 2890 107
rect 2894 103 2897 107
rect 2902 103 2904 107
rect 2542 62 2545 78
rect 2822 62 2825 68
rect 2910 62 2913 98
rect 2934 62 2937 138
rect 3094 82 3097 148
rect 3382 92 3385 238
rect 3400 203 3402 207
rect 3406 203 3409 207
rect 3414 203 3416 207
rect 3390 62 3393 88
rect 3430 72 3433 78
rect 3438 72 3441 398
rect 3494 372 3497 678
rect 3486 272 3489 278
rect 3494 192 3497 368
rect 3494 152 3497 188
rect 3462 112 3465 138
rect 3470 92 3473 98
rect 3490 88 3494 91
rect 3502 82 3505 548
rect 3510 362 3513 1028
rect 3526 842 3529 1198
rect 3534 1072 3537 2068
rect 3542 1952 3545 2458
rect 3550 2292 3553 2538
rect 3558 2292 3561 2328
rect 3550 2252 3553 2258
rect 3566 2252 3569 2828
rect 3574 2742 3577 3348
rect 3582 2982 3585 3908
rect 3590 3772 3593 3848
rect 3590 3422 3593 3768
rect 3598 3752 3601 4238
rect 3606 3941 3609 4718
rect 3674 4708 3681 4711
rect 3634 4638 3641 4641
rect 3638 4432 3641 4638
rect 3638 4422 3641 4428
rect 3630 4062 3633 4178
rect 3618 3988 3625 3991
rect 3606 3938 3614 3941
rect 3622 3892 3625 3988
rect 3638 3982 3641 4168
rect 3598 3682 3601 3688
rect 3590 2702 3593 2718
rect 3574 2462 3577 2478
rect 3574 2272 3577 2408
rect 3582 2312 3585 2388
rect 3590 2282 3593 2528
rect 3598 2482 3601 3408
rect 3606 3332 3609 3338
rect 3606 3172 3609 3228
rect 3630 3112 3633 3858
rect 3638 3612 3641 3958
rect 3646 3952 3649 4088
rect 3654 3942 3657 4658
rect 3662 4372 3665 4518
rect 3662 4182 3665 4368
rect 3678 4261 3681 4708
rect 3686 4502 3689 4788
rect 3702 4752 3705 4948
rect 3726 4632 3729 4948
rect 3690 4498 3697 4501
rect 3694 4332 3697 4498
rect 3678 4258 3686 4261
rect 3690 4258 3697 4261
rect 3646 3472 3649 3888
rect 3654 3232 3657 3918
rect 3662 3672 3665 3688
rect 3626 3058 3630 3061
rect 3606 2672 3609 2678
rect 3606 2652 3609 2668
rect 3542 1938 3550 1941
rect 3542 1892 3545 1938
rect 3546 1868 3550 1871
rect 3550 1752 3553 1828
rect 3546 1748 3550 1751
rect 3542 1562 3545 1578
rect 3542 1161 3545 1378
rect 3550 1181 3553 1688
rect 3558 1332 3561 2068
rect 3558 1222 3561 1328
rect 3550 1178 3558 1181
rect 3542 1158 3550 1161
rect 3566 1161 3569 1738
rect 3574 1592 3577 1878
rect 3590 1832 3593 2128
rect 3598 2072 3601 2368
rect 3606 2172 3609 2638
rect 3614 2462 3617 2478
rect 3614 2362 3617 2388
rect 3614 2292 3617 2318
rect 3598 2052 3601 2058
rect 3606 1952 3609 2168
rect 3614 2072 3617 2078
rect 3622 1991 3625 2838
rect 3638 2782 3641 2928
rect 3646 2922 3649 3058
rect 3654 2882 3657 3228
rect 3662 3072 3665 3078
rect 3638 2692 3641 2778
rect 3670 2682 3673 4218
rect 3678 3572 3681 3968
rect 3686 3882 3689 3938
rect 3694 3902 3697 4258
rect 3702 4022 3705 4188
rect 3710 4052 3713 4398
rect 3718 4082 3721 4478
rect 3734 4472 3737 4548
rect 3726 4468 3734 4471
rect 3726 4452 3729 4468
rect 3726 4042 3729 4448
rect 3742 4272 3745 4728
rect 3830 4708 3838 4711
rect 3782 4352 3785 4618
rect 3830 4402 3833 4708
rect 3846 4551 3849 4928
rect 3920 4903 3922 4907
rect 3926 4903 3929 4907
rect 3934 4903 3936 4907
rect 3920 4703 3922 4707
rect 3926 4703 3929 4707
rect 3934 4703 3936 4707
rect 3886 4562 3889 4578
rect 3842 4548 3849 4551
rect 3870 4542 3873 4558
rect 3942 4552 3945 4558
rect 3838 4442 3841 4458
rect 3830 4328 3838 4331
rect 3830 4312 3833 4328
rect 3734 4268 3742 4271
rect 3722 3948 3726 3951
rect 3734 3932 3737 4268
rect 3678 3522 3681 3528
rect 3678 3152 3681 3328
rect 3686 3322 3689 3818
rect 3694 3592 3697 3878
rect 3702 3582 3705 3658
rect 3702 3562 3705 3568
rect 3694 3482 3697 3528
rect 3678 3072 3681 3088
rect 3694 3072 3697 3478
rect 3702 2982 3705 3558
rect 3718 3492 3721 3858
rect 3734 3682 3737 3728
rect 3726 3561 3729 3588
rect 3726 3558 3734 3561
rect 3726 3382 3729 3468
rect 3718 3342 3721 3368
rect 3710 3272 3713 3288
rect 3686 2882 3689 2978
rect 3654 2662 3657 2668
rect 3642 2658 3646 2661
rect 3646 2502 3649 2568
rect 3630 2482 3633 2498
rect 3646 2352 3649 2428
rect 3642 2348 3646 2351
rect 3634 2268 3638 2271
rect 3662 2262 3665 2658
rect 3686 2592 3689 2878
rect 3718 2742 3721 2768
rect 3726 2692 3729 3268
rect 3734 3152 3737 3308
rect 3742 3172 3745 4138
rect 3758 3772 3761 4198
rect 3774 3962 3777 4048
rect 3790 3972 3793 4188
rect 3766 3732 3769 3868
rect 3758 3562 3761 3698
rect 3750 3462 3753 3538
rect 3734 2822 3737 3148
rect 3742 3052 3745 3058
rect 3726 2672 3729 2688
rect 3734 2622 3737 2638
rect 3678 2332 3681 2348
rect 3678 2252 3681 2278
rect 3614 1988 3625 1991
rect 3574 1202 3577 1588
rect 3582 1332 3585 1798
rect 3582 1262 3585 1328
rect 3590 1322 3593 1618
rect 3598 1382 3601 1898
rect 3614 1882 3617 1988
rect 3614 1452 3617 1458
rect 3598 1368 3606 1371
rect 3566 1158 3574 1161
rect 3550 1051 3553 1158
rect 3598 1142 3601 1368
rect 3622 1151 3625 1978
rect 3670 1962 3673 2108
rect 3686 2082 3689 2588
rect 3694 2112 3697 2288
rect 3710 2182 3713 2588
rect 3686 2048 3694 2051
rect 3686 2032 3689 2048
rect 3670 1928 3678 1931
rect 3662 1872 3665 1898
rect 3634 1868 3638 1871
rect 3654 1782 3657 1858
rect 3670 1802 3673 1928
rect 3630 1182 3633 1538
rect 3630 1162 3633 1178
rect 3622 1148 3633 1151
rect 3546 1048 3561 1051
rect 3526 662 3529 838
rect 3542 652 3545 658
rect 3542 622 3545 648
rect 3550 472 3553 808
rect 3558 592 3561 1048
rect 3566 752 3569 788
rect 3542 462 3545 468
rect 3538 448 3542 451
rect 3526 412 3529 448
rect 3546 348 3550 351
rect 3566 272 3569 458
rect 3530 268 3534 271
rect 3534 62 3537 128
rect 3566 62 3569 268
rect 3574 252 3577 498
rect 3606 392 3609 1118
rect 3622 672 3625 1138
rect 3622 352 3625 668
rect 3630 632 3633 1148
rect 3638 1112 3641 1728
rect 3654 1702 3657 1738
rect 3646 1668 3654 1671
rect 3646 1652 3649 1668
rect 3654 1472 3657 1658
rect 3650 1458 3654 1461
rect 3638 1051 3641 1108
rect 3638 1048 3646 1051
rect 3654 862 3657 868
rect 3638 702 3641 808
rect 3638 532 3641 548
rect 3662 452 3665 1558
rect 3674 1358 3678 1361
rect 3686 1052 3689 1978
rect 3710 1942 3713 2178
rect 3718 2172 3721 2598
rect 3730 2468 3734 2471
rect 3734 2422 3737 2448
rect 3734 2362 3737 2398
rect 3726 2182 3729 2268
rect 3734 2142 3737 2148
rect 3722 2058 3726 2061
rect 3710 1842 3713 1848
rect 3726 1792 3729 2048
rect 3742 2042 3745 2718
rect 3750 2642 3753 3458
rect 3758 2722 3761 2758
rect 3766 2692 3769 3728
rect 3774 3531 3777 3958
rect 3790 3952 3793 3968
rect 3798 3852 3801 3868
rect 3810 3848 3814 3851
rect 3774 3528 3785 3531
rect 3750 1922 3753 2598
rect 3766 2372 3769 2688
rect 3774 2572 3777 3478
rect 3782 2772 3785 3528
rect 3806 3522 3809 3528
rect 3822 3492 3825 4188
rect 3830 4182 3833 4308
rect 3854 4142 3857 4348
rect 3790 3182 3793 3328
rect 3814 3242 3817 3258
rect 3798 2782 3801 2968
rect 3782 2662 3785 2768
rect 3802 2728 3809 2731
rect 3806 2712 3809 2728
rect 3798 2672 3801 2678
rect 3790 2662 3793 2668
rect 3774 2542 3777 2558
rect 3782 2512 3785 2608
rect 3794 2548 3798 2551
rect 3758 2102 3761 2328
rect 3758 2081 3761 2098
rect 3774 2082 3777 2258
rect 3758 2078 3766 2081
rect 3698 1538 3702 1541
rect 3678 871 3681 908
rect 3674 868 3681 871
rect 3686 452 3689 598
rect 3694 552 3697 1158
rect 3702 582 3705 1358
rect 3726 1172 3729 1238
rect 3726 942 3729 1118
rect 3734 972 3737 1468
rect 3742 1392 3745 1438
rect 3750 1382 3753 1918
rect 3766 1822 3769 2058
rect 3778 1878 3782 1881
rect 3790 1762 3793 2308
rect 3766 1312 3769 1638
rect 3742 1232 3745 1238
rect 3710 751 3713 938
rect 3730 858 3734 861
rect 3718 842 3721 858
rect 3710 748 3718 751
rect 3710 472 3713 688
rect 3742 542 3745 1098
rect 3758 1071 3761 1258
rect 3774 1162 3777 1588
rect 3790 1372 3793 1758
rect 3798 1441 3801 2368
rect 3806 2102 3809 2708
rect 3814 2612 3817 3238
rect 3822 2552 3825 3308
rect 3830 2852 3833 3558
rect 3830 2632 3833 2658
rect 3814 2262 3817 2508
rect 3822 2392 3825 2548
rect 3838 2472 3841 3238
rect 3846 3152 3849 3158
rect 3854 2842 3857 4028
rect 3862 3252 3865 3958
rect 3862 2762 3865 3068
rect 3870 2902 3873 4538
rect 3920 4503 3922 4507
rect 3926 4503 3929 4507
rect 3934 4503 3936 4507
rect 3942 4491 3945 4508
rect 3938 4488 3945 4491
rect 3934 4352 3937 4368
rect 3882 4348 3889 4351
rect 3886 4342 3889 4348
rect 3920 4303 3922 4307
rect 3926 4303 3929 4307
rect 3934 4303 3936 4307
rect 3902 4122 3905 4158
rect 3910 4112 3913 4118
rect 3920 4103 3922 4107
rect 3926 4103 3929 4107
rect 3934 4103 3936 4107
rect 3890 4078 3894 4081
rect 3894 3982 3897 4038
rect 3910 3952 3913 4078
rect 3920 3903 3922 3907
rect 3926 3903 3929 3907
rect 3934 3903 3936 3907
rect 3882 3848 3886 3851
rect 3898 3708 3902 3711
rect 3920 3703 3922 3707
rect 3926 3703 3929 3707
rect 3934 3703 3936 3707
rect 3942 3692 3945 4478
rect 3894 3672 3897 3678
rect 3920 3503 3922 3507
rect 3926 3503 3929 3507
rect 3934 3503 3936 3507
rect 3894 2992 3897 3148
rect 3902 3072 3905 3348
rect 3920 3303 3922 3307
rect 3926 3303 3929 3307
rect 3934 3303 3936 3307
rect 3942 3192 3945 3528
rect 3920 3103 3922 3107
rect 3926 3103 3929 3107
rect 3934 3103 3936 3107
rect 3910 3062 3913 3098
rect 3942 3072 3945 3098
rect 3838 2442 3841 2468
rect 3846 2322 3849 2758
rect 3826 2268 3830 2271
rect 3854 2241 3857 2698
rect 3862 2682 3865 2758
rect 3854 2238 3862 2241
rect 3806 2052 3809 2058
rect 3810 1548 3814 1551
rect 3798 1438 3809 1441
rect 3782 1292 3785 1298
rect 3798 1292 3801 1428
rect 3782 1152 3785 1178
rect 3770 1148 3774 1151
rect 3754 1068 3761 1071
rect 3750 972 3753 978
rect 3766 902 3769 1058
rect 3774 712 3777 1078
rect 3774 552 3777 708
rect 3662 372 3665 448
rect 3574 92 3577 118
rect 3606 62 3609 148
rect 3646 142 3649 218
rect 3654 212 3657 338
rect 3662 282 3665 368
rect 3702 362 3705 468
rect 3638 102 3641 128
rect 3710 92 3713 278
rect 3734 72 3737 478
rect 3774 412 3777 548
rect 3782 452 3785 1078
rect 3790 972 3793 1258
rect 3798 952 3801 1288
rect 3806 1162 3809 1438
rect 3814 1302 3817 1308
rect 3798 562 3801 868
rect 3806 732 3809 868
rect 3814 752 3817 1168
rect 3822 902 3825 2168
rect 3838 2152 3841 2188
rect 3830 1532 3833 2138
rect 3846 1592 3849 2098
rect 3854 1732 3857 2038
rect 3870 1931 3873 2898
rect 3886 2732 3889 2988
rect 3878 2728 3886 2731
rect 3878 2472 3881 2728
rect 3886 2462 3889 2688
rect 3894 2412 3897 2928
rect 3902 2582 3905 2908
rect 3920 2903 3922 2907
rect 3926 2903 3929 2907
rect 3934 2903 3936 2907
rect 3920 2703 3922 2707
rect 3926 2703 3929 2707
rect 3934 2703 3936 2707
rect 3910 2512 3913 2548
rect 3920 2503 3922 2507
rect 3926 2503 3929 2507
rect 3934 2503 3936 2507
rect 3950 2492 3953 5048
rect 4078 4792 4081 5058
rect 4518 5018 4526 5021
rect 4094 4892 4097 4948
rect 4126 4832 4129 4938
rect 4134 4922 4137 5018
rect 4424 5003 4426 5007
rect 4430 5003 4433 5007
rect 4438 5003 4440 5007
rect 4190 4942 4193 4978
rect 4134 4852 4137 4858
rect 4030 4702 4033 4738
rect 3962 4548 3966 4551
rect 3962 4538 3966 4541
rect 3974 4032 3977 4448
rect 3958 3132 3961 3498
rect 3902 2412 3905 2448
rect 3958 2372 3961 3018
rect 3966 2862 3969 3508
rect 3974 3222 3977 4028
rect 3998 3882 4001 4528
rect 4030 4462 4033 4698
rect 4038 4462 4041 4788
rect 4006 4212 4009 4438
rect 3994 3758 3998 3761
rect 4006 3742 4009 3758
rect 3998 3722 4001 3728
rect 3982 3652 3985 3718
rect 3990 3592 3993 3608
rect 3998 3482 4001 3708
rect 4006 3572 4009 3658
rect 4014 3572 4017 3708
rect 3982 3302 3985 3308
rect 3966 2442 3969 2808
rect 3886 2202 3889 2328
rect 3894 2192 3897 2358
rect 3910 2272 3913 2308
rect 3920 2303 3922 2307
rect 3926 2303 3929 2307
rect 3934 2303 3936 2307
rect 3974 2301 3977 2708
rect 3982 2532 3985 2938
rect 3982 2352 3985 2378
rect 3990 2312 3993 2958
rect 3998 2802 4001 3478
rect 4006 2502 4009 3448
rect 4022 3442 4025 3948
rect 4030 3902 4033 4458
rect 4038 4128 4046 4131
rect 4038 4122 4041 4128
rect 4054 4082 4057 4588
rect 4062 4332 4065 4338
rect 4062 4302 4065 4328
rect 4070 4252 4073 4688
rect 4078 4552 4081 4558
rect 4094 4502 4097 4738
rect 4102 4538 4110 4541
rect 4102 4532 4105 4538
rect 4098 4468 4105 4471
rect 4102 4442 4105 4468
rect 4078 4062 4081 4298
rect 4086 4062 4089 4358
rect 4102 4288 4110 4291
rect 4094 4152 4097 4208
rect 4070 4022 4073 4048
rect 4030 3532 4033 3608
rect 4030 3482 4033 3528
rect 3974 2298 3982 2301
rect 3998 2282 4001 2308
rect 3866 1928 3873 1931
rect 3862 1832 3865 1918
rect 3830 1302 3833 1318
rect 3830 1032 3833 1048
rect 3822 892 3825 898
rect 3822 852 3825 888
rect 3814 722 3817 748
rect 3814 672 3817 718
rect 3806 362 3809 588
rect 3830 522 3833 1028
rect 3838 682 3841 1568
rect 3846 1522 3849 1548
rect 3854 1452 3857 1488
rect 3870 1482 3873 1828
rect 3854 1322 3857 1418
rect 3854 762 3857 1318
rect 3870 1272 3873 1278
rect 3878 1072 3881 2138
rect 3894 2092 3897 2148
rect 3942 2112 3945 2148
rect 3920 2103 3922 2107
rect 3926 2103 3929 2107
rect 3934 2103 3936 2107
rect 3886 2042 3889 2048
rect 3894 1922 3897 2058
rect 3920 1903 3922 1907
rect 3926 1903 3929 1907
rect 3934 1903 3936 1907
rect 3942 1892 3945 1898
rect 3902 1582 3905 1698
rect 3910 1692 3913 1858
rect 3920 1703 3922 1707
rect 3926 1703 3929 1707
rect 3934 1703 3936 1707
rect 3910 1571 3913 1688
rect 3906 1568 3913 1571
rect 3902 1552 3905 1558
rect 3890 1548 3894 1551
rect 3920 1503 3922 1507
rect 3926 1503 3929 1507
rect 3934 1503 3936 1507
rect 3942 1402 3945 1738
rect 3886 1262 3889 1278
rect 3866 858 3870 861
rect 3886 812 3889 1018
rect 3902 892 3905 1338
rect 3950 1332 3953 1808
rect 3920 1303 3922 1307
rect 3926 1303 3929 1307
rect 3934 1303 3936 1307
rect 3910 1292 3913 1298
rect 3934 1122 3937 1138
rect 3920 1103 3922 1107
rect 3926 1103 3929 1107
rect 3934 1103 3936 1107
rect 3910 912 3913 918
rect 3920 903 3922 907
rect 3926 903 3929 907
rect 3934 903 3936 907
rect 3838 562 3841 678
rect 3910 572 3913 738
rect 3920 703 3922 707
rect 3926 703 3929 707
rect 3934 703 3936 707
rect 3942 632 3945 1248
rect 3950 852 3953 1328
rect 3958 1132 3961 1868
rect 3966 1782 3969 2198
rect 3974 1872 3977 1898
rect 3978 1858 3982 1861
rect 3966 1462 3969 1778
rect 3978 1748 3982 1751
rect 3958 1092 3961 1128
rect 3958 912 3961 988
rect 3966 862 3969 1378
rect 3974 1232 3977 1448
rect 3990 1382 3993 1898
rect 3998 1672 4001 1878
rect 3942 582 3945 628
rect 3974 582 3977 948
rect 3982 752 3985 1318
rect 3990 1282 3993 1298
rect 3990 862 3993 1218
rect 3998 1062 4001 1558
rect 4006 1162 4009 2368
rect 4014 2062 4017 3438
rect 4026 3268 4030 3271
rect 4026 3088 4030 3091
rect 4038 3062 4041 3968
rect 4070 3882 4073 3928
rect 4054 3492 4057 3758
rect 4062 3542 4065 3558
rect 4070 3542 4073 3548
rect 4022 3002 4025 3058
rect 4022 2632 4025 2998
rect 4046 2952 4049 3468
rect 4062 3262 4065 3298
rect 4062 3152 4065 3258
rect 4046 2862 4049 2908
rect 4038 2858 4046 2861
rect 4030 2522 4033 2778
rect 4038 2592 4041 2858
rect 4054 2592 4057 2628
rect 4054 2552 4057 2588
rect 4038 2472 4041 2518
rect 4046 2452 4049 2478
rect 4014 1852 4017 1878
rect 4022 1852 4025 2318
rect 4022 1602 4025 1688
rect 4014 1352 4017 1378
rect 4006 972 4009 1158
rect 3826 458 3830 461
rect 3838 352 3841 358
rect 3746 258 3750 261
rect 3894 212 3897 528
rect 3902 472 3905 558
rect 3910 472 3913 568
rect 3920 503 3922 507
rect 3926 503 3929 507
rect 3934 503 3936 507
rect 3982 472 3985 668
rect 3998 662 4001 858
rect 4014 752 4017 1348
rect 4030 1272 4033 2258
rect 4038 2242 4041 2258
rect 4038 2072 4041 2128
rect 4046 2002 4049 2448
rect 4054 2032 4057 2238
rect 4062 2082 4065 3108
rect 4070 2422 4073 3338
rect 4078 2962 4081 3878
rect 4086 3622 4089 3948
rect 4094 3662 4097 4148
rect 4102 4112 4105 4288
rect 4118 4262 4121 4568
rect 4126 4342 4129 4828
rect 4134 4792 4137 4828
rect 4150 4752 4153 4798
rect 4134 4372 4137 4728
rect 4142 4562 4145 4568
rect 4142 4532 4145 4538
rect 4150 4452 4153 4748
rect 4170 4558 4174 4561
rect 4182 4442 4185 4918
rect 4134 4272 4137 4368
rect 4090 3618 4097 3621
rect 4094 3432 4097 3618
rect 4102 3362 4105 3918
rect 4102 3322 4105 3348
rect 4086 3272 4089 3278
rect 4110 3212 4113 3788
rect 4118 3192 4121 3928
rect 4126 3912 4129 3958
rect 4142 3911 4145 4078
rect 4138 3908 4145 3911
rect 4142 3472 4145 3908
rect 4134 3172 4137 3218
rect 4086 3072 4089 3108
rect 4082 2748 4086 2751
rect 4078 2692 4081 2708
rect 4070 2362 4073 2408
rect 4078 2192 4081 2498
rect 4086 2222 4089 2738
rect 4094 2462 4097 2988
rect 4114 2838 4118 2841
rect 4126 2832 4129 3148
rect 4134 2822 4137 3168
rect 4142 3022 4145 3428
rect 4150 3162 4153 4368
rect 4158 4262 4161 4268
rect 4158 4192 4161 4258
rect 4166 4142 4169 4418
rect 4190 4352 4193 4938
rect 4218 4848 4225 4851
rect 4222 4842 4225 4848
rect 4206 4572 4209 4718
rect 4214 4562 4217 4818
rect 4202 4528 4206 4531
rect 4182 4292 4185 4338
rect 4158 3552 4161 4018
rect 4158 3262 4161 3518
rect 4150 2952 4153 3058
rect 4078 2011 4081 2188
rect 4094 2162 4097 2458
rect 4102 2362 4105 2748
rect 4110 2612 4113 2748
rect 4110 2472 4113 2498
rect 4094 2062 4097 2098
rect 4078 2008 4089 2011
rect 4078 1942 4081 1998
rect 4066 1938 4073 1941
rect 4070 1922 4073 1938
rect 4050 1868 4054 1871
rect 4070 1772 4073 1918
rect 4086 1772 4089 2008
rect 4054 1482 4057 1498
rect 4054 1342 4057 1428
rect 4022 1152 4025 1158
rect 4030 762 4033 778
rect 3978 468 3982 471
rect 3920 303 3922 307
rect 3926 303 3929 307
rect 3934 303 3936 307
rect 3998 272 4001 658
rect 4014 552 4017 668
rect 4026 528 4030 531
rect 4030 352 4033 418
rect 4038 402 4041 658
rect 4046 482 4049 1068
rect 4054 692 4057 868
rect 4062 682 4065 1618
rect 4070 772 4073 1688
rect 4094 1652 4097 1928
rect 4102 1572 4105 2338
rect 4110 1992 4113 2038
rect 4110 1542 4113 1628
rect 4110 1522 4113 1538
rect 4078 952 4081 1258
rect 4086 1062 4089 1098
rect 4078 862 4081 948
rect 4086 898 4094 901
rect 4086 732 4089 898
rect 4102 892 4105 1508
rect 4110 1252 4113 1258
rect 4082 648 4086 651
rect 4094 512 4097 848
rect 4118 662 4121 2548
rect 4126 982 4129 2698
rect 4134 2652 4137 2818
rect 4142 2702 4145 2928
rect 4134 2552 4137 2558
rect 4142 2482 4145 2698
rect 4134 1152 4137 2268
rect 4142 2112 4145 2478
rect 4158 2392 4161 3258
rect 4166 3002 4169 3668
rect 4174 3092 4177 3618
rect 4182 3422 4185 4208
rect 4190 4132 4193 4148
rect 4206 3872 4209 4348
rect 4214 4272 4217 4358
rect 4214 4132 4217 4248
rect 4230 4072 4233 4678
rect 4238 4122 4241 4538
rect 4246 4452 4249 4458
rect 4254 4272 4257 4688
rect 4238 4052 4241 4068
rect 4238 4038 4246 4041
rect 4190 3672 4193 3698
rect 4198 3642 4201 3658
rect 4190 3532 4193 3628
rect 4206 3542 4209 3638
rect 4190 3432 4193 3528
rect 4190 3392 4193 3418
rect 4198 3232 4201 3308
rect 4174 3062 4177 3068
rect 4174 2892 4177 2938
rect 4174 2142 4177 2748
rect 4174 2072 4177 2078
rect 4146 2068 4150 2071
rect 4146 2038 4150 2041
rect 4142 1612 4145 1758
rect 4150 1662 4153 1908
rect 4158 1562 4161 1868
rect 4170 1818 4174 1821
rect 4182 1802 4185 3188
rect 4198 3032 4201 3228
rect 4190 2962 4193 3008
rect 4190 2862 4193 2938
rect 4190 2682 4193 2858
rect 4206 2832 4209 3518
rect 4214 3332 4217 3688
rect 4214 3252 4217 3258
rect 4222 2782 4225 3628
rect 4230 3071 4233 3818
rect 4238 3682 4241 4038
rect 4230 3068 4241 3071
rect 4238 2772 4241 3068
rect 4246 2852 4249 3858
rect 4254 3652 4257 4118
rect 4262 4102 4265 4328
rect 4270 3952 4273 4848
rect 4278 4552 4281 4558
rect 4278 4122 4281 4548
rect 4286 4072 4289 4908
rect 4398 4572 4401 4798
rect 4406 4552 4409 4868
rect 4424 4803 4426 4807
rect 4430 4803 4433 4807
rect 4438 4803 4440 4807
rect 4414 4622 4417 4698
rect 4414 4562 4417 4618
rect 4424 4603 4426 4607
rect 4430 4603 4433 4607
rect 4438 4603 4440 4607
rect 4294 4062 4297 4368
rect 4262 3948 4270 3951
rect 4262 3092 4265 3948
rect 4274 3658 4278 3661
rect 4254 3052 4257 3058
rect 4214 2662 4217 2668
rect 4206 2658 4214 2661
rect 4190 2482 4193 2618
rect 4190 2262 4193 2268
rect 4190 2062 4193 2138
rect 4190 1982 4193 2058
rect 4190 1902 4193 1908
rect 4178 1758 4182 1761
rect 4142 1538 4150 1541
rect 4142 1492 4145 1538
rect 4158 1392 4161 1558
rect 4166 1472 4169 1718
rect 4174 1682 4177 1718
rect 4174 1252 4177 1678
rect 4190 1652 4193 1748
rect 4198 1662 4201 2468
rect 4198 1562 4201 1658
rect 4194 1538 4198 1541
rect 4186 1468 4190 1471
rect 4166 1152 4169 1188
rect 4174 1071 4177 1168
rect 4174 1068 4182 1071
rect 4178 1048 4182 1051
rect 4134 1042 4137 1048
rect 4142 1038 4150 1041
rect 4142 1032 4145 1038
rect 4174 812 4177 838
rect 4166 802 4169 808
rect 4150 772 4153 798
rect 4114 458 4118 461
rect 3998 262 4001 268
rect 3894 92 3897 208
rect 4102 162 4105 408
rect 4126 362 4129 668
rect 4134 492 4137 588
rect 4150 552 4153 758
rect 4166 502 4169 798
rect 3978 138 3982 141
rect 4066 138 4070 141
rect 3920 103 3922 107
rect 3926 103 3929 107
rect 3934 103 3936 107
rect 3942 92 3945 108
rect 4118 91 4121 158
rect 4118 88 4126 91
rect 3914 68 3918 71
rect 4150 62 4153 488
rect 4166 442 4169 448
rect 4174 342 4177 698
rect 4190 682 4193 1468
rect 4206 1132 4209 2658
rect 4214 1992 4217 2468
rect 4230 2412 4233 2498
rect 4238 2372 4241 2488
rect 4246 2432 4249 2828
rect 4262 2682 4265 3058
rect 4270 2472 4273 3238
rect 4278 2752 4281 3558
rect 4286 3532 4289 4048
rect 4302 3982 4305 4338
rect 4302 2942 4305 3808
rect 4310 3612 4313 3628
rect 4318 3592 4321 4168
rect 4342 4162 4345 4358
rect 4350 4232 4353 4398
rect 4310 3502 4313 3548
rect 4310 3462 4313 3498
rect 4310 3082 4313 3278
rect 4318 3252 4321 3528
rect 4286 2862 4289 2878
rect 4278 2532 4281 2538
rect 4254 2452 4257 2458
rect 4286 2452 4289 2578
rect 4294 2472 4297 2888
rect 4302 2702 4305 2708
rect 4302 2642 4305 2648
rect 4234 2278 4241 2281
rect 4238 2262 4241 2278
rect 4222 1872 4225 2068
rect 4214 1562 4217 1828
rect 4222 1762 4225 1788
rect 4230 1571 4233 1998
rect 4238 1722 4241 2048
rect 4246 1962 4249 2098
rect 4246 1832 4249 1858
rect 4238 1642 4241 1678
rect 4242 1638 4246 1641
rect 4230 1568 4238 1571
rect 4222 1362 4225 1508
rect 4218 1348 4222 1351
rect 4206 1092 4209 1128
rect 4230 1062 4233 1558
rect 4242 1538 4246 1541
rect 4246 1022 4249 1478
rect 4206 962 4209 988
rect 4198 471 4201 908
rect 4238 862 4241 988
rect 4254 882 4257 2128
rect 4262 1511 4265 2208
rect 4270 1892 4273 2438
rect 4270 1742 4273 1758
rect 4278 1592 4281 2208
rect 4286 2152 4289 2318
rect 4294 1832 4297 2428
rect 4302 2322 4305 2528
rect 4310 2522 4313 2948
rect 4318 2932 4321 3248
rect 4326 3192 4329 4138
rect 4358 4091 4361 4188
rect 4358 4088 4366 4091
rect 4358 4012 4361 4088
rect 4350 3961 4353 3988
rect 4346 3958 4353 3961
rect 4342 3861 4345 3878
rect 4338 3858 4345 3861
rect 4334 3562 4337 3758
rect 4350 3732 4353 3958
rect 4358 3692 4361 3998
rect 4390 3932 4393 4478
rect 4424 4403 4426 4407
rect 4430 4403 4433 4407
rect 4438 4403 4440 4407
rect 4402 4288 4406 4291
rect 4398 4202 4401 4238
rect 4374 3822 4377 3848
rect 4366 3662 4369 3788
rect 4374 3642 4377 3748
rect 4334 3262 4337 3268
rect 4334 2972 4337 3248
rect 4366 3212 4369 3548
rect 4382 3532 4385 3768
rect 4398 3741 4401 4128
rect 4390 3738 4401 3741
rect 4346 3168 4353 3171
rect 4350 2952 4353 3168
rect 4374 3082 4377 3338
rect 4318 2652 4321 2928
rect 4326 2532 4329 2858
rect 4346 2768 4350 2771
rect 4310 2352 4313 2518
rect 4302 2152 4305 2318
rect 4302 1552 4305 2098
rect 4318 2092 4321 2328
rect 4326 2152 4329 2478
rect 4334 2292 4337 2718
rect 4350 2672 4353 2758
rect 4358 2672 4361 3078
rect 4366 2952 4369 2958
rect 4342 2532 4345 2648
rect 4358 2632 4361 2668
rect 4350 2422 4353 2468
rect 4310 1892 4313 2028
rect 4318 1842 4321 1958
rect 4318 1832 4321 1838
rect 4262 1508 4270 1511
rect 4310 1472 4313 1718
rect 4318 1552 4321 1568
rect 4270 1322 4273 1458
rect 4278 1322 4281 1328
rect 4282 1278 4286 1281
rect 4262 1262 4265 1278
rect 4294 1142 4297 1148
rect 4262 1022 4265 1068
rect 4266 848 4270 851
rect 4206 652 4209 658
rect 4198 468 4206 471
rect 4198 262 4201 348
rect 4214 272 4217 548
rect 4222 342 4225 728
rect 4302 662 4305 1198
rect 4310 1032 4313 1338
rect 4318 922 4321 1538
rect 4326 1312 4329 2088
rect 4342 2072 4345 2108
rect 4342 2062 4345 2068
rect 4350 2032 4353 2348
rect 4358 2232 4361 2618
rect 4350 1782 4353 1938
rect 4334 1562 4337 1568
rect 4330 1268 4334 1271
rect 4326 1252 4329 1258
rect 4342 1252 4345 1718
rect 4350 1492 4353 1768
rect 4358 1542 4361 2228
rect 4366 2092 4369 2658
rect 4374 2622 4377 3058
rect 4382 2592 4385 3318
rect 4390 2972 4393 3738
rect 4398 3662 4401 3678
rect 4398 3032 4401 3548
rect 4406 3012 4409 4278
rect 4414 4072 4417 4288
rect 4424 4203 4426 4207
rect 4430 4203 4433 4207
rect 4438 4203 4440 4207
rect 4424 4003 4426 4007
rect 4430 4003 4433 4007
rect 4438 4003 4440 4007
rect 4424 3803 4426 3807
rect 4430 3803 4433 3807
rect 4438 3803 4440 3807
rect 4414 3612 4417 3768
rect 4446 3622 4449 4728
rect 4454 3882 4457 4358
rect 4478 4282 4481 4628
rect 4502 4552 4505 4788
rect 4462 3892 4465 4038
rect 4462 3862 4465 3888
rect 4414 3462 4417 3608
rect 4424 3603 4426 3607
rect 4430 3603 4433 3607
rect 4438 3603 4440 3607
rect 4424 3403 4426 3407
rect 4430 3403 4433 3407
rect 4438 3403 4440 3407
rect 4424 3203 4426 3207
rect 4430 3203 4433 3207
rect 4438 3203 4440 3207
rect 4414 3152 4417 3158
rect 4446 3152 4449 3588
rect 4470 3542 4473 4148
rect 4470 3412 4473 3468
rect 4478 3372 4481 4208
rect 4486 4142 4489 4338
rect 4494 4022 4497 4348
rect 4486 3452 4489 4018
rect 4494 3962 4497 3978
rect 4502 3912 4505 4408
rect 4510 3961 4513 4098
rect 4518 4022 4521 5018
rect 4526 4372 4529 4948
rect 4526 4202 4529 4368
rect 4510 3958 4521 3961
rect 4494 3532 4497 3538
rect 4502 3532 4505 3548
rect 4510 3422 4513 3948
rect 4518 3462 4521 3958
rect 4534 3912 4537 4838
rect 4550 4798 4558 4801
rect 4550 4662 4553 4798
rect 4570 4748 4574 4751
rect 4542 3782 4545 4298
rect 4562 4258 4566 4261
rect 4550 3762 4553 4248
rect 4530 3548 4534 3551
rect 4414 3122 4417 3128
rect 4424 3003 4426 3007
rect 4430 3003 4433 3007
rect 4438 3003 4440 3007
rect 4398 2958 4406 2961
rect 4390 2752 4393 2948
rect 4398 2942 4401 2958
rect 4390 2672 4393 2678
rect 4398 2601 4401 2878
rect 4390 2598 4401 2601
rect 4374 2152 4377 2518
rect 4390 2472 4393 2598
rect 4382 2112 4385 2138
rect 4378 2038 4382 2041
rect 4366 1962 4369 1998
rect 4366 1532 4369 1958
rect 4374 1542 4377 1928
rect 4390 1922 4393 2188
rect 4398 2012 4401 2588
rect 4406 2402 4409 2708
rect 4414 2652 4417 2978
rect 4422 2952 4425 2958
rect 4424 2803 4426 2807
rect 4430 2803 4433 2807
rect 4438 2803 4440 2807
rect 4424 2603 4426 2607
rect 4430 2603 4433 2607
rect 4438 2603 4440 2607
rect 4426 2538 4430 2541
rect 4414 2472 4417 2478
rect 4430 2462 4433 2468
rect 4406 2212 4409 2398
rect 4398 1582 4401 2008
rect 4406 1822 4409 2138
rect 4414 2112 4417 2448
rect 4424 2403 4426 2407
rect 4430 2403 4433 2407
rect 4438 2403 4440 2407
rect 4438 2232 4441 2288
rect 4446 2212 4449 2968
rect 4454 2732 4457 3268
rect 4462 3102 4465 3358
rect 4486 3292 4489 3358
rect 4502 3341 4505 3348
rect 4498 3338 4505 3341
rect 4506 3268 4510 3271
rect 4494 3262 4497 3268
rect 4482 3258 4486 3261
rect 4518 3202 4521 3358
rect 4534 3261 4537 3318
rect 4530 3258 4537 3261
rect 4518 3122 4521 3168
rect 4526 3152 4529 3178
rect 4534 3152 4537 3248
rect 4462 2661 4465 2718
rect 4470 2712 4473 3098
rect 4458 2658 4465 2661
rect 4470 2612 4473 2688
rect 4424 2203 4426 2207
rect 4430 2203 4433 2207
rect 4438 2203 4440 2207
rect 4414 2082 4417 2108
rect 4424 2003 4426 2007
rect 4430 2003 4433 2007
rect 4438 2003 4440 2007
rect 4414 1812 4417 1968
rect 4424 1803 4426 1807
rect 4430 1803 4433 1807
rect 4438 1803 4440 1807
rect 4406 1612 4409 1618
rect 4358 1502 4361 1508
rect 4374 1432 4377 1538
rect 4382 1492 4385 1578
rect 4398 1542 4401 1568
rect 4382 1352 4385 1398
rect 4390 1312 4393 1538
rect 4406 1512 4409 1548
rect 4398 1452 4401 1498
rect 4406 1342 4409 1478
rect 4414 1362 4417 1798
rect 4424 1603 4426 1607
rect 4430 1603 4433 1607
rect 4438 1603 4440 1607
rect 4424 1403 4426 1407
rect 4430 1403 4433 1407
rect 4438 1403 4440 1407
rect 4446 1362 4449 2148
rect 4454 2132 4457 2548
rect 4462 2432 4465 2528
rect 4462 2272 4465 2428
rect 4454 2002 4457 2098
rect 4454 1662 4457 1758
rect 4454 1412 4457 1488
rect 4390 1252 4393 1308
rect 4326 1192 4329 1248
rect 4350 1128 4358 1131
rect 4214 152 4217 268
rect 4310 142 4313 668
rect 4326 662 4329 718
rect 4342 542 4345 908
rect 4350 792 4353 1128
rect 4362 1118 4366 1121
rect 4374 1062 4377 1068
rect 4390 872 4393 1248
rect 4398 1052 4401 1248
rect 4390 862 4393 868
rect 2730 58 2734 61
rect 2962 58 2966 61
rect 4246 61 4249 108
rect 4374 92 4377 768
rect 4398 702 4401 938
rect 4406 512 4409 1328
rect 4446 1262 4449 1298
rect 4424 1203 4426 1207
rect 4430 1203 4433 1207
rect 4438 1203 4440 1207
rect 4424 1003 4426 1007
rect 4430 1003 4433 1007
rect 4438 1003 4440 1007
rect 4414 962 4417 998
rect 4446 992 4449 1258
rect 4454 1122 4457 1198
rect 4424 803 4426 807
rect 4430 803 4433 807
rect 4438 803 4440 807
rect 4446 732 4449 828
rect 4454 722 4457 1028
rect 4462 822 4465 2258
rect 4470 1562 4473 2548
rect 4478 2262 4481 3008
rect 4490 2958 4494 2961
rect 4486 2582 4489 2858
rect 4470 1462 4473 1468
rect 4470 1362 4473 1368
rect 4478 951 4481 2078
rect 4486 1032 4489 2558
rect 4494 2552 4497 2938
rect 4510 2912 4513 2938
rect 4526 2932 4529 2938
rect 4542 2882 4545 3758
rect 4566 3532 4569 3578
rect 4526 2852 4529 2868
rect 4538 2858 4542 2861
rect 4502 2662 4505 2678
rect 4534 2662 4537 2858
rect 4550 2851 4553 3378
rect 4558 3302 4561 3508
rect 4574 3342 4577 4598
rect 4582 3572 4585 4798
rect 4606 4582 4609 4858
rect 4590 3902 4593 4398
rect 4606 4132 4609 4438
rect 4614 3962 4617 4968
rect 4678 4732 4681 4898
rect 4638 4591 4641 4698
rect 4634 4588 4641 4591
rect 4626 4458 4630 4461
rect 4646 4362 4649 4598
rect 4654 4592 4657 4678
rect 4666 4658 4670 4661
rect 4678 4562 4681 4728
rect 4622 4332 4625 4338
rect 4642 4288 4646 4291
rect 4610 3948 4617 3951
rect 4614 3942 4617 3948
rect 4558 3222 4561 3238
rect 4566 3162 4569 3168
rect 4542 2848 4553 2851
rect 4494 1662 4497 2098
rect 4502 2052 4505 2598
rect 4510 2052 4513 2078
rect 4518 2042 4521 2468
rect 4502 1742 4505 1778
rect 4526 1672 4529 2608
rect 4534 2262 4537 2648
rect 4542 2452 4545 2848
rect 4534 2092 4537 2258
rect 4534 1842 4537 1878
rect 4494 1542 4497 1658
rect 4498 1508 4502 1511
rect 4526 1482 4529 1668
rect 4474 948 4481 951
rect 4486 942 4489 948
rect 4470 938 4478 941
rect 4470 832 4473 938
rect 4494 872 4497 1468
rect 4502 1378 4510 1381
rect 4486 868 4494 871
rect 4390 462 4393 478
rect 4406 202 4409 468
rect 4414 222 4417 718
rect 4424 603 4426 607
rect 4430 603 4433 607
rect 4438 603 4440 607
rect 4424 403 4426 407
rect 4430 403 4433 407
rect 4438 403 4440 407
rect 4424 203 4426 207
rect 4430 203 4433 207
rect 4438 203 4440 207
rect 4406 72 4409 198
rect 4430 112 4433 128
rect 4438 82 4441 108
rect 4446 82 4449 628
rect 4486 332 4489 868
rect 4502 802 4505 1378
rect 4514 1358 4518 1361
rect 4534 1262 4537 1418
rect 4542 1402 4545 2408
rect 4550 1952 4553 2688
rect 4558 2442 4561 3158
rect 4574 3152 4577 3318
rect 4558 2282 4561 2288
rect 4554 1948 4561 1951
rect 4558 1472 4561 1948
rect 4566 1612 4569 3148
rect 4574 3052 4577 3078
rect 4574 2792 4577 3048
rect 4582 2992 4585 3258
rect 4582 2772 4585 2908
rect 4578 2678 4582 2681
rect 4590 2562 4593 3878
rect 4606 3662 4609 3928
rect 4630 3762 4633 4238
rect 4638 4142 4641 4228
rect 4622 3748 4630 3751
rect 4598 2862 4601 3458
rect 4606 3162 4609 3658
rect 4606 3062 4609 3068
rect 4582 2252 4585 2258
rect 4566 1502 4569 1568
rect 4562 1418 4566 1421
rect 4574 1362 4577 1828
rect 4582 1682 4585 2048
rect 4590 1882 4593 1888
rect 4598 1702 4601 2778
rect 4614 2692 4617 3458
rect 4614 2582 4617 2588
rect 4614 2541 4617 2568
rect 4610 2538 4617 2541
rect 4614 2352 4617 2388
rect 4610 2248 4614 2251
rect 4622 2102 4625 3748
rect 4630 3642 4633 3668
rect 4646 3642 4649 4068
rect 4634 3548 4638 3551
rect 4654 3462 4657 4448
rect 4662 4122 4665 4528
rect 4670 4282 4673 4298
rect 4670 4172 4673 4278
rect 4630 3092 4633 3418
rect 4630 2461 4633 2718
rect 4630 2458 4638 2461
rect 4610 2058 4614 2061
rect 4606 1751 4609 2018
rect 4606 1748 4614 1751
rect 4594 1568 4598 1571
rect 4582 1382 4585 1558
rect 4598 1542 4601 1548
rect 4606 1362 4609 1738
rect 4614 1352 4617 1578
rect 4622 1571 4625 1998
rect 4630 1632 4633 2358
rect 4638 2142 4641 2438
rect 4638 2062 4641 2138
rect 4646 1652 4649 3048
rect 4654 2902 4657 3438
rect 4662 3382 4665 3548
rect 4670 2982 4673 3638
rect 4678 3462 4681 3748
rect 4686 3472 4689 4768
rect 4706 4558 4710 4561
rect 4726 4341 4729 4818
rect 4722 4338 4729 4341
rect 4734 4242 4737 4508
rect 4694 3842 4697 4158
rect 4734 4152 4737 4238
rect 4710 4112 4713 4118
rect 4678 3442 4681 3448
rect 4662 2742 4665 2968
rect 4658 2738 4662 2741
rect 4670 2191 4673 2978
rect 4686 2762 4689 3458
rect 4694 3022 4697 3638
rect 4702 3062 4705 3398
rect 4710 3052 4713 4108
rect 4686 2652 4689 2738
rect 4686 2362 4689 2398
rect 4694 2262 4697 3018
rect 4702 2962 4705 2978
rect 4718 2842 4721 3798
rect 4726 3362 4729 3978
rect 4670 2188 4681 2191
rect 4654 1632 4657 2148
rect 4678 2072 4681 2188
rect 4662 1792 4665 2058
rect 4670 2052 4673 2058
rect 4622 1568 4633 1571
rect 4662 1571 4665 1588
rect 4670 1582 4673 1848
rect 4678 1822 4681 2068
rect 4702 2012 4705 2738
rect 4710 2432 4713 2768
rect 4710 2222 4713 2378
rect 4718 2052 4721 2058
rect 4726 2002 4729 3148
rect 4734 2972 4737 4148
rect 4742 3222 4745 3488
rect 4750 3172 4753 4278
rect 4758 3972 4761 4968
rect 4758 3392 4761 3738
rect 4758 3142 4761 3388
rect 4742 2722 4745 3138
rect 4758 3052 4761 3108
rect 4758 2652 4761 2758
rect 4766 2682 4769 4738
rect 4774 3662 4777 3708
rect 4774 2662 4777 3658
rect 4782 2772 4785 4748
rect 4854 4462 4857 4688
rect 4862 4541 4865 4918
rect 4862 4538 4870 4541
rect 4834 4258 4838 4261
rect 4822 4252 4825 4258
rect 4806 4242 4809 4248
rect 4790 3271 4793 3428
rect 4790 3268 4798 3271
rect 4790 2852 4793 3188
rect 4806 3141 4809 3938
rect 4814 3262 4817 4218
rect 4822 3162 4825 3538
rect 4802 3138 4809 3141
rect 4786 2748 4793 2751
rect 4770 2658 4774 2661
rect 4746 2448 4753 2451
rect 4734 2442 4737 2448
rect 4750 2432 4753 2448
rect 4742 2071 4745 2268
rect 4758 2232 4761 2488
rect 4778 2448 4782 2451
rect 4790 2442 4793 2748
rect 4798 2592 4801 3138
rect 4818 2918 4822 2921
rect 4830 2882 4833 3348
rect 4838 3302 4841 4198
rect 4854 3822 4857 4238
rect 4846 3732 4849 3748
rect 4854 3372 4857 3818
rect 4842 3278 4846 3281
rect 4842 3248 4849 3251
rect 4846 3232 4849 3248
rect 4854 2922 4857 3358
rect 4870 3271 4873 3818
rect 4878 3512 4881 4268
rect 4886 4162 4889 4418
rect 4890 4158 4897 4161
rect 4886 3932 4889 3948
rect 4894 3942 4897 4158
rect 4894 3842 4897 3848
rect 4886 3292 4889 3638
rect 4862 3268 4873 3271
rect 4862 3252 4865 3268
rect 4870 3252 4873 3258
rect 4862 3232 4865 3238
rect 4870 3202 4873 3238
rect 4866 3148 4870 3151
rect 4862 2952 4865 3138
rect 4878 2962 4881 3268
rect 4886 3162 4889 3288
rect 4874 2938 4881 2941
rect 4830 2862 4833 2868
rect 4798 2452 4801 2478
rect 4766 2272 4769 2278
rect 4762 2128 4766 2131
rect 4738 2068 4745 2071
rect 4706 1958 4710 1961
rect 4710 1802 4713 1848
rect 4710 1762 4713 1798
rect 4702 1758 4710 1761
rect 4690 1658 4694 1661
rect 4658 1568 4665 1571
rect 4702 1572 4705 1758
rect 4718 1692 4721 1998
rect 4718 1662 4721 1688
rect 4622 1552 4625 1558
rect 4622 1502 4625 1508
rect 4622 1362 4625 1388
rect 4574 1281 4577 1288
rect 4570 1278 4577 1281
rect 4550 1151 4553 1178
rect 4546 1148 4553 1151
rect 4538 1068 4545 1071
rect 4534 1042 4537 1048
rect 4510 842 4513 948
rect 4494 622 4497 798
rect 4526 492 4529 678
rect 4534 482 4537 898
rect 4542 502 4545 1068
rect 4574 682 4577 1278
rect 4590 1132 4593 1188
rect 4590 852 4593 998
rect 4598 882 4601 1138
rect 4586 548 4590 551
rect 4538 278 4542 281
rect 4526 82 4529 228
rect 4246 58 4254 61
rect 4534 12 4537 278
rect 4550 232 4553 518
rect 4574 382 4577 548
rect 4598 422 4601 878
rect 4606 752 4609 1338
rect 4630 1062 4633 1568
rect 4638 1142 4641 1528
rect 4650 1338 4657 1341
rect 4646 1142 4649 1168
rect 4654 1132 4657 1338
rect 4614 692 4617 928
rect 4622 772 4625 948
rect 4606 642 4609 678
rect 4654 662 4657 668
rect 4662 582 4665 1568
rect 4694 1552 4697 1558
rect 4682 1258 4686 1261
rect 4670 1142 4673 1148
rect 4678 882 4681 1078
rect 4674 678 4678 681
rect 4598 402 4601 418
rect 4574 172 4577 378
rect 4582 272 4585 358
rect 4686 352 4689 418
rect 4686 182 4689 348
rect 4694 342 4697 1508
rect 4718 1392 4721 1518
rect 4718 1352 4721 1358
rect 4706 968 4710 971
rect 4726 812 4729 1778
rect 4734 1152 4737 1488
rect 4742 1421 4745 1518
rect 4742 1418 4750 1421
rect 4734 742 4737 1128
rect 4742 922 4745 1318
rect 4750 1132 4753 1388
rect 4766 1362 4769 1568
rect 4774 1422 4777 2418
rect 4782 1932 4785 2148
rect 4790 1852 4793 2358
rect 4758 1012 4761 1348
rect 4754 958 4758 961
rect 4766 752 4769 1108
rect 4774 1092 4777 1338
rect 4782 1042 4785 1468
rect 4710 622 4713 658
rect 4710 422 4713 618
rect 4702 348 4710 351
rect 4702 172 4705 348
rect 4574 72 4577 168
rect 4726 62 4729 688
rect 4734 552 4737 738
rect 4758 151 4761 508
rect 4754 148 4761 151
rect 4766 52 4769 578
rect 4774 252 4777 448
rect 4798 112 4801 2438
rect 4806 2262 4809 2338
rect 4814 2152 4817 2648
rect 4822 1882 4825 2858
rect 4830 2702 4833 2848
rect 4830 2672 4833 2698
rect 4838 2602 4841 2908
rect 4846 1902 4849 2858
rect 4854 1982 4857 2898
rect 4862 2712 4865 2918
rect 4878 2852 4881 2938
rect 4886 2862 4889 2868
rect 4870 1982 4873 2768
rect 4894 2762 4897 3838
rect 4878 2662 4881 2758
rect 4878 2242 4881 2548
rect 4886 2212 4889 2618
rect 4894 2382 4897 2718
rect 4854 1892 4857 1898
rect 4854 1832 4857 1858
rect 4854 1682 4857 1828
rect 4814 1461 4817 1578
rect 4810 1458 4817 1461
rect 4810 1418 4814 1421
rect 4806 1361 4809 1368
rect 4806 1358 4814 1361
rect 4814 912 4817 1278
rect 4814 762 4817 908
rect 4830 222 4833 1678
rect 4862 1652 4865 1968
rect 4894 1742 4897 2158
rect 4874 1658 4878 1661
rect 4862 1552 4865 1648
rect 4894 1222 4897 1468
rect 4894 1142 4897 1218
rect 4866 748 4870 751
rect 4838 462 4841 478
rect 4870 132 4873 608
rect 4830 92 4833 118
rect 4878 92 4881 918
rect 4886 692 4889 1118
rect 4894 842 4897 938
rect 4894 662 4897 818
rect 4890 658 4894 661
rect 4890 558 4894 561
rect 4890 478 4894 481
rect 4902 272 4905 5058
rect 4926 5052 4929 5058
rect 4910 5042 4913 5048
rect 5014 4942 5017 5038
rect 5146 5018 5150 5021
rect 4910 4472 4913 4938
rect 5006 4922 5009 4928
rect 4936 4903 4938 4907
rect 4942 4903 4945 4907
rect 4950 4903 4952 4907
rect 4926 4692 4929 4708
rect 4936 4703 4938 4707
rect 4942 4703 4945 4707
rect 4950 4703 4952 4707
rect 4910 3662 4913 4318
rect 4918 3962 4921 4588
rect 4936 4503 4938 4507
rect 4942 4503 4945 4507
rect 4950 4503 4952 4507
rect 4962 4478 4966 4481
rect 4926 4142 4929 4308
rect 4936 4303 4938 4307
rect 4942 4303 4945 4307
rect 4950 4303 4952 4307
rect 4936 4103 4938 4107
rect 4942 4103 4945 4107
rect 4950 4103 4952 4107
rect 4936 3903 4938 3907
rect 4942 3903 4945 3907
rect 4950 3903 4952 3907
rect 4926 3552 4929 3748
rect 4958 3722 4961 3918
rect 4936 3703 4938 3707
rect 4942 3703 4945 3707
rect 4950 3703 4952 3707
rect 4958 3692 4961 3718
rect 4950 3682 4953 3688
rect 4936 3503 4938 3507
rect 4942 3503 4945 3507
rect 4950 3503 4952 3507
rect 4958 3452 4961 3688
rect 4910 3272 4913 3278
rect 4910 3152 4913 3158
rect 4910 3082 4913 3088
rect 4910 2992 4913 3028
rect 4910 2752 4913 2758
rect 4918 2752 4921 3368
rect 4910 1252 4913 2748
rect 4918 2722 4921 2748
rect 4918 2382 4921 2698
rect 4926 2232 4929 3368
rect 4936 3303 4938 3307
rect 4942 3303 4945 3307
rect 4950 3303 4952 3307
rect 4936 3103 4938 3107
rect 4942 3103 4945 3107
rect 4950 3103 4952 3107
rect 4958 3062 4961 3448
rect 4966 3122 4969 3548
rect 4936 2903 4938 2907
rect 4942 2903 4945 2907
rect 4950 2903 4952 2907
rect 4950 2732 4953 2888
rect 4936 2703 4938 2707
rect 4942 2703 4945 2707
rect 4950 2703 4952 2707
rect 4936 2503 4938 2507
rect 4942 2503 4945 2507
rect 4950 2503 4952 2507
rect 4958 2352 4961 2878
rect 4966 2442 4969 2738
rect 4936 2303 4938 2307
rect 4942 2303 4945 2307
rect 4950 2303 4952 2307
rect 4966 2222 4969 2348
rect 4918 2112 4921 2148
rect 4936 2103 4938 2107
rect 4942 2103 4945 2107
rect 4950 2103 4952 2107
rect 4918 1362 4921 1938
rect 4936 1903 4938 1907
rect 4942 1903 4945 1907
rect 4950 1903 4952 1907
rect 4936 1703 4938 1707
rect 4942 1703 4945 1707
rect 4950 1703 4952 1707
rect 4926 1572 4929 1678
rect 4936 1503 4938 1507
rect 4942 1503 4945 1507
rect 4950 1503 4952 1507
rect 4930 1468 4934 1471
rect 4922 1338 4929 1341
rect 4910 1072 4913 1148
rect 4910 672 4913 1068
rect 4910 362 4913 668
rect 4918 572 4921 1248
rect 4926 1082 4929 1338
rect 4936 1303 4938 1307
rect 4942 1303 4945 1307
rect 4950 1303 4952 1307
rect 4934 1122 4937 1248
rect 4936 1103 4938 1107
rect 4942 1103 4945 1107
rect 4950 1103 4952 1107
rect 4930 958 4937 961
rect 4934 952 4937 958
rect 4936 903 4938 907
rect 4942 903 4945 907
rect 4950 903 4952 907
rect 4936 703 4938 707
rect 4942 703 4945 707
rect 4950 703 4952 707
rect 4930 678 4934 681
rect 4936 503 4938 507
rect 4942 503 4945 507
rect 4950 503 4952 507
rect 4930 478 4934 481
rect 4958 322 4961 1808
rect 4974 1682 4977 4788
rect 4994 4558 4998 4561
rect 4998 4532 5001 4538
rect 4982 3962 4985 4508
rect 4990 4172 4993 4498
rect 4998 3952 5001 4438
rect 5006 4282 5009 4808
rect 4986 3948 4990 3951
rect 4982 3852 4985 3938
rect 4990 3762 4993 3938
rect 4998 3872 5001 3928
rect 4998 3751 5001 3868
rect 4990 3748 5001 3751
rect 4982 3412 4985 3748
rect 4990 3402 4993 3748
rect 4998 3472 5001 3718
rect 5006 3591 5009 4168
rect 5014 3692 5017 4938
rect 5022 4918 5030 4921
rect 5022 4832 5025 4918
rect 5022 4262 5025 4638
rect 5030 4292 5033 4878
rect 5038 4382 5041 4748
rect 5046 4592 5049 4888
rect 5054 4861 5057 5018
rect 5066 4868 5070 4871
rect 5054 4858 5065 4861
rect 5022 3922 5025 3928
rect 5030 3872 5033 4278
rect 5038 3962 5041 4368
rect 5046 4072 5049 4578
rect 5054 4272 5057 4718
rect 5054 4262 5057 4268
rect 5042 3948 5046 3951
rect 5006 3588 5017 3591
rect 4982 3092 4985 3398
rect 4990 3202 4993 3378
rect 5006 3372 5009 3578
rect 4982 1982 4985 3048
rect 4990 2632 4993 3188
rect 5014 3132 5017 3588
rect 5002 2918 5006 2921
rect 5014 2762 5017 3118
rect 5022 3012 5025 3758
rect 5038 3662 5041 3848
rect 5046 3622 5049 3938
rect 5038 3232 5041 3488
rect 5038 3221 5041 3228
rect 5030 3218 5041 3221
rect 5022 2822 5025 2988
rect 4990 2162 4993 2598
rect 4994 2058 4998 2061
rect 5006 1932 5009 2648
rect 5014 2302 5017 2658
rect 5014 2052 5017 2168
rect 5022 2152 5025 2448
rect 5030 2392 5033 3218
rect 5046 3172 5049 3378
rect 5038 2732 5041 2938
rect 5038 2362 5041 2728
rect 5046 2692 5049 3158
rect 5030 2162 5033 2168
rect 5046 2132 5049 2668
rect 5054 2372 5057 3968
rect 5062 2822 5065 4858
rect 5062 2722 5065 2808
rect 4982 1671 4985 1848
rect 4974 1668 4985 1671
rect 4966 1372 4969 1378
rect 4966 1122 4969 1358
rect 4974 952 4977 1668
rect 5006 1532 5009 1678
rect 4966 452 4969 748
rect 4974 742 4977 948
rect 4982 932 4985 1138
rect 4974 342 4977 628
rect 4926 282 4929 318
rect 4936 303 4938 307
rect 4942 303 4945 307
rect 4950 303 4952 307
rect 4890 128 4894 131
rect 4936 103 4938 107
rect 4942 103 4945 107
rect 4950 103 4952 107
rect 4910 81 4913 88
rect 4910 78 4918 81
rect 4822 72 4825 78
rect 4958 62 4961 278
rect 4982 162 4985 868
rect 4990 862 4993 1138
rect 4990 742 4993 748
rect 4990 472 4993 478
rect 4998 292 5001 1428
rect 5006 692 5009 758
rect 5006 342 5009 668
rect 5014 462 5017 738
rect 5022 282 5025 1968
rect 5030 1772 5033 2018
rect 5038 1882 5041 2068
rect 5046 2058 5054 2061
rect 5038 1862 5041 1868
rect 5030 1552 5033 1768
rect 5030 1322 5033 1428
rect 5030 652 5033 838
rect 5038 822 5041 1848
rect 5046 1532 5049 2058
rect 5046 732 5049 1398
rect 5054 1142 5057 1888
rect 5062 1752 5065 2358
rect 5070 1912 5073 4848
rect 5078 3192 5081 4768
rect 5086 2842 5089 4918
rect 5094 4132 5097 4928
rect 5102 4352 5105 4698
rect 5094 3442 5097 4118
rect 5102 3222 5105 4338
rect 5110 4002 5113 4868
rect 5118 4362 5121 4968
rect 5110 3772 5113 3988
rect 5118 3952 5121 4348
rect 5126 4102 5129 4938
rect 5134 4122 5137 4858
rect 5142 4422 5145 4658
rect 5150 4632 5153 4638
rect 5150 4472 5153 4548
rect 5142 4242 5145 4378
rect 5150 4112 5153 4358
rect 5158 4302 5161 4688
rect 5166 4552 5169 5068
rect 5178 4718 5182 4721
rect 5166 4282 5169 4528
rect 5174 4322 5177 4708
rect 5182 4462 5185 4548
rect 5182 4452 5185 4458
rect 5178 4308 5182 4311
rect 5126 3988 5134 3991
rect 5126 3822 5129 3988
rect 5094 2832 5097 3178
rect 5086 2722 5089 2768
rect 5086 2682 5089 2698
rect 5078 2252 5081 2638
rect 5086 2592 5089 2678
rect 5086 2252 5089 2518
rect 5070 1551 5073 1568
rect 5066 1548 5073 1551
rect 5062 1062 5065 1488
rect 5070 1232 5073 1348
rect 5046 682 5049 728
rect 5042 658 5046 661
rect 5038 462 5041 488
rect 5054 462 5057 748
rect 5062 672 5065 1058
rect 5070 742 5073 958
rect 4998 262 5001 268
rect 5062 262 5065 668
rect 5070 662 5073 668
rect 5078 622 5081 2058
rect 5086 1232 5089 2238
rect 5094 2172 5097 2818
rect 5102 2552 5105 3208
rect 5110 3102 5113 3738
rect 5118 3692 5121 3798
rect 5130 3758 5134 3761
rect 5134 3722 5137 3728
rect 5130 3708 5137 3711
rect 5118 3152 5121 3678
rect 5126 3512 5129 3698
rect 5126 3462 5129 3468
rect 5134 3442 5137 3708
rect 5110 2852 5113 3018
rect 5102 2392 5105 2428
rect 5110 2192 5113 2828
rect 5118 2562 5121 2978
rect 5094 1962 5097 2158
rect 5094 1922 5097 1928
rect 5102 1882 5105 2098
rect 5094 1742 5097 1758
rect 5102 1722 5105 1858
rect 5110 1442 5113 2108
rect 5118 1892 5121 2548
rect 5126 2312 5129 3358
rect 5134 3212 5137 3338
rect 5134 2992 5137 3188
rect 5086 812 5089 1198
rect 5094 1122 5097 1348
rect 5102 1282 5105 1338
rect 5094 852 5097 1108
rect 5086 772 5089 808
rect 5102 802 5105 1208
rect 5110 1042 5113 1428
rect 5118 1322 5121 1878
rect 5126 1732 5129 2188
rect 5126 1362 5129 1718
rect 5118 1052 5121 1148
rect 5102 752 5105 798
rect 5094 292 5097 498
rect 5102 492 5105 728
rect 5110 512 5113 1008
rect 5118 762 5121 1048
rect 5126 982 5129 1308
rect 5134 1142 5137 2968
rect 5142 2862 5145 4098
rect 5158 4002 5161 4208
rect 5150 2972 5153 3838
rect 5158 3702 5161 3958
rect 5166 3942 5169 4048
rect 5166 3862 5169 3928
rect 5174 3872 5177 4298
rect 5182 4112 5185 4278
rect 5182 4072 5185 4078
rect 5190 3861 5193 4888
rect 5198 4332 5201 4338
rect 5198 4012 5201 4318
rect 5182 3858 5193 3861
rect 5142 2492 5145 2848
rect 5150 2272 5153 2948
rect 5158 2382 5161 3688
rect 5166 2892 5169 3708
rect 5174 3562 5177 3678
rect 5174 2812 5177 3538
rect 5166 2572 5169 2748
rect 5174 2561 5177 2798
rect 5166 2558 5177 2561
rect 5142 2142 5145 2248
rect 5018 258 5022 261
rect 5062 232 5065 258
rect 5082 188 5086 191
rect 4982 42 4985 158
rect 5034 78 5038 81
rect 5126 62 5129 788
rect 5134 572 5137 578
rect 5142 72 5145 1918
rect 5150 1142 5153 1498
rect 5158 1432 5161 2348
rect 5166 1892 5169 2558
rect 5174 2322 5177 2338
rect 5182 2192 5185 3858
rect 5190 3742 5193 3848
rect 5190 3032 5193 3738
rect 5198 3662 5201 3858
rect 5198 3172 5201 3518
rect 5190 2832 5193 3018
rect 5198 2921 5201 3128
rect 5206 2931 5209 5078
rect 5230 4792 5233 4918
rect 5238 4702 5241 5058
rect 5214 4132 5217 4558
rect 5214 3272 5217 4108
rect 5214 2952 5217 3178
rect 5206 2928 5217 2931
rect 5198 2918 5209 2921
rect 5198 2822 5201 2898
rect 5206 2862 5209 2918
rect 5190 2562 5193 2568
rect 5190 2502 5193 2508
rect 5182 2152 5185 2168
rect 5182 2132 5185 2138
rect 5166 1462 5169 1668
rect 5158 1082 5161 1418
rect 5166 1172 5169 1348
rect 5174 1161 5177 1658
rect 5182 1502 5185 2108
rect 5190 2072 5193 2488
rect 5198 2222 5201 2808
rect 5206 1711 5209 2848
rect 5198 1708 5209 1711
rect 5182 1462 5185 1478
rect 5182 1262 5185 1338
rect 5170 1158 5177 1161
rect 5190 1172 5193 1468
rect 5198 1451 5201 1708
rect 5206 1692 5209 1698
rect 5198 1448 5209 1451
rect 5198 1312 5201 1438
rect 5190 1162 5193 1168
rect 5166 1152 5169 1158
rect 5150 352 5153 958
rect 5158 332 5161 1068
rect 5166 392 5169 1088
rect 5174 532 5177 1138
rect 5182 872 5185 918
rect 5182 862 5185 868
rect 5182 732 5185 768
rect 5182 492 5185 648
rect 5170 58 5174 61
rect 5182 52 5185 458
rect 5190 362 5193 978
rect 5198 382 5201 1168
rect 5206 482 5209 1448
rect 5214 962 5217 2928
rect 5222 2852 5225 4418
rect 5230 3422 5233 4588
rect 5246 4342 5249 4878
rect 5254 4862 5257 4868
rect 5246 3872 5249 4318
rect 5242 3858 5246 3861
rect 5242 3558 5249 3561
rect 5246 3522 5249 3558
rect 5230 3122 5233 3128
rect 5230 3022 5233 3088
rect 5222 2112 5225 2838
rect 5222 1522 5225 2098
rect 5230 1311 5233 3008
rect 5238 2552 5241 3458
rect 5246 2652 5249 3508
rect 5254 2942 5257 4848
rect 5246 2552 5249 2558
rect 5238 2132 5241 2538
rect 5254 2522 5257 2938
rect 5246 2332 5249 2338
rect 5262 2291 5265 4878
rect 5270 3932 5273 4838
rect 5278 4172 5281 4818
rect 5270 3642 5273 3928
rect 5278 3682 5281 3688
rect 5270 2322 5273 3558
rect 5258 2288 5265 2291
rect 5246 2122 5249 2218
rect 5254 1872 5257 2138
rect 5238 1692 5241 1858
rect 5238 1532 5241 1678
rect 5222 1308 5233 1311
rect 5214 322 5217 948
rect 5202 288 5206 291
rect 5214 282 5217 308
rect 5222 262 5225 1308
rect 5230 462 5233 1188
rect 5238 902 5241 1518
rect 5230 172 5233 438
rect 5238 312 5241 888
rect 5246 292 5249 1178
rect 5254 922 5257 1858
rect 5262 1662 5265 2208
rect 5254 372 5257 908
rect 5262 822 5265 1568
rect 5270 1022 5273 2308
rect 5278 2202 5281 3528
rect 5286 2822 5289 4808
rect 5294 3272 5297 3538
rect 5294 3252 5297 3258
rect 5294 2892 5297 2948
rect 5286 2412 5289 2568
rect 5286 2372 5289 2388
rect 5294 2352 5297 2418
rect 5278 2062 5281 2068
rect 5270 992 5273 998
rect 5278 982 5281 1948
rect 5286 1162 5289 2168
rect 5294 1932 5297 2318
rect 5302 2272 5305 4788
rect 5302 2242 5305 2248
rect 5262 342 5265 768
rect 5270 732 5273 758
rect 5270 472 5273 478
rect 5278 322 5281 968
rect 5286 402 5289 1148
rect 5294 532 5297 1908
rect 5286 282 5289 318
rect 5302 272 5305 2228
rect 5246 152 5249 158
rect 5274 148 5278 151
rect 5262 132 5265 138
rect 5226 68 5230 71
rect 328 3 330 7
rect 334 3 337 7
rect 342 3 344 7
rect 1352 3 1354 7
rect 1358 3 1361 7
rect 1366 3 1368 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2398 3 2400 7
rect 3400 3 3402 7
rect 3406 3 3409 7
rect 3414 3 3416 7
rect 4424 3 4426 7
rect 4430 3 4433 7
rect 4438 3 4440 7
<< m5contact >>
rect 850 5103 854 5107
rect 857 5103 858 5107
rect 858 5103 861 5107
rect 1874 5103 1878 5107
rect 1881 5103 1882 5107
rect 1882 5103 1885 5107
rect 2890 5103 2894 5107
rect 2897 5103 2898 5107
rect 2898 5103 2901 5107
rect 3922 5103 3926 5107
rect 3929 5103 3930 5107
rect 3930 5103 3933 5107
rect 4938 5103 4942 5107
rect 4945 5103 4946 5107
rect 4946 5103 4949 5107
rect 166 5058 170 5062
rect 198 5058 202 5062
rect 330 5003 334 5007
rect 337 5003 338 5007
rect 338 5003 341 5007
rect 190 4948 194 4952
rect 198 4928 202 4932
rect 246 4848 250 4852
rect 330 4803 334 4807
rect 337 4803 338 4807
rect 338 4803 341 4807
rect 470 4958 474 4962
rect 542 4878 546 4882
rect 430 4758 434 4762
rect 134 4348 138 4352
rect 110 3838 114 3842
rect 54 3748 58 3752
rect 86 3748 90 3752
rect 206 4278 210 4282
rect 330 4603 334 4607
rect 337 4603 338 4607
rect 338 4603 341 4607
rect 330 4403 334 4407
rect 337 4403 338 4407
rect 338 4403 341 4407
rect 318 4328 322 4332
rect 214 3838 218 3842
rect 374 4538 378 4542
rect 358 4248 362 4252
rect 350 4228 354 4232
rect 330 4203 334 4207
rect 337 4203 338 4207
rect 338 4203 341 4207
rect 446 4558 450 4562
rect 438 4538 442 4542
rect 486 4338 490 4342
rect 382 4178 386 4182
rect 330 4003 334 4007
rect 337 4003 338 4007
rect 338 4003 341 4007
rect 526 4178 530 4182
rect 330 3803 334 3807
rect 337 3803 338 3807
rect 338 3803 341 3807
rect 150 3568 154 3572
rect 46 2858 50 2862
rect 86 2668 90 2672
rect 118 2668 122 2672
rect 330 3603 334 3607
rect 337 3603 338 3607
rect 338 3603 341 3607
rect 462 3838 466 3842
rect 702 4878 706 4882
rect 638 4758 642 4762
rect 638 4728 642 4732
rect 582 4608 586 4612
rect 598 4558 602 4562
rect 742 4958 746 4962
rect 774 4948 778 4952
rect 790 4858 794 4862
rect 734 4848 738 4852
rect 734 4768 738 4772
rect 694 4618 698 4622
rect 702 4338 706 4342
rect 566 4328 570 4332
rect 614 4278 618 4282
rect 550 4078 554 4082
rect 638 4268 642 4272
rect 598 4258 602 4262
rect 646 4248 650 4252
rect 574 3978 578 3982
rect 598 3978 602 3982
rect 718 4458 722 4462
rect 870 4928 874 4932
rect 850 4903 854 4907
rect 857 4903 858 4907
rect 858 4903 861 4907
rect 870 4858 874 4862
rect 910 4728 914 4732
rect 850 4703 854 4707
rect 857 4703 858 4707
rect 858 4703 861 4707
rect 850 4503 854 4507
rect 857 4503 858 4507
rect 858 4503 861 4507
rect 886 4448 890 4452
rect 798 4348 802 4352
rect 850 4303 854 4307
rect 857 4303 858 4307
rect 858 4303 861 4307
rect 734 4268 738 4272
rect 782 4258 786 4262
rect 774 4248 778 4252
rect 830 4248 834 4252
rect 814 4228 818 4232
rect 1070 4458 1074 4462
rect 1354 5003 1358 5007
rect 1361 5003 1362 5007
rect 1362 5003 1365 5007
rect 1462 4948 1466 4952
rect 1150 4548 1154 4552
rect 850 4103 854 4107
rect 857 4103 858 4107
rect 858 4103 861 4107
rect 630 3668 634 3672
rect 462 3588 466 3592
rect 398 3448 402 3452
rect 330 3403 334 3407
rect 337 3403 338 3407
rect 338 3403 341 3407
rect 262 2858 266 2862
rect 262 2748 266 2752
rect 214 2698 218 2702
rect 158 2148 162 2152
rect 30 1818 34 1822
rect 54 718 58 722
rect 214 1518 218 1522
rect 294 2268 298 2272
rect 470 3528 474 3532
rect 566 3528 570 3532
rect 510 3418 514 3422
rect 566 3358 570 3362
rect 430 3338 434 3342
rect 446 3328 450 3332
rect 470 3228 474 3232
rect 406 3218 410 3222
rect 330 3203 334 3207
rect 337 3203 338 3207
rect 338 3203 341 3207
rect 330 3003 334 3007
rect 337 3003 338 3007
rect 338 3003 341 3007
rect 358 2818 362 2822
rect 330 2803 334 2807
rect 337 2803 338 2807
rect 338 2803 341 2807
rect 310 2698 314 2702
rect 330 2603 334 2607
rect 337 2603 338 2607
rect 338 2603 341 2607
rect 330 2403 334 2407
rect 337 2403 338 2407
rect 338 2403 341 2407
rect 310 2278 314 2282
rect 238 1258 242 1262
rect 318 2258 322 2262
rect 330 2203 334 2207
rect 337 2203 338 2207
rect 338 2203 341 2207
rect 330 2003 334 2007
rect 337 2003 338 2007
rect 338 2003 341 2007
rect 398 2668 402 2672
rect 374 2268 378 2272
rect 318 1818 322 1822
rect 206 538 210 542
rect 330 1803 334 1807
rect 337 1803 338 1807
rect 338 1803 341 1807
rect 330 1603 334 1607
rect 337 1603 338 1607
rect 338 1603 341 1607
rect 590 3268 594 3272
rect 590 3128 594 3132
rect 454 2888 458 2892
rect 494 2688 498 2692
rect 430 2428 434 2432
rect 342 1438 346 1442
rect 330 1403 334 1407
rect 337 1403 338 1407
rect 338 1403 341 1407
rect 330 1203 334 1207
rect 337 1203 338 1207
rect 338 1203 341 1207
rect 330 1003 334 1007
rect 337 1003 338 1007
rect 338 1003 341 1007
rect 318 938 322 942
rect 150 258 154 262
rect 262 258 266 262
rect 414 1558 418 1562
rect 406 1538 410 1542
rect 406 1458 410 1462
rect 398 1348 402 1352
rect 406 1268 410 1272
rect 422 1348 426 1352
rect 510 2848 514 2852
rect 598 2878 602 2882
rect 526 2678 530 2682
rect 550 2668 554 2672
rect 582 2488 586 2492
rect 534 2368 538 2372
rect 518 2358 522 2362
rect 550 2348 554 2352
rect 454 2338 458 2342
rect 542 2078 546 2082
rect 510 2048 514 2052
rect 454 1578 458 1582
rect 330 803 334 807
rect 337 803 338 807
rect 338 803 341 807
rect 438 1248 442 1252
rect 414 728 418 732
rect 470 1058 474 1062
rect 478 988 482 992
rect 330 603 334 607
rect 337 603 338 607
rect 338 603 341 607
rect 342 558 346 562
rect 330 403 334 407
rect 337 403 338 407
rect 338 403 341 407
rect 334 348 338 352
rect 330 203 334 207
rect 337 203 338 207
rect 338 203 341 207
rect 558 2228 562 2232
rect 566 1168 570 1172
rect 590 1938 594 1942
rect 606 2748 610 2752
rect 718 3658 722 3662
rect 974 4028 978 4032
rect 934 3918 938 3922
rect 850 3903 854 3907
rect 857 3903 858 3907
rect 858 3903 861 3907
rect 966 3858 970 3862
rect 918 3728 922 3732
rect 850 3703 854 3707
rect 857 3703 858 3707
rect 858 3703 861 3707
rect 750 3648 754 3652
rect 782 3538 786 3542
rect 646 3468 650 3472
rect 862 3528 866 3532
rect 850 3503 854 3507
rect 857 3503 858 3507
rect 858 3503 861 3507
rect 654 3428 658 3432
rect 766 3358 770 3362
rect 734 3318 738 3322
rect 726 3258 730 3262
rect 638 2688 642 2692
rect 622 2608 626 2612
rect 654 2528 658 2532
rect 662 2368 666 2372
rect 662 2188 666 2192
rect 678 2938 682 2942
rect 718 2868 722 2872
rect 702 2838 706 2842
rect 718 2758 722 2762
rect 710 2678 714 2682
rect 702 2468 706 2472
rect 694 2348 698 2352
rect 622 2048 626 2052
rect 606 1758 610 1762
rect 598 1528 602 1532
rect 654 1938 658 1942
rect 662 1938 666 1942
rect 646 1878 650 1882
rect 630 1548 634 1552
rect 662 1548 666 1552
rect 638 1538 642 1542
rect 614 1458 618 1462
rect 590 978 594 982
rect 718 2338 722 2342
rect 710 1858 714 1862
rect 694 1828 698 1832
rect 750 3268 754 3272
rect 750 2868 754 2872
rect 734 2818 738 2822
rect 734 2758 738 2762
rect 742 2368 746 2372
rect 734 2168 738 2172
rect 798 3348 802 3352
rect 790 2948 794 2952
rect 782 2798 786 2802
rect 758 2598 762 2602
rect 758 2268 762 2272
rect 710 1768 714 1772
rect 702 1528 706 1532
rect 686 1438 690 1442
rect 678 1288 682 1292
rect 718 1548 722 1552
rect 782 2058 786 2062
rect 814 2888 818 2892
rect 806 2868 810 2872
rect 850 3303 854 3307
rect 857 3303 858 3307
rect 858 3303 861 3307
rect 838 3128 842 3132
rect 850 3103 854 3107
rect 857 3103 858 3107
rect 858 3103 861 3107
rect 830 2778 834 2782
rect 850 2903 854 2907
rect 857 2903 858 2907
rect 858 2903 861 2907
rect 998 3818 1002 3822
rect 894 3458 898 3462
rect 886 3348 890 3352
rect 886 2738 890 2742
rect 850 2703 854 2707
rect 857 2703 858 2707
rect 858 2703 861 2707
rect 850 2503 854 2507
rect 857 2503 858 2507
rect 858 2503 861 2507
rect 854 2468 858 2472
rect 814 2288 818 2292
rect 798 2268 802 2272
rect 758 1758 762 1762
rect 614 868 618 872
rect 582 858 586 862
rect 574 718 578 722
rect 702 948 706 952
rect 782 1818 786 1822
rect 790 1468 794 1472
rect 798 1288 802 1292
rect 494 618 498 622
rect 534 588 538 592
rect 670 548 674 552
rect 678 378 682 382
rect 850 2303 854 2307
rect 857 2303 858 2307
rect 858 2303 861 2307
rect 838 2238 842 2242
rect 822 1948 826 1952
rect 850 2103 854 2107
rect 857 2103 858 2107
rect 858 2103 861 2107
rect 850 1903 854 1907
rect 857 1903 858 1907
rect 858 1903 861 1907
rect 846 1868 850 1872
rect 850 1703 854 1707
rect 857 1703 858 1707
rect 858 1703 861 1707
rect 850 1503 854 1507
rect 857 1503 858 1507
rect 858 1503 861 1507
rect 910 3088 914 3092
rect 894 2508 898 2512
rect 878 2448 882 2452
rect 894 2418 898 2422
rect 902 2408 906 2412
rect 902 2068 906 2072
rect 870 1328 874 1332
rect 850 1303 854 1307
rect 857 1303 858 1307
rect 858 1303 861 1307
rect 854 1268 858 1272
rect 838 1158 842 1162
rect 850 1103 854 1107
rect 857 1103 858 1107
rect 858 1103 861 1107
rect 814 958 818 962
rect 806 468 810 472
rect 798 348 802 352
rect 814 368 818 372
rect 846 978 850 982
rect 850 903 854 907
rect 857 903 858 907
rect 858 903 861 907
rect 850 703 854 707
rect 857 703 858 707
rect 858 703 861 707
rect 878 698 882 702
rect 870 688 874 692
rect 850 503 854 507
rect 857 503 858 507
rect 858 503 861 507
rect 850 303 854 307
rect 857 303 858 307
rect 858 303 861 307
rect 926 3158 930 3162
rect 942 3138 946 3142
rect 966 2918 970 2922
rect 942 2758 946 2762
rect 974 2748 978 2752
rect 934 2508 938 2512
rect 934 2358 938 2362
rect 918 2348 922 2352
rect 934 2338 938 2342
rect 974 2428 978 2432
rect 974 2268 978 2272
rect 926 1668 930 1672
rect 918 1188 922 1192
rect 910 938 914 942
rect 950 2148 954 2152
rect 950 1998 954 2002
rect 990 2258 994 2262
rect 1022 3528 1026 3532
rect 1014 3328 1018 3332
rect 1062 3898 1066 3902
rect 1086 3868 1090 3872
rect 1062 3708 1066 3712
rect 1118 3658 1122 3662
rect 1054 3638 1058 3642
rect 1190 4448 1194 4452
rect 1354 4803 1358 4807
rect 1361 4803 1362 4807
rect 1362 4803 1365 4807
rect 1454 4748 1458 4752
rect 1354 4603 1358 4607
rect 1361 4603 1362 4607
rect 1362 4603 1365 4607
rect 1782 5048 1786 5052
rect 2386 5003 2390 5007
rect 2393 5003 2394 5007
rect 2394 5003 2397 5007
rect 1726 4948 1730 4952
rect 1874 4903 1878 4907
rect 1881 4903 1882 4907
rect 1882 4903 1885 4907
rect 1358 4558 1362 4562
rect 1278 4138 1282 4142
rect 1294 4118 1298 4122
rect 1166 3878 1170 3882
rect 1182 3868 1186 3872
rect 1038 2948 1042 2952
rect 1038 2788 1042 2792
rect 1046 2768 1050 2772
rect 1006 2438 1010 2442
rect 1014 2278 1018 2282
rect 1006 2128 1010 2132
rect 1094 3018 1098 3022
rect 1086 2908 1090 2912
rect 1174 3558 1178 3562
rect 1174 3488 1178 3492
rect 1150 3338 1154 3342
rect 1142 3308 1146 3312
rect 1134 3128 1138 3132
rect 1102 2798 1106 2802
rect 1102 2678 1106 2682
rect 1222 3888 1226 3892
rect 1238 3878 1242 3882
rect 1254 3738 1258 3742
rect 1214 3678 1218 3682
rect 1198 3448 1202 3452
rect 1182 3148 1186 3152
rect 1174 2948 1178 2952
rect 1166 2888 1170 2892
rect 1110 2608 1114 2612
rect 1054 2248 1058 2252
rect 1038 2118 1042 2122
rect 974 1568 978 1572
rect 998 1488 1002 1492
rect 982 1388 986 1392
rect 966 1268 970 1272
rect 958 1258 962 1262
rect 950 968 954 972
rect 942 878 946 882
rect 934 868 938 872
rect 918 818 922 822
rect 934 728 938 732
rect 950 528 954 532
rect 902 478 906 482
rect 982 988 986 992
rect 998 1088 1002 1092
rect 998 758 1002 762
rect 1014 1168 1018 1172
rect 1022 938 1026 942
rect 1022 858 1026 862
rect 1022 568 1026 572
rect 990 338 994 342
rect 1102 2308 1106 2312
rect 1062 1578 1066 1582
rect 1102 1898 1106 1902
rect 1102 1728 1106 1732
rect 1094 948 1098 952
rect 1094 928 1098 932
rect 1182 2718 1186 2722
rect 1150 2688 1154 2692
rect 1118 2568 1122 2572
rect 1134 2338 1138 2342
rect 1118 1908 1122 1912
rect 1126 1888 1130 1892
rect 1142 1868 1146 1872
rect 1110 1538 1114 1542
rect 1118 1528 1122 1532
rect 1166 2348 1170 2352
rect 1222 3068 1226 3072
rect 1190 2308 1194 2312
rect 1182 2258 1186 2262
rect 1166 2148 1170 2152
rect 1158 1838 1162 1842
rect 1142 1668 1146 1672
rect 1174 2078 1178 2082
rect 1190 2108 1194 2112
rect 1174 2018 1178 2022
rect 1166 1448 1170 1452
rect 1214 2338 1218 2342
rect 1286 3918 1290 3922
rect 1278 3728 1282 3732
rect 1246 3668 1250 3672
rect 1270 3458 1274 3462
rect 1246 3368 1250 3372
rect 1238 2548 1242 2552
rect 1230 2438 1234 2442
rect 1238 2278 1242 2282
rect 1254 2878 1258 2882
rect 1262 2578 1266 2582
rect 1318 3868 1322 3872
rect 1334 3628 1338 3632
rect 1326 3338 1330 3342
rect 1354 4403 1358 4407
rect 1361 4403 1362 4407
rect 1362 4403 1365 4407
rect 1454 4368 1458 4372
rect 1462 4288 1466 4292
rect 1354 4203 1358 4207
rect 1361 4203 1362 4207
rect 1362 4203 1365 4207
rect 1478 4148 1482 4152
rect 1354 4003 1358 4007
rect 1361 4003 1362 4007
rect 1362 4003 1365 4007
rect 1350 3868 1354 3872
rect 1446 4038 1450 4042
rect 1354 3803 1358 3807
rect 1361 3803 1362 3807
rect 1362 3803 1365 3807
rect 1350 3688 1354 3692
rect 1414 3828 1418 3832
rect 1354 3603 1358 3607
rect 1361 3603 1362 3607
rect 1362 3603 1365 3607
rect 1310 3078 1314 3082
rect 1294 2988 1298 2992
rect 1278 2898 1282 2902
rect 1286 2858 1290 2862
rect 1278 2348 1282 2352
rect 1270 2318 1274 2322
rect 1246 2258 1250 2262
rect 1222 2138 1226 2142
rect 1230 1988 1234 1992
rect 1134 1078 1138 1082
rect 1166 1018 1170 1022
rect 1118 958 1122 962
rect 1174 958 1178 962
rect 1126 948 1130 952
rect 1062 788 1066 792
rect 1190 1228 1194 1232
rect 1118 668 1122 672
rect 1222 1738 1226 1742
rect 1206 1628 1210 1632
rect 1238 1588 1242 1592
rect 1230 1548 1234 1552
rect 1230 1528 1234 1532
rect 1214 1358 1218 1362
rect 1222 1328 1226 1332
rect 1262 1518 1266 1522
rect 1278 1468 1282 1472
rect 1270 1458 1274 1462
rect 1278 1268 1282 1272
rect 1254 1038 1258 1042
rect 1246 858 1250 862
rect 1246 818 1250 822
rect 1222 758 1226 762
rect 1262 558 1266 562
rect 1302 2848 1306 2852
rect 1318 2848 1322 2852
rect 1334 3058 1338 3062
rect 1326 2638 1330 2642
rect 1326 2588 1330 2592
rect 1354 3403 1358 3407
rect 1361 3403 1362 3407
rect 1362 3403 1365 3407
rect 1354 3203 1358 3207
rect 1361 3203 1362 3207
rect 1362 3203 1365 3207
rect 1406 3168 1410 3172
rect 1406 3128 1410 3132
rect 1354 3003 1358 3007
rect 1361 3003 1362 3007
rect 1362 3003 1365 3007
rect 1374 2918 1378 2922
rect 1354 2803 1358 2807
rect 1361 2803 1362 2807
rect 1362 2803 1365 2807
rect 1342 2628 1346 2632
rect 1354 2603 1358 2607
rect 1361 2603 1362 2607
rect 1362 2603 1365 2607
rect 1614 4748 1618 4752
rect 1718 4748 1722 4752
rect 1678 4268 1682 4272
rect 1670 4258 1674 4262
rect 1454 3998 1458 4002
rect 1422 3738 1426 3742
rect 1430 3258 1434 3262
rect 1454 3438 1458 3442
rect 1534 3728 1538 3732
rect 1526 3558 1530 3562
rect 1510 3438 1514 3442
rect 1462 3248 1466 3252
rect 1470 3218 1474 3222
rect 1438 3088 1442 3092
rect 1430 2708 1434 2712
rect 1414 2518 1418 2522
rect 1342 2408 1346 2412
rect 1354 2403 1358 2407
rect 1361 2403 1362 2407
rect 1362 2403 1365 2407
rect 1390 2398 1394 2402
rect 1302 2258 1306 2262
rect 1302 2158 1306 2162
rect 1374 2288 1378 2292
rect 1334 2178 1338 2182
rect 1326 2068 1330 2072
rect 1366 2218 1370 2222
rect 1354 2203 1358 2207
rect 1361 2203 1362 2207
rect 1362 2203 1365 2207
rect 1398 2338 1402 2342
rect 1430 2358 1434 2362
rect 1422 2328 1426 2332
rect 1382 2058 1386 2062
rect 1354 2003 1358 2007
rect 1361 2003 1362 2007
rect 1362 2003 1365 2007
rect 1374 1908 1378 1912
rect 1374 1808 1378 1812
rect 1354 1803 1358 1807
rect 1361 1803 1362 1807
rect 1362 1803 1365 1807
rect 1354 1603 1358 1607
rect 1361 1603 1362 1607
rect 1362 1603 1365 1607
rect 1382 1798 1386 1802
rect 1462 3138 1466 3142
rect 1454 3048 1458 3052
rect 1494 3238 1498 3242
rect 1542 3518 1546 3522
rect 1534 3508 1538 3512
rect 1550 3408 1554 3412
rect 1534 3308 1538 3312
rect 1534 3248 1538 3252
rect 1494 3128 1498 3132
rect 1462 2968 1466 2972
rect 1478 2868 1482 2872
rect 1446 2598 1450 2602
rect 1406 2058 1410 2062
rect 1422 2038 1426 2042
rect 1422 1958 1426 1962
rect 1414 1748 1418 1752
rect 1422 1668 1426 1672
rect 1398 1648 1402 1652
rect 1354 1403 1358 1407
rect 1361 1403 1362 1407
rect 1362 1403 1365 1407
rect 1310 1208 1314 1212
rect 1326 1158 1330 1162
rect 1278 558 1282 562
rect 1294 538 1298 542
rect 1294 438 1298 442
rect 1354 1203 1358 1207
rect 1361 1203 1362 1207
rect 1362 1203 1365 1207
rect 1354 1003 1358 1007
rect 1361 1003 1362 1007
rect 1362 1003 1365 1007
rect 1354 803 1358 807
rect 1361 803 1362 807
rect 1362 803 1365 807
rect 1430 1598 1434 1602
rect 1414 1578 1418 1582
rect 1414 1478 1418 1482
rect 1406 1268 1410 1272
rect 1414 958 1418 962
rect 1382 698 1386 702
rect 1374 668 1378 672
rect 1354 603 1358 607
rect 1361 603 1362 607
rect 1362 603 1365 607
rect 1342 588 1346 592
rect 1430 1288 1434 1292
rect 1462 2568 1466 2572
rect 1470 2418 1474 2422
rect 1454 2388 1458 2392
rect 1446 1948 1450 1952
rect 1462 2188 1466 2192
rect 1518 3108 1522 3112
rect 1502 2728 1506 2732
rect 1502 2468 1506 2472
rect 1486 2288 1490 2292
rect 1478 2218 1482 2222
rect 1486 2208 1490 2212
rect 1486 2128 1490 2132
rect 1462 1968 1466 1972
rect 1462 1718 1466 1722
rect 1502 2008 1506 2012
rect 1478 1688 1482 1692
rect 1470 1638 1474 1642
rect 1446 1468 1450 1472
rect 1542 2848 1546 2852
rect 1526 2578 1530 2582
rect 1518 2498 1522 2502
rect 1534 2508 1538 2512
rect 1606 3748 1610 3752
rect 1574 3358 1578 3362
rect 1622 3738 1626 3742
rect 1630 3628 1634 3632
rect 1638 3578 1642 3582
rect 1630 3568 1634 3572
rect 1614 3528 1618 3532
rect 1622 3518 1626 3522
rect 1574 3318 1578 3322
rect 1582 3278 1586 3282
rect 1566 3088 1570 3092
rect 1598 3058 1602 3062
rect 1558 2988 1562 2992
rect 1558 2858 1562 2862
rect 1590 2898 1594 2902
rect 1582 2828 1586 2832
rect 1558 2808 1562 2812
rect 1558 2778 1562 2782
rect 1566 2708 1570 2712
rect 1558 2678 1562 2682
rect 1558 2478 1562 2482
rect 1614 3238 1618 3242
rect 1630 3158 1634 3162
rect 1630 3138 1634 3142
rect 1662 3568 1666 3572
rect 1694 4058 1698 4062
rect 1686 3538 1690 3542
rect 1694 3538 1698 3542
rect 1662 3518 1666 3522
rect 1678 3518 1682 3522
rect 1686 3518 1690 3522
rect 1670 3158 1674 3162
rect 1694 3138 1698 3142
rect 1662 3118 1666 3122
rect 1654 3078 1658 3082
rect 1630 2978 1634 2982
rect 1646 2968 1650 2972
rect 1638 2928 1642 2932
rect 1606 2878 1610 2882
rect 1630 2858 1634 2862
rect 1590 2708 1594 2712
rect 1654 2958 1658 2962
rect 1646 2838 1650 2842
rect 1518 2328 1522 2332
rect 1550 2318 1554 2322
rect 1542 2148 1546 2152
rect 1534 2138 1538 2142
rect 1574 2458 1578 2462
rect 1582 2378 1586 2382
rect 1638 2368 1642 2372
rect 1638 2338 1642 2342
rect 1598 2318 1602 2322
rect 1606 2288 1610 2292
rect 1590 2188 1594 2192
rect 1566 2068 1570 2072
rect 1606 2048 1610 2052
rect 1646 2138 1650 2142
rect 1582 1938 1586 1942
rect 1590 1938 1594 1942
rect 1606 1938 1610 1942
rect 1582 1918 1586 1922
rect 1566 1888 1570 1892
rect 1630 1898 1634 1902
rect 1622 1878 1626 1882
rect 1574 1848 1578 1852
rect 1614 1848 1618 1852
rect 1526 1818 1530 1822
rect 1470 1518 1474 1522
rect 1510 1558 1514 1562
rect 1526 1528 1530 1532
rect 1470 1468 1474 1472
rect 1462 1388 1466 1392
rect 1422 618 1426 622
rect 1354 403 1358 407
rect 1361 403 1362 407
rect 1362 403 1365 407
rect 1510 1458 1514 1462
rect 1518 1428 1522 1432
rect 1494 1338 1498 1342
rect 1486 1248 1490 1252
rect 1478 1118 1482 1122
rect 1486 848 1490 852
rect 1526 1158 1530 1162
rect 1542 1488 1546 1492
rect 1574 1518 1578 1522
rect 1574 1468 1578 1472
rect 1606 1348 1610 1352
rect 1646 1928 1650 1932
rect 1630 1468 1634 1472
rect 1622 1148 1626 1152
rect 1638 1078 1642 1082
rect 1494 688 1498 692
rect 1454 658 1458 662
rect 1354 203 1358 207
rect 1361 203 1362 207
rect 1362 203 1365 207
rect 850 103 854 107
rect 857 103 858 107
rect 858 103 861 107
rect 1654 1248 1658 1252
rect 1718 4068 1722 4072
rect 1734 4058 1738 4062
rect 1742 3938 1746 3942
rect 1742 3888 1746 3892
rect 1742 3838 1746 3842
rect 1710 3448 1714 3452
rect 1702 3108 1706 3112
rect 1686 3028 1690 3032
rect 1678 2758 1682 2762
rect 1678 2638 1682 2642
rect 1670 2388 1674 2392
rect 1670 2358 1674 2362
rect 1670 1748 1674 1752
rect 1686 2588 1690 2592
rect 1718 3178 1722 3182
rect 1742 3288 1746 3292
rect 1726 3088 1730 3092
rect 1734 2978 1738 2982
rect 1710 2748 1714 2752
rect 1710 2718 1714 2722
rect 1726 2628 1730 2632
rect 1702 2348 1706 2352
rect 1694 2228 1698 2232
rect 1718 2218 1722 2222
rect 1726 2198 1730 2202
rect 1702 2128 1706 2132
rect 1686 2118 1690 2122
rect 1718 2118 1722 2122
rect 1726 1988 1730 1992
rect 1702 1958 1706 1962
rect 1726 1958 1730 1962
rect 1678 1648 1682 1652
rect 1670 1258 1674 1262
rect 1662 968 1666 972
rect 1670 958 1674 962
rect 1678 928 1682 932
rect 1726 1918 1730 1922
rect 1710 1488 1714 1492
rect 1702 1458 1706 1462
rect 1782 3878 1786 3882
rect 1790 3648 1794 3652
rect 1798 3588 1802 3592
rect 1790 3558 1794 3562
rect 1798 3558 1802 3562
rect 1790 3538 1794 3542
rect 1874 4703 1878 4707
rect 1881 4703 1882 4707
rect 1882 4703 1885 4707
rect 1874 4503 1878 4507
rect 1881 4503 1882 4507
rect 1882 4503 1885 4507
rect 1874 4303 1878 4307
rect 1881 4303 1882 4307
rect 1882 4303 1885 4307
rect 1878 4118 1882 4122
rect 1874 4103 1878 4107
rect 1881 4103 1882 4107
rect 1882 4103 1885 4107
rect 1822 3858 1826 3862
rect 1838 3688 1842 3692
rect 1822 3508 1826 3512
rect 1806 3498 1810 3502
rect 1822 3498 1826 3502
rect 1790 3468 1794 3472
rect 1782 3438 1786 3442
rect 1774 3338 1778 3342
rect 1790 3268 1794 3272
rect 1782 3138 1786 3142
rect 1782 2988 1786 2992
rect 1766 2978 1770 2982
rect 1758 2838 1762 2842
rect 1758 2768 1762 2772
rect 1758 2748 1762 2752
rect 1758 2578 1762 2582
rect 1782 2718 1786 2722
rect 1806 3458 1810 3462
rect 1814 2938 1818 2942
rect 1854 4038 1858 4042
rect 1902 4138 1906 4142
rect 1926 4108 1930 4112
rect 1918 4088 1922 4092
rect 1918 4058 1922 4062
rect 1874 3903 1878 3907
rect 1881 3903 1882 3907
rect 1882 3903 1885 3907
rect 1934 4068 1938 4072
rect 1942 4058 1946 4062
rect 1926 3858 1930 3862
rect 1894 3848 1898 3852
rect 1942 3788 1946 3792
rect 1910 3738 1914 3742
rect 1934 3718 1938 3722
rect 1874 3703 1878 3707
rect 1881 3703 1882 3707
rect 1882 3703 1885 3707
rect 1854 3678 1858 3682
rect 1846 3548 1850 3552
rect 1874 3503 1878 3507
rect 1881 3503 1882 3507
rect 1882 3503 1885 3507
rect 1854 3458 1858 3462
rect 1798 2898 1802 2902
rect 1806 2878 1810 2882
rect 1798 2728 1802 2732
rect 1742 2198 1746 2202
rect 1766 2088 1770 2092
rect 1758 2068 1762 2072
rect 1750 2008 1754 2012
rect 1750 1928 1754 1932
rect 1750 1888 1754 1892
rect 1782 1998 1786 2002
rect 1782 1978 1786 1982
rect 1830 2728 1834 2732
rect 1798 2358 1802 2362
rect 1790 1758 1794 1762
rect 1766 1628 1770 1632
rect 1742 1548 1746 1552
rect 1758 1488 1762 1492
rect 1750 1468 1754 1472
rect 1726 1438 1730 1442
rect 1710 1348 1714 1352
rect 1574 488 1578 492
rect 1590 378 1594 382
rect 1534 368 1538 372
rect 1710 858 1714 862
rect 1694 478 1698 482
rect 1774 1518 1778 1522
rect 1766 1338 1770 1342
rect 1790 1358 1794 1362
rect 1782 1348 1786 1352
rect 1830 2548 1834 2552
rect 1814 2258 1818 2262
rect 1814 1798 1818 1802
rect 1838 2408 1842 2412
rect 1830 2388 1834 2392
rect 1942 3378 1946 3382
rect 1902 3358 1906 3362
rect 1874 3303 1878 3307
rect 1881 3303 1882 3307
rect 1882 3303 1885 3307
rect 1874 3103 1878 3107
rect 1881 3103 1882 3107
rect 1882 3103 1885 3107
rect 1894 3068 1898 3072
rect 1854 3058 1858 3062
rect 1918 3128 1922 3132
rect 1870 3048 1874 3052
rect 1854 3008 1858 3012
rect 1874 2903 1878 2907
rect 1881 2903 1882 2907
rect 1882 2903 1885 2907
rect 1862 2718 1866 2722
rect 1874 2703 1878 2707
rect 1881 2703 1882 2707
rect 1882 2703 1885 2707
rect 1854 2658 1858 2662
rect 1874 2503 1878 2507
rect 1881 2503 1882 2507
rect 1882 2503 1885 2507
rect 1878 2468 1882 2472
rect 1918 3038 1922 3042
rect 1918 2908 1922 2912
rect 1902 2748 1906 2752
rect 1902 2558 1906 2562
rect 1902 2468 1906 2472
rect 1846 2378 1850 2382
rect 1838 2338 1842 2342
rect 1878 2338 1882 2342
rect 1830 2328 1834 2332
rect 1846 2328 1850 2332
rect 1918 2768 1922 2772
rect 1990 4448 1994 4452
rect 1998 4238 2002 4242
rect 1966 4068 1970 4072
rect 1958 2978 1962 2982
rect 1950 2958 1954 2962
rect 1958 2958 1962 2962
rect 1982 3498 1986 3502
rect 1966 2948 1970 2952
rect 1974 2948 1978 2952
rect 1934 2708 1938 2712
rect 1934 2598 1938 2602
rect 1918 2548 1922 2552
rect 1942 2548 1946 2552
rect 1942 2508 1946 2512
rect 1926 2458 1930 2462
rect 1918 2448 1922 2452
rect 1934 2448 1938 2452
rect 1966 2598 1970 2602
rect 1958 2438 1962 2442
rect 1910 2318 1914 2322
rect 1874 2303 1878 2307
rect 1881 2303 1882 2307
rect 1882 2303 1885 2307
rect 1862 2288 1866 2292
rect 1846 2058 1850 2062
rect 1830 2028 1834 2032
rect 1822 1618 1826 1622
rect 1806 1458 1810 1462
rect 1782 728 1786 732
rect 1830 1498 1834 1502
rect 1830 1408 1834 1412
rect 1854 1988 1858 1992
rect 1926 2228 1930 2232
rect 1942 2228 1946 2232
rect 1874 2103 1878 2107
rect 1881 2103 1882 2107
rect 1882 2103 1885 2107
rect 1934 2148 1938 2152
rect 1926 2078 1930 2082
rect 1878 2068 1882 2072
rect 1862 1978 1866 1982
rect 1910 1948 1914 1952
rect 1934 2058 1938 2062
rect 1934 2038 1938 2042
rect 1886 1938 1890 1942
rect 1918 1938 1922 1942
rect 1846 1758 1850 1762
rect 1958 2348 1962 2352
rect 1966 2348 1970 2352
rect 1982 2848 1986 2852
rect 2022 4448 2026 4452
rect 2046 4298 2050 4302
rect 2014 3918 2018 3922
rect 2006 3868 2010 3872
rect 1990 2758 1994 2762
rect 2070 4458 2074 4462
rect 2054 4258 2058 4262
rect 2094 4348 2098 4352
rect 2086 4258 2090 4262
rect 2038 3958 2042 3962
rect 2038 3938 2042 3942
rect 2038 3858 2042 3862
rect 2014 3638 2018 3642
rect 2022 3428 2026 3432
rect 2014 3228 2018 3232
rect 2022 3228 2026 3232
rect 2006 3158 2010 3162
rect 2006 3148 2010 3152
rect 1990 2738 1994 2742
rect 1998 2738 2002 2742
rect 1958 2298 1962 2302
rect 1894 1908 1898 1912
rect 1874 1903 1878 1907
rect 1881 1903 1882 1907
rect 1882 1903 1885 1907
rect 1918 1788 1922 1792
rect 1874 1703 1878 1707
rect 1881 1703 1882 1707
rect 1882 1703 1885 1707
rect 1862 1678 1866 1682
rect 1846 1558 1850 1562
rect 1874 1503 1878 1507
rect 1881 1503 1882 1507
rect 1882 1503 1885 1507
rect 1886 1468 1890 1472
rect 1902 1448 1906 1452
rect 1910 1448 1914 1452
rect 1894 1438 1898 1442
rect 1894 1358 1898 1362
rect 1874 1303 1878 1307
rect 1881 1303 1882 1307
rect 1882 1303 1885 1307
rect 1870 1258 1874 1262
rect 1798 558 1802 562
rect 1782 538 1786 542
rect 1790 538 1794 542
rect 1774 478 1778 482
rect 1758 338 1762 342
rect 1814 628 1818 632
rect 1874 1103 1878 1107
rect 1881 1103 1882 1107
rect 1882 1103 1885 1107
rect 1874 903 1878 907
rect 1881 903 1882 907
rect 1882 903 1885 907
rect 1950 1818 1954 1822
rect 1934 1498 1938 1502
rect 1934 1468 1938 1472
rect 1974 1948 1978 1952
rect 1934 1448 1938 1452
rect 1934 1048 1938 1052
rect 1918 988 1922 992
rect 1910 978 1914 982
rect 1874 703 1878 707
rect 1881 703 1882 707
rect 1882 703 1885 707
rect 1874 503 1878 507
rect 1881 503 1882 507
rect 1882 503 1885 507
rect 1894 478 1898 482
rect 1934 488 1938 492
rect 1958 1238 1962 1242
rect 1966 1038 1970 1042
rect 1966 948 1970 952
rect 1958 728 1962 732
rect 1958 698 1962 702
rect 2038 3238 2042 3242
rect 2030 3148 2034 3152
rect 2022 3058 2026 3062
rect 2022 2748 2026 2752
rect 2022 2458 2026 2462
rect 2014 2438 2018 2442
rect 2022 2278 2026 2282
rect 2006 2228 2010 2232
rect 1990 2018 1994 2022
rect 2022 2208 2026 2212
rect 2014 2028 2018 2032
rect 1998 1558 2002 1562
rect 1990 1528 1994 1532
rect 1990 1508 1994 1512
rect 2014 1658 2018 1662
rect 2014 1528 2018 1532
rect 2006 1448 2010 1452
rect 2078 3948 2082 3952
rect 2118 4138 2122 4142
rect 2118 4088 2122 4092
rect 2086 3758 2090 3762
rect 2086 3748 2090 3752
rect 2078 3718 2082 3722
rect 2070 3708 2074 3712
rect 2062 3638 2066 3642
rect 2062 3598 2066 3602
rect 2054 3418 2058 3422
rect 2062 3358 2066 3362
rect 2078 3338 2082 3342
rect 2062 3298 2066 3302
rect 2054 3258 2058 3262
rect 2134 3958 2138 3962
rect 2134 3928 2138 3932
rect 2142 3878 2146 3882
rect 2102 3628 2106 3632
rect 2086 3238 2090 3242
rect 2046 2838 2050 2842
rect 2126 3368 2130 3372
rect 2134 3348 2138 3352
rect 2126 3338 2130 3342
rect 2094 2808 2098 2812
rect 2118 3148 2122 3152
rect 2126 3108 2130 3112
rect 2046 2698 2050 2702
rect 2062 2688 2066 2692
rect 2054 2668 2058 2672
rect 2054 2468 2058 2472
rect 2046 2418 2050 2422
rect 2054 2398 2058 2402
rect 2054 2368 2058 2372
rect 2078 2678 2082 2682
rect 2102 2568 2106 2572
rect 2086 2558 2090 2562
rect 2086 2498 2090 2502
rect 2102 2518 2106 2522
rect 2070 2378 2074 2382
rect 2062 2308 2066 2312
rect 2054 2278 2058 2282
rect 2070 2238 2074 2242
rect 2038 2028 2042 2032
rect 2030 2018 2034 2022
rect 2038 1868 2042 1872
rect 2070 2168 2074 2172
rect 2070 2108 2074 2112
rect 2054 2048 2058 2052
rect 2094 2448 2098 2452
rect 2118 2668 2122 2672
rect 2118 2568 2122 2572
rect 2134 3028 2138 3032
rect 2174 4148 2178 4152
rect 2158 3718 2162 3722
rect 2386 4803 2390 4807
rect 2393 4803 2394 4807
rect 2394 4803 2397 4807
rect 2198 4148 2202 4152
rect 2190 3938 2194 3942
rect 2166 3618 2170 3622
rect 2190 3668 2194 3672
rect 2150 3178 2154 3182
rect 2142 2978 2146 2982
rect 2158 2878 2162 2882
rect 2150 2868 2154 2872
rect 2150 2678 2154 2682
rect 2142 2658 2146 2662
rect 2174 2948 2178 2952
rect 2150 2648 2154 2652
rect 2158 2638 2162 2642
rect 2126 2528 2130 2532
rect 2126 2468 2130 2472
rect 2102 2358 2106 2362
rect 2118 2358 2122 2362
rect 2094 2308 2098 2312
rect 2110 2208 2114 2212
rect 2086 2168 2090 2172
rect 2102 2058 2106 2062
rect 2078 1938 2082 1942
rect 2054 1898 2058 1902
rect 2062 1868 2066 1872
rect 2142 2458 2146 2462
rect 2142 2438 2146 2442
rect 2126 2258 2130 2262
rect 2118 1978 2122 1982
rect 2110 1928 2114 1932
rect 2094 1878 2098 1882
rect 2110 1878 2114 1882
rect 2078 1868 2082 1872
rect 2070 1808 2074 1812
rect 2070 1788 2074 1792
rect 2038 1778 2042 1782
rect 2030 1698 2034 1702
rect 2046 1628 2050 1632
rect 2070 1588 2074 1592
rect 2102 1748 2106 1752
rect 2038 1498 2042 1502
rect 1982 388 1986 392
rect 2070 1338 2074 1342
rect 2062 1258 2066 1262
rect 1782 148 1786 152
rect 1874 303 1878 307
rect 1881 303 1882 307
rect 1882 303 1885 307
rect 1966 268 1970 272
rect 2046 558 2050 562
rect 2102 1588 2106 1592
rect 2118 1778 2122 1782
rect 2182 2758 2186 2762
rect 2182 2698 2186 2702
rect 2182 2668 2186 2672
rect 2182 2588 2186 2592
rect 2174 2558 2178 2562
rect 2174 2488 2178 2492
rect 2158 2478 2162 2482
rect 2174 2348 2178 2352
rect 2158 2218 2162 2222
rect 2166 2068 2170 2072
rect 2158 1968 2162 1972
rect 2094 1278 2098 1282
rect 2094 1248 2098 1252
rect 2086 1158 2090 1162
rect 2118 1148 2122 1152
rect 2142 1238 2146 1242
rect 2142 1028 2146 1032
rect 2030 248 2034 252
rect 1838 148 1842 152
rect 1874 103 1878 107
rect 1881 103 1882 107
rect 1882 103 1885 107
rect 2206 3188 2210 3192
rect 2198 3088 2202 3092
rect 2198 2788 2202 2792
rect 2206 2778 2210 2782
rect 2198 2678 2202 2682
rect 2254 4138 2258 4142
rect 2222 3098 2226 3102
rect 2262 3778 2266 3782
rect 2254 3628 2258 3632
rect 2262 3568 2266 3572
rect 2246 3488 2250 3492
rect 2246 3418 2250 3422
rect 2246 3378 2250 3382
rect 2238 3358 2242 3362
rect 2238 3148 2242 3152
rect 2222 2688 2226 2692
rect 2214 2638 2218 2642
rect 2198 2598 2202 2602
rect 2206 2538 2210 2542
rect 2214 2538 2218 2542
rect 2198 2488 2202 2492
rect 2198 2428 2202 2432
rect 2190 2308 2194 2312
rect 2174 1798 2178 1802
rect 2174 1678 2178 1682
rect 2254 3318 2258 3322
rect 2270 3298 2274 3302
rect 2278 3148 2282 3152
rect 2270 3128 2274 3132
rect 2278 3008 2282 3012
rect 2270 2818 2274 2822
rect 2278 2818 2282 2822
rect 2278 2738 2282 2742
rect 2246 2608 2250 2612
rect 2246 2568 2250 2572
rect 2222 2308 2226 2312
rect 2206 2208 2210 2212
rect 2206 2188 2210 2192
rect 2270 2668 2274 2672
rect 2262 2378 2266 2382
rect 2386 4603 2390 4607
rect 2393 4603 2394 4607
rect 2394 4603 2397 4607
rect 2386 4403 2390 4407
rect 2393 4403 2394 4407
rect 2394 4403 2397 4407
rect 2386 4203 2390 4207
rect 2393 4203 2394 4207
rect 2394 4203 2397 4207
rect 2386 4003 2390 4007
rect 2393 4003 2394 4007
rect 2394 4003 2397 4007
rect 2318 3328 2322 3332
rect 2302 2968 2306 2972
rect 2310 2968 2314 2972
rect 2302 2918 2306 2922
rect 2286 2698 2290 2702
rect 2278 2318 2282 2322
rect 2254 2258 2258 2262
rect 2246 2228 2250 2232
rect 2238 2198 2242 2202
rect 2230 2158 2234 2162
rect 2230 2098 2234 2102
rect 2222 2068 2226 2072
rect 2214 1998 2218 2002
rect 2206 1828 2210 1832
rect 2166 1578 2170 1582
rect 2182 1488 2186 1492
rect 2166 1468 2170 1472
rect 2166 1188 2170 1192
rect 2166 1158 2170 1162
rect 2166 1108 2170 1112
rect 2158 548 2162 552
rect 2190 698 2194 702
rect 2230 1848 2234 1852
rect 2238 1768 2242 1772
rect 2262 2198 2266 2202
rect 2286 2228 2290 2232
rect 2278 2198 2282 2202
rect 2270 2118 2274 2122
rect 2262 1978 2266 1982
rect 2254 1958 2258 1962
rect 2262 1958 2266 1962
rect 2230 1378 2234 1382
rect 2230 1348 2234 1352
rect 2174 538 2178 542
rect 2302 2778 2306 2782
rect 2310 2658 2314 2662
rect 2302 2508 2306 2512
rect 2326 3308 2330 3312
rect 2334 2798 2338 2802
rect 2334 2658 2338 2662
rect 2334 2638 2338 2642
rect 2386 3803 2390 3807
rect 2393 3803 2394 3807
rect 2394 3803 2397 3807
rect 2390 3788 2394 3792
rect 2366 3768 2370 3772
rect 2438 4228 2442 4232
rect 2414 3678 2418 3682
rect 2386 3603 2390 3607
rect 2393 3603 2394 3607
rect 2394 3603 2397 3607
rect 2358 2988 2362 2992
rect 2366 2988 2370 2992
rect 2326 2448 2330 2452
rect 2366 2778 2370 2782
rect 2406 3408 2410 3412
rect 2386 3403 2390 3407
rect 2393 3403 2394 3407
rect 2394 3403 2397 3407
rect 2406 3378 2410 3382
rect 2406 3208 2410 3212
rect 2386 3203 2390 3207
rect 2393 3203 2394 3207
rect 2394 3203 2397 3207
rect 2406 3158 2410 3162
rect 2386 3003 2390 3007
rect 2393 3003 2394 3007
rect 2394 3003 2397 3007
rect 2414 2908 2418 2912
rect 2386 2803 2390 2807
rect 2393 2803 2394 2807
rect 2394 2803 2397 2807
rect 2386 2603 2390 2607
rect 2393 2603 2394 2607
rect 2394 2603 2397 2607
rect 2398 2558 2402 2562
rect 2366 2458 2370 2462
rect 2374 2458 2378 2462
rect 2342 2438 2346 2442
rect 2366 2388 2370 2392
rect 2358 2338 2362 2342
rect 2326 2328 2330 2332
rect 2342 2308 2346 2312
rect 2358 2278 2362 2282
rect 2350 2268 2354 2272
rect 2294 2148 2298 2152
rect 2294 2138 2298 2142
rect 2294 2048 2298 2052
rect 2270 1738 2274 1742
rect 2278 1708 2282 1712
rect 2262 1598 2266 1602
rect 2270 1438 2274 1442
rect 2294 1478 2298 1482
rect 2262 1388 2266 1392
rect 2342 2178 2346 2182
rect 2318 2008 2322 2012
rect 2334 1898 2338 1902
rect 2326 1878 2330 1882
rect 2310 1408 2314 1412
rect 2386 2403 2390 2407
rect 2393 2403 2394 2407
rect 2394 2403 2397 2407
rect 2406 2258 2410 2262
rect 2386 2203 2390 2207
rect 2393 2203 2394 2207
rect 2394 2203 2397 2207
rect 2374 2188 2378 2192
rect 2374 2128 2378 2132
rect 2374 2108 2378 2112
rect 2358 2038 2362 2042
rect 2358 1938 2362 1942
rect 2350 1648 2354 1652
rect 2278 1188 2282 1192
rect 2262 958 2266 962
rect 2294 948 2298 952
rect 2238 748 2242 752
rect 2238 548 2242 552
rect 2318 1268 2322 1272
rect 2318 868 2322 872
rect 2310 788 2314 792
rect 2318 768 2322 772
rect 2254 568 2258 572
rect 2478 4748 2482 4752
rect 2558 4368 2562 4372
rect 2518 4338 2522 4342
rect 2470 4268 2474 4272
rect 2454 4168 2458 4172
rect 2462 3868 2466 3872
rect 2446 3708 2450 3712
rect 2438 3648 2442 3652
rect 2438 3358 2442 3362
rect 2438 3278 2442 3282
rect 2446 3158 2450 3162
rect 2518 3838 2522 3842
rect 2494 3778 2498 3782
rect 2502 3508 2506 3512
rect 2502 3378 2506 3382
rect 2486 3288 2490 3292
rect 2470 3198 2474 3202
rect 2486 3078 2490 3082
rect 2486 3068 2490 3072
rect 2486 2958 2490 2962
rect 2422 2568 2426 2572
rect 2438 2548 2442 2552
rect 2446 2468 2450 2472
rect 2462 2778 2466 2782
rect 2478 2698 2482 2702
rect 2462 2448 2466 2452
rect 2438 2418 2442 2422
rect 2386 2003 2390 2007
rect 2393 2003 2394 2007
rect 2394 2003 2397 2007
rect 2386 1803 2390 1807
rect 2393 1803 2394 1807
rect 2394 1803 2397 1807
rect 2422 1828 2426 1832
rect 2406 1638 2410 1642
rect 2414 1638 2418 1642
rect 2406 1608 2410 1612
rect 2386 1603 2390 1607
rect 2393 1603 2394 1607
rect 2394 1603 2397 1607
rect 2406 1438 2410 1442
rect 2386 1403 2390 1407
rect 2393 1403 2394 1407
rect 2394 1403 2397 1407
rect 2502 2978 2506 2982
rect 2502 2808 2506 2812
rect 2494 2448 2498 2452
rect 2526 3068 2530 3072
rect 2510 2698 2514 2702
rect 2510 2608 2514 2612
rect 2518 2458 2522 2462
rect 2542 4038 2546 4042
rect 2550 3268 2554 3272
rect 2542 3198 2546 3202
rect 2542 2738 2546 2742
rect 2534 2588 2538 2592
rect 2526 2368 2530 2372
rect 2486 2278 2490 2282
rect 2470 2268 2474 2272
rect 2454 2258 2458 2262
rect 2462 2238 2466 2242
rect 2486 2178 2490 2182
rect 2478 2118 2482 2122
rect 2462 2078 2466 2082
rect 2478 1978 2482 1982
rect 2462 1878 2466 1882
rect 2454 1868 2458 1872
rect 2486 1858 2490 1862
rect 2486 1668 2490 1672
rect 2486 1648 2490 1652
rect 2430 1598 2434 1602
rect 2454 1548 2458 1552
rect 2414 1358 2418 1362
rect 2454 1468 2458 1472
rect 2386 1203 2390 1207
rect 2393 1203 2394 1207
rect 2394 1203 2397 1207
rect 2386 1003 2390 1007
rect 2393 1003 2394 1007
rect 2394 1003 2397 1007
rect 2422 1208 2426 1212
rect 2414 998 2418 1002
rect 2422 958 2426 962
rect 2414 878 2418 882
rect 2374 838 2378 842
rect 2358 658 2362 662
rect 2334 648 2338 652
rect 2386 803 2390 807
rect 2393 803 2394 807
rect 2394 803 2397 807
rect 2386 603 2390 607
rect 2393 603 2394 607
rect 2394 603 2397 607
rect 2386 403 2390 407
rect 2393 403 2394 407
rect 2394 403 2397 407
rect 2486 1258 2490 1262
rect 2478 1148 2482 1152
rect 2510 2188 2514 2192
rect 2502 1898 2506 1902
rect 2502 1878 2506 1882
rect 2542 2418 2546 2422
rect 2542 2298 2546 2302
rect 2534 2218 2538 2222
rect 2526 2168 2530 2172
rect 2526 2118 2530 2122
rect 2518 2058 2522 2062
rect 2518 1868 2522 1872
rect 2518 1848 2522 1852
rect 2510 1568 2514 1572
rect 2518 1348 2522 1352
rect 2518 1278 2522 1282
rect 2486 858 2490 862
rect 2478 848 2482 852
rect 2494 818 2498 822
rect 2478 568 2482 572
rect 2566 4218 2570 4222
rect 2566 3618 2570 3622
rect 2574 3558 2578 3562
rect 2614 4138 2618 4142
rect 2606 3618 2610 3622
rect 2590 3548 2594 3552
rect 2598 3448 2602 3452
rect 2558 3008 2562 3012
rect 2582 2978 2586 2982
rect 2574 2948 2578 2952
rect 2582 2728 2586 2732
rect 2598 3108 2602 3112
rect 2638 3388 2642 3392
rect 2622 3338 2626 3342
rect 2590 2698 2594 2702
rect 2566 2568 2570 2572
rect 2566 2548 2570 2552
rect 2558 2538 2562 2542
rect 2558 2458 2562 2462
rect 2558 2398 2562 2402
rect 2558 2228 2562 2232
rect 2550 2188 2554 2192
rect 2550 1948 2554 1952
rect 2534 1658 2538 1662
rect 2574 2238 2578 2242
rect 2574 2188 2578 2192
rect 2606 2858 2610 2862
rect 2622 3138 2626 3142
rect 2622 3098 2626 3102
rect 2614 2708 2618 2712
rect 2654 3698 2658 3702
rect 2686 4428 2690 4432
rect 2686 4008 2690 4012
rect 2678 3868 2682 3872
rect 2662 3678 2666 3682
rect 2662 3638 2666 3642
rect 2654 3198 2658 3202
rect 2654 3128 2658 3132
rect 2646 3018 2650 3022
rect 2686 3678 2690 3682
rect 2686 3638 2690 3642
rect 2678 3548 2682 3552
rect 2670 3498 2674 3502
rect 4502 5078 4506 5082
rect 4486 5068 4490 5072
rect 4582 5058 4586 5062
rect 3950 5048 3954 5052
rect 2890 4903 2894 4907
rect 2897 4903 2898 4907
rect 2898 4903 2901 4907
rect 3262 4858 3266 4862
rect 2862 4728 2866 4732
rect 2878 4728 2882 4732
rect 2890 4703 2894 4707
rect 2897 4703 2898 4707
rect 2898 4703 2901 4707
rect 2902 4668 2906 4672
rect 2870 4658 2874 4662
rect 2790 4548 2794 4552
rect 2710 3728 2714 3732
rect 2710 3698 2714 3702
rect 2742 3608 2746 3612
rect 2710 3478 2714 3482
rect 2678 3178 2682 3182
rect 2670 2958 2674 2962
rect 2670 2938 2674 2942
rect 2654 2908 2658 2912
rect 2662 2858 2666 2862
rect 2590 2168 2594 2172
rect 2566 1818 2570 1822
rect 2566 1778 2570 1782
rect 2590 1858 2594 1862
rect 2558 1508 2562 1512
rect 2550 1458 2554 1462
rect 2550 1418 2554 1422
rect 2542 1358 2546 1362
rect 2550 1338 2554 1342
rect 2534 1258 2538 1262
rect 2574 1288 2578 1292
rect 2526 478 2530 482
rect 2614 2358 2618 2362
rect 2606 2168 2610 2172
rect 2622 2158 2626 2162
rect 2598 1128 2602 1132
rect 2662 2808 2666 2812
rect 2678 2828 2682 2832
rect 2766 4128 2770 4132
rect 2782 3748 2786 3752
rect 2766 3668 2770 3672
rect 2774 3608 2778 3612
rect 2710 3318 2714 3322
rect 2734 3318 2738 3322
rect 2702 3088 2706 3092
rect 2694 2928 2698 2932
rect 2678 2808 2682 2812
rect 2702 2768 2706 2772
rect 2662 2468 2666 2472
rect 2662 2418 2666 2422
rect 2654 2378 2658 2382
rect 2670 2308 2674 2312
rect 2646 2258 2650 2262
rect 2654 2258 2658 2262
rect 2670 2108 2674 2112
rect 2630 2028 2634 2032
rect 2630 1908 2634 1912
rect 2630 1808 2634 1812
rect 2622 1618 2626 1622
rect 2622 1478 2626 1482
rect 2694 2508 2698 2512
rect 2694 2398 2698 2402
rect 2694 2378 2698 2382
rect 2686 2298 2690 2302
rect 2646 1998 2650 2002
rect 2678 1998 2682 2002
rect 2678 1948 2682 1952
rect 2662 1938 2666 1942
rect 2654 1878 2658 1882
rect 2646 1718 2650 1722
rect 2670 1848 2674 1852
rect 2662 1798 2666 1802
rect 2646 1458 2650 1462
rect 2638 1388 2642 1392
rect 2630 1088 2634 1092
rect 2678 1668 2682 1672
rect 2710 2688 2714 2692
rect 2718 2528 2722 2532
rect 2742 3268 2746 3272
rect 2734 3068 2738 3072
rect 2758 3328 2762 3332
rect 2750 2898 2754 2902
rect 2790 3398 2794 3402
rect 2782 3188 2786 3192
rect 2766 2948 2770 2952
rect 2758 2828 2762 2832
rect 2726 2518 2730 2522
rect 2726 2408 2730 2412
rect 2718 2318 2722 2322
rect 2710 2248 2714 2252
rect 2726 2248 2730 2252
rect 2710 2048 2714 2052
rect 2830 4538 2834 4542
rect 2862 4518 2866 4522
rect 2838 4298 2842 4302
rect 2830 4278 2834 4282
rect 2822 4108 2826 4112
rect 2854 4188 2858 4192
rect 2854 4038 2858 4042
rect 2950 4548 2954 4552
rect 2890 4503 2894 4507
rect 2897 4503 2898 4507
rect 2898 4503 2901 4507
rect 2890 4303 2894 4307
rect 2897 4303 2898 4307
rect 2898 4303 2901 4307
rect 2886 4278 2890 4282
rect 2890 4103 2894 4107
rect 2897 4103 2898 4107
rect 2898 4103 2901 4107
rect 2926 4148 2930 4152
rect 2918 4038 2922 4042
rect 2870 4008 2874 4012
rect 2854 3968 2858 3972
rect 2854 3928 2858 3932
rect 2806 3398 2810 3402
rect 2838 3268 2842 3272
rect 2838 3248 2842 3252
rect 2798 3198 2802 3202
rect 2790 3048 2794 3052
rect 2798 2748 2802 2752
rect 2822 3168 2826 3172
rect 2838 3148 2842 3152
rect 2806 2668 2810 2672
rect 2798 2658 2802 2662
rect 2790 2638 2794 2642
rect 2838 3108 2842 3112
rect 2830 3068 2834 3072
rect 2854 3628 2858 3632
rect 2854 3298 2858 3302
rect 2890 3903 2894 3907
rect 2897 3903 2898 3907
rect 2898 3903 2901 3907
rect 2878 3828 2882 3832
rect 2890 3703 2894 3707
rect 2897 3703 2898 3707
rect 2898 3703 2901 3707
rect 2890 3503 2894 3507
rect 2897 3503 2898 3507
rect 2898 3503 2901 3507
rect 2910 3378 2914 3382
rect 2890 3303 2894 3307
rect 2897 3303 2898 3307
rect 2898 3303 2901 3307
rect 2902 3228 2906 3232
rect 2910 3178 2914 3182
rect 2870 3158 2874 3162
rect 2854 3118 2858 3122
rect 2758 2568 2762 2572
rect 2758 2468 2762 2472
rect 2822 2548 2826 2552
rect 2774 2518 2778 2522
rect 2782 2518 2786 2522
rect 2766 2458 2770 2462
rect 2742 2428 2746 2432
rect 2742 2248 2746 2252
rect 2798 2508 2802 2512
rect 2790 2498 2794 2502
rect 2782 2458 2786 2462
rect 2790 2368 2794 2372
rect 2814 2368 2818 2372
rect 2838 2408 2842 2412
rect 2806 2338 2810 2342
rect 2742 2208 2746 2212
rect 2734 2018 2738 2022
rect 2758 2118 2762 2122
rect 2742 1958 2746 1962
rect 2694 1628 2698 1632
rect 2710 1778 2714 1782
rect 2710 1658 2714 1662
rect 2702 1218 2706 1222
rect 2686 1168 2690 1172
rect 2670 1068 2674 1072
rect 2726 1168 2730 1172
rect 2726 1068 2730 1072
rect 2702 1018 2706 1022
rect 2710 968 2714 972
rect 2710 948 2714 952
rect 2326 248 2330 252
rect 2386 203 2390 207
rect 2393 203 2394 207
rect 2394 203 2397 207
rect 2750 1858 2754 1862
rect 2750 1768 2754 1772
rect 2774 1958 2778 1962
rect 2766 1928 2770 1932
rect 2766 1918 2770 1922
rect 2758 1688 2762 1692
rect 2774 1318 2778 1322
rect 2846 2278 2850 2282
rect 2822 2248 2826 2252
rect 2838 2198 2842 2202
rect 2806 2078 2810 2082
rect 2806 2068 2810 2072
rect 2806 1978 2810 1982
rect 2798 1968 2802 1972
rect 2798 1588 2802 1592
rect 2798 1348 2802 1352
rect 2790 988 2794 992
rect 2822 1888 2826 1892
rect 2822 1858 2826 1862
rect 2782 938 2786 942
rect 2890 3103 2894 3107
rect 2897 3103 2898 3107
rect 2898 3103 2901 3107
rect 2878 3068 2882 3072
rect 2934 3778 2938 3782
rect 3070 4748 3074 4752
rect 2950 4248 2954 4252
rect 2958 4238 2962 4242
rect 2926 3728 2930 3732
rect 2910 2968 2914 2972
rect 2890 2903 2894 2907
rect 2897 2903 2898 2907
rect 2898 2903 2901 2907
rect 2910 2888 2914 2892
rect 2870 2828 2874 2832
rect 2910 2828 2914 2832
rect 2862 2448 2866 2452
rect 2862 2358 2866 2362
rect 2890 2703 2894 2707
rect 2897 2703 2898 2707
rect 2898 2703 2901 2707
rect 2878 2678 2882 2682
rect 2902 2558 2906 2562
rect 2886 2528 2890 2532
rect 2890 2503 2894 2507
rect 2897 2503 2898 2507
rect 2898 2503 2901 2507
rect 2878 2478 2882 2482
rect 2894 2428 2898 2432
rect 2886 2338 2890 2342
rect 2890 2303 2894 2307
rect 2897 2303 2898 2307
rect 2898 2303 2901 2307
rect 2934 3668 2938 3672
rect 2942 3358 2946 3362
rect 2942 3188 2946 3192
rect 2934 3098 2938 3102
rect 2934 3048 2938 3052
rect 2918 2488 2922 2492
rect 2918 2268 2922 2272
rect 2846 1958 2850 1962
rect 2862 1848 2866 1852
rect 2870 1838 2874 1842
rect 2838 1518 2842 1522
rect 2870 1728 2874 1732
rect 2910 2118 2914 2122
rect 2890 2103 2894 2107
rect 2897 2103 2898 2107
rect 2898 2103 2901 2107
rect 2942 2858 2946 2862
rect 3038 4148 3042 4152
rect 3030 4138 3034 4142
rect 2990 3718 2994 3722
rect 2966 3688 2970 3692
rect 2990 3698 2994 3702
rect 2982 3648 2986 3652
rect 2966 3528 2970 3532
rect 2982 3378 2986 3382
rect 2958 2778 2962 2782
rect 2958 2738 2962 2742
rect 2990 3088 2994 3092
rect 2990 2938 2994 2942
rect 3014 4058 3018 4062
rect 3054 4028 3058 4032
rect 3054 4018 3058 4022
rect 3046 3758 3050 3762
rect 3046 3678 3050 3682
rect 3030 3668 3034 3672
rect 3038 3658 3042 3662
rect 3030 3578 3034 3582
rect 3014 3418 3018 3422
rect 3014 3318 3018 3322
rect 3006 2918 3010 2922
rect 2998 2868 3002 2872
rect 3006 2868 3010 2872
rect 2990 2838 2994 2842
rect 2958 2648 2962 2652
rect 2950 2548 2954 2552
rect 2934 2458 2938 2462
rect 2990 2638 2994 2642
rect 2990 2568 2994 2572
rect 2982 2558 2986 2562
rect 2982 2488 2986 2492
rect 2974 2458 2978 2462
rect 2966 2398 2970 2402
rect 2950 2348 2954 2352
rect 2974 2388 2978 2392
rect 2926 2098 2930 2102
rect 2890 1903 2894 1907
rect 2897 1903 2898 1907
rect 2898 1903 2901 1907
rect 2918 1838 2922 1842
rect 2890 1703 2894 1707
rect 2897 1703 2898 1707
rect 2898 1703 2901 1707
rect 2918 1688 2922 1692
rect 2918 1608 2922 1612
rect 2958 2078 2962 2082
rect 2990 2298 2994 2302
rect 3038 3408 3042 3412
rect 3070 3838 3074 3842
rect 3038 3348 3042 3352
rect 3030 3158 3034 3162
rect 3046 3148 3050 3152
rect 3054 3028 3058 3032
rect 3062 3028 3066 3032
rect 3030 2978 3034 2982
rect 3046 2968 3050 2972
rect 3038 2948 3042 2952
rect 3030 2928 3034 2932
rect 3118 4458 3122 4462
rect 3126 4358 3130 4362
rect 3086 4008 3090 4012
rect 3078 3728 3082 3732
rect 3102 3538 3106 3542
rect 3102 3508 3106 3512
rect 3094 3328 3098 3332
rect 3086 3058 3090 3062
rect 3062 2818 3066 2822
rect 3054 2728 3058 2732
rect 3022 2638 3026 2642
rect 3006 2548 3010 2552
rect 3030 2548 3034 2552
rect 3006 2508 3010 2512
rect 3022 2508 3026 2512
rect 3014 2498 3018 2502
rect 3030 2488 3034 2492
rect 3006 2428 3010 2432
rect 2990 2278 2994 2282
rect 2998 2278 3002 2282
rect 3030 2348 3034 2352
rect 3022 2328 3026 2332
rect 3030 2278 3034 2282
rect 3006 2108 3010 2112
rect 2982 2068 2986 2072
rect 2958 1958 2962 1962
rect 2934 1748 2938 1752
rect 2918 1588 2922 1592
rect 2890 1503 2894 1507
rect 2897 1503 2898 1507
rect 2898 1503 2901 1507
rect 2910 1458 2914 1462
rect 2854 1338 2858 1342
rect 2846 1178 2850 1182
rect 2890 1303 2894 1307
rect 2897 1303 2898 1307
rect 2898 1303 2901 1307
rect 2950 1748 2954 1752
rect 2958 1648 2962 1652
rect 2958 1298 2962 1302
rect 2958 1258 2962 1262
rect 2890 1103 2894 1107
rect 2897 1103 2898 1107
rect 2898 1103 2901 1107
rect 2878 988 2882 992
rect 2890 903 2894 907
rect 2897 903 2898 907
rect 2898 903 2901 907
rect 2890 703 2894 707
rect 2897 703 2898 707
rect 2898 703 2901 707
rect 2942 1108 2946 1112
rect 2918 1058 2922 1062
rect 2942 1048 2946 1052
rect 2926 898 2930 902
rect 3022 2048 3026 2052
rect 3070 2808 3074 2812
rect 3086 2608 3090 2612
rect 3174 4268 3178 4272
rect 3150 3748 3154 3752
rect 3126 3568 3130 3572
rect 3110 3438 3114 3442
rect 3110 3398 3114 3402
rect 3102 3178 3106 3182
rect 3150 3578 3154 3582
rect 3150 3468 3154 3472
rect 3142 3438 3146 3442
rect 3182 3978 3186 3982
rect 3174 3888 3178 3892
rect 3206 4348 3210 4352
rect 3206 4288 3210 4292
rect 3206 4008 3210 4012
rect 3206 3828 3210 3832
rect 3206 3758 3210 3762
rect 3214 3758 3218 3762
rect 3174 3648 3178 3652
rect 3214 3648 3218 3652
rect 3174 3468 3178 3472
rect 3142 3208 3146 3212
rect 3110 2798 3114 2802
rect 3102 2628 3106 2632
rect 3094 2598 3098 2602
rect 3046 2468 3050 2472
rect 3046 2368 3050 2372
rect 3038 2038 3042 2042
rect 3030 1808 3034 1812
rect 3022 1738 3026 1742
rect 2998 1648 3002 1652
rect 3022 1518 3026 1522
rect 2998 1448 3002 1452
rect 3006 1388 3010 1392
rect 3006 1368 3010 1372
rect 2982 1338 2986 1342
rect 3006 1318 3010 1322
rect 2990 1258 2994 1262
rect 3022 1338 3026 1342
rect 3014 1168 3018 1172
rect 3038 1228 3042 1232
rect 3030 1158 3034 1162
rect 3038 1158 3042 1162
rect 3014 1138 3018 1142
rect 3030 1128 3034 1132
rect 2886 558 2890 562
rect 2890 503 2894 507
rect 2897 503 2898 507
rect 2898 503 2901 507
rect 2702 448 2706 452
rect 2782 468 2786 472
rect 2870 458 2874 462
rect 2890 303 2894 307
rect 2897 303 2898 307
rect 2898 303 2901 307
rect 2974 728 2978 732
rect 2990 1068 2994 1072
rect 2990 868 2994 872
rect 2990 848 2994 852
rect 3030 888 3034 892
rect 3070 2588 3074 2592
rect 3062 2578 3066 2582
rect 3078 2558 3082 2562
rect 3086 2538 3090 2542
rect 3102 2548 3106 2552
rect 3062 2408 3066 2412
rect 3102 2398 3106 2402
rect 3078 2388 3082 2392
rect 3062 2358 3066 2362
rect 3078 2108 3082 2112
rect 3078 1978 3082 1982
rect 3142 2978 3146 2982
rect 3142 2698 3146 2702
rect 3110 2338 3114 2342
rect 3134 2508 3138 2512
rect 3150 2438 3154 2442
rect 3150 2428 3154 2432
rect 3134 2318 3138 2322
rect 3134 2258 3138 2262
rect 3150 1868 3154 1872
rect 3110 1818 3114 1822
rect 3070 1598 3074 1602
rect 3062 1418 3066 1422
rect 3094 1568 3098 1572
rect 3086 1528 3090 1532
rect 3022 768 3026 772
rect 3030 758 3034 762
rect 3006 448 3010 452
rect 3054 818 3058 822
rect 3110 1658 3114 1662
rect 3150 1688 3154 1692
rect 3142 1668 3146 1672
rect 3150 1668 3154 1672
rect 3118 1558 3122 1562
rect 3110 1538 3114 1542
rect 3142 1528 3146 1532
rect 3102 1448 3106 1452
rect 3118 1448 3122 1452
rect 3062 648 3066 652
rect 3038 628 3042 632
rect 3110 1148 3114 1152
rect 3126 1278 3130 1282
rect 3134 1268 3138 1272
rect 3206 3538 3210 3542
rect 3254 4438 3258 4442
rect 3222 3588 3226 3592
rect 3198 3528 3202 3532
rect 3206 3478 3210 3482
rect 3206 3448 3210 3452
rect 3198 3168 3202 3172
rect 3182 3118 3186 3122
rect 3174 2968 3178 2972
rect 3206 2988 3210 2992
rect 3166 2748 3170 2752
rect 3190 2838 3194 2842
rect 3174 2518 3178 2522
rect 3166 2348 3170 2352
rect 3182 2468 3186 2472
rect 3402 5003 3406 5007
rect 3409 5003 3410 5007
rect 3410 5003 3413 5007
rect 3402 4803 3406 4807
rect 3409 4803 3410 4807
rect 3410 4803 3413 4807
rect 3366 4668 3370 4672
rect 3402 4603 3406 4607
rect 3409 4603 3410 4607
rect 3410 4603 3413 4607
rect 3402 4403 3406 4407
rect 3409 4403 3410 4407
rect 3410 4403 3413 4407
rect 3342 4348 3346 4352
rect 3398 4348 3402 4352
rect 3334 4328 3338 4332
rect 3294 3858 3298 3862
rect 3270 3848 3274 3852
rect 3262 3738 3266 3742
rect 3254 3628 3258 3632
rect 3238 3498 3242 3502
rect 3230 3428 3234 3432
rect 3230 3398 3234 3402
rect 3294 3628 3298 3632
rect 3262 3308 3266 3312
rect 3262 3068 3266 3072
rect 3254 2958 3258 2962
rect 3246 2848 3250 2852
rect 3222 2728 3226 2732
rect 3238 2618 3242 2622
rect 3198 2488 3202 2492
rect 3246 2608 3250 2612
rect 3238 2478 3242 2482
rect 3222 2458 3226 2462
rect 3166 1788 3170 1792
rect 3150 1078 3154 1082
rect 3142 918 3146 922
rect 3166 1288 3170 1292
rect 3166 1168 3170 1172
rect 3190 2398 3194 2402
rect 3222 2358 3226 2362
rect 3198 2338 3202 2342
rect 3238 2448 3242 2452
rect 3214 2288 3218 2292
rect 3222 2288 3226 2292
rect 3230 2258 3234 2262
rect 3206 2248 3210 2252
rect 3206 1978 3210 1982
rect 3198 1928 3202 1932
rect 3182 1878 3186 1882
rect 3190 1828 3194 1832
rect 3174 948 3178 952
rect 3198 1728 3202 1732
rect 3158 528 3162 532
rect 3054 388 3058 392
rect 3230 1688 3234 1692
rect 3222 1658 3226 1662
rect 3222 1278 3226 1282
rect 3238 1678 3242 1682
rect 3310 3678 3314 3682
rect 3310 3568 3314 3572
rect 3382 3988 3386 3992
rect 3402 4203 3406 4207
rect 3409 4203 3410 4207
rect 3410 4203 3413 4207
rect 3402 4003 3406 4007
rect 3409 4003 3410 4007
rect 3410 4003 3413 4007
rect 3398 3918 3402 3922
rect 3382 3818 3386 3822
rect 3374 3748 3378 3752
rect 3342 3728 3346 3732
rect 3302 3278 3306 3282
rect 3302 3268 3306 3272
rect 3302 3008 3306 3012
rect 3286 2748 3290 2752
rect 3334 3038 3338 3042
rect 3326 2758 3330 2762
rect 3318 2648 3322 2652
rect 3302 2618 3306 2622
rect 3294 2528 3298 2532
rect 3278 2488 3282 2492
rect 3278 2208 3282 2212
rect 3286 2148 3290 2152
rect 3286 2048 3290 2052
rect 3286 2038 3290 2042
rect 3278 1988 3282 1992
rect 3270 1948 3274 1952
rect 3270 1938 3274 1942
rect 3278 1578 3282 1582
rect 3262 1538 3266 1542
rect 3254 1448 3258 1452
rect 3334 2528 3338 2532
rect 3310 2508 3314 2512
rect 3326 2508 3330 2512
rect 3358 3708 3362 3712
rect 3350 3678 3354 3682
rect 3366 3658 3370 3662
rect 3366 3478 3370 3482
rect 3350 3268 3354 3272
rect 3382 3368 3386 3372
rect 3402 3803 3406 3807
rect 3409 3803 3410 3807
rect 3410 3803 3413 3807
rect 3438 4838 3442 4842
rect 3462 4528 3466 4532
rect 3454 4448 3458 4452
rect 3430 3878 3434 3882
rect 3402 3603 3406 3607
rect 3409 3603 3410 3607
rect 3410 3603 3413 3607
rect 3446 3608 3450 3612
rect 3438 3548 3442 3552
rect 3446 3528 3450 3532
rect 3402 3403 3406 3407
rect 3409 3403 3410 3407
rect 3410 3403 3413 3407
rect 3402 3203 3406 3207
rect 3409 3203 3410 3207
rect 3410 3203 3413 3207
rect 3374 3198 3378 3202
rect 3358 2708 3362 2712
rect 3350 2518 3354 2522
rect 3326 2468 3330 2472
rect 3342 2468 3346 2472
rect 3342 2438 3346 2442
rect 3334 2408 3338 2412
rect 3318 2368 3322 2372
rect 3334 2368 3338 2372
rect 3342 2338 3346 2342
rect 3326 2328 3330 2332
rect 3302 2198 3306 2202
rect 3326 2198 3330 2202
rect 3302 2188 3306 2192
rect 3310 2038 3314 2042
rect 3342 2188 3346 2192
rect 3334 2138 3338 2142
rect 3302 1908 3306 1912
rect 3286 1438 3290 1442
rect 3302 1768 3306 1772
rect 3302 1458 3306 1462
rect 3294 1338 3298 1342
rect 3278 1278 3282 1282
rect 3270 1148 3274 1152
rect 3230 1088 3234 1092
rect 3222 1048 3226 1052
rect 3222 958 3226 962
rect 3294 1098 3298 1102
rect 3334 1558 3338 1562
rect 3318 1208 3322 1212
rect 3310 1158 3314 1162
rect 3382 3018 3386 3022
rect 3402 3003 3406 3007
rect 3409 3003 3410 3007
rect 3410 3003 3413 3007
rect 3390 2938 3394 2942
rect 3446 3338 3450 3342
rect 3534 4548 3538 4552
rect 3526 4458 3530 4462
rect 3486 4218 3490 4222
rect 3526 4258 3530 4262
rect 3550 4258 3554 4262
rect 3510 4058 3514 4062
rect 3486 3948 3490 3952
rect 3486 3668 3490 3672
rect 3470 3508 3474 3512
rect 3518 3888 3522 3892
rect 3462 3218 3466 3222
rect 3454 3158 3458 3162
rect 3430 3028 3434 3032
rect 3422 2918 3426 2922
rect 3402 2803 3406 2807
rect 3409 2803 3410 2807
rect 3410 2803 3413 2807
rect 3402 2603 3406 2607
rect 3409 2603 3410 2607
rect 3410 2603 3413 2607
rect 3406 2558 3410 2562
rect 3390 2518 3394 2522
rect 3402 2403 3406 2407
rect 3409 2403 3410 2407
rect 3410 2403 3413 2407
rect 3414 2338 3418 2342
rect 3398 2328 3402 2332
rect 3406 2318 3410 2322
rect 3390 2308 3394 2312
rect 3382 2258 3386 2262
rect 3374 2238 3378 2242
rect 3402 2203 3406 2207
rect 3409 2203 3410 2207
rect 3410 2203 3413 2207
rect 3366 2148 3370 2152
rect 3462 2918 3466 2922
rect 3462 2818 3466 2822
rect 3462 2718 3466 2722
rect 3454 2638 3458 2642
rect 3446 2378 3450 2382
rect 3446 2358 3450 2362
rect 3438 2288 3442 2292
rect 3454 2228 3458 2232
rect 3414 2068 3418 2072
rect 3350 1878 3354 1882
rect 3342 1548 3346 1552
rect 3382 1798 3386 1802
rect 3402 2003 3406 2007
rect 3409 2003 3410 2007
rect 3410 2003 3413 2007
rect 3430 1968 3434 1972
rect 3414 1958 3418 1962
rect 3402 1803 3406 1807
rect 3409 1803 3410 1807
rect 3410 1803 3413 1807
rect 3398 1658 3402 1662
rect 3402 1603 3406 1607
rect 3409 1603 3410 1607
rect 3410 1603 3413 1607
rect 3430 1548 3434 1552
rect 3402 1403 3406 1407
rect 3409 1403 3410 1407
rect 3410 1403 3413 1407
rect 3350 1368 3354 1372
rect 3582 4828 3586 4832
rect 3598 4238 3602 4242
rect 3526 3848 3530 3852
rect 3534 3738 3538 3742
rect 3542 3698 3546 3702
rect 3518 3318 3522 3322
rect 3558 3618 3562 3622
rect 3494 2748 3498 2752
rect 3502 2688 3506 2692
rect 3494 2678 3498 2682
rect 3486 2668 3490 2672
rect 3470 2468 3474 2472
rect 3470 2298 3474 2302
rect 3470 2258 3474 2262
rect 3438 1428 3442 1432
rect 3334 1138 3338 1142
rect 3294 728 3298 732
rect 3318 658 3322 662
rect 3390 1208 3394 1212
rect 3358 1198 3362 1202
rect 3358 1138 3362 1142
rect 3358 1118 3362 1122
rect 3358 868 3362 872
rect 3402 1203 3406 1207
rect 3409 1203 3410 1207
rect 3410 1203 3413 1207
rect 3402 1003 3406 1007
rect 3409 1003 3410 1007
rect 3410 1003 3413 1007
rect 3454 1608 3458 1612
rect 3454 1588 3458 1592
rect 3486 2408 3490 2412
rect 3486 2338 3490 2342
rect 3486 2328 3490 2332
rect 3518 2448 3522 2452
rect 3510 2368 3514 2372
rect 3502 2348 3506 2352
rect 3518 2318 3522 2322
rect 3542 2828 3546 2832
rect 3542 2658 3546 2662
rect 3534 2608 3538 2612
rect 3566 3558 3570 3562
rect 3574 3498 3578 3502
rect 3566 3488 3570 3492
rect 3574 3488 3578 3492
rect 3574 3348 3578 3352
rect 3558 2968 3562 2972
rect 3566 2828 3570 2832
rect 3558 2768 3562 2772
rect 3558 2588 3562 2592
rect 3534 2278 3538 2282
rect 3518 2268 3522 2272
rect 3518 2068 3522 2072
rect 3502 1948 3506 1952
rect 3494 1858 3498 1862
rect 3470 1538 3474 1542
rect 3462 1388 3466 1392
rect 3494 1468 3498 1472
rect 3502 1388 3506 1392
rect 3526 1308 3530 1312
rect 3526 1198 3530 1202
rect 3414 868 3418 872
rect 3402 803 3406 807
rect 3409 803 3410 807
rect 3410 803 3413 807
rect 3494 758 3498 762
rect 3454 688 3458 692
rect 3402 603 3406 607
rect 3409 603 3410 607
rect 3410 603 3413 607
rect 3470 448 3474 452
rect 3402 403 3406 407
rect 3409 403 3410 407
rect 3410 403 3413 407
rect 3278 358 3282 362
rect 3198 348 3202 352
rect 2990 148 2994 152
rect 3078 148 3082 152
rect 3102 148 3106 152
rect 2890 103 2894 107
rect 2897 103 2898 107
rect 2898 103 2901 107
rect 2542 78 2546 82
rect 2822 68 2826 72
rect 3402 203 3406 207
rect 3409 203 3410 207
rect 3410 203 3413 207
rect 3094 78 3098 82
rect 3486 268 3490 272
rect 3470 98 3474 102
rect 3486 88 3490 92
rect 3558 2328 3562 2332
rect 3550 2288 3554 2292
rect 3550 2258 3554 2262
rect 3590 3768 3594 3772
rect 3638 4428 3642 4432
rect 3638 3978 3642 3982
rect 3598 3748 3602 3752
rect 3598 3678 3602 3682
rect 3590 2718 3594 2722
rect 3574 2478 3578 2482
rect 3582 2388 3586 2392
rect 3606 3328 3610 3332
rect 3646 3468 3650 3472
rect 3662 3688 3666 3692
rect 3654 3228 3658 3232
rect 3630 3058 3634 3062
rect 3606 2678 3610 2682
rect 3606 2648 3610 2652
rect 3598 2478 3602 2482
rect 3558 2068 3562 2072
rect 3542 1948 3546 1952
rect 3542 1888 3546 1892
rect 3542 1868 3546 1872
rect 3550 1828 3554 1832
rect 3542 1748 3546 1752
rect 3542 1578 3546 1582
rect 3566 1738 3570 1742
rect 3558 1218 3562 1222
rect 3614 2458 3618 2462
rect 3614 2388 3618 2392
rect 3614 2288 3618 2292
rect 3606 2168 3610 2172
rect 3598 2068 3602 2072
rect 3598 2048 3602 2052
rect 3614 2068 3618 2072
rect 3662 3068 3666 3072
rect 3638 2688 3642 2692
rect 3686 3938 3690 3942
rect 3922 4903 3926 4907
rect 3929 4903 3930 4907
rect 3930 4903 3933 4907
rect 3922 4703 3926 4707
rect 3929 4703 3930 4707
rect 3930 4703 3933 4707
rect 3942 4558 3946 4562
rect 3870 4538 3874 4542
rect 3838 4438 3842 4442
rect 3726 3948 3730 3952
rect 3678 3528 3682 3532
rect 3718 3858 3722 3862
rect 3702 3578 3706 3582
rect 3702 3568 3706 3572
rect 3678 3088 3682 3092
rect 3734 3678 3738 3682
rect 3726 3588 3730 3592
rect 3726 3378 3730 3382
rect 3718 3368 3722 3372
rect 3710 3268 3714 3272
rect 3646 2658 3650 2662
rect 3654 2658 3658 2662
rect 3646 2568 3650 2572
rect 3630 2498 3634 2502
rect 3638 2348 3642 2352
rect 3638 2268 3642 2272
rect 3790 3968 3794 3972
rect 3774 3958 3778 3962
rect 3766 3868 3770 3872
rect 3750 3538 3754 3542
rect 3742 3048 3746 3052
rect 3734 2818 3738 2822
rect 3726 2688 3730 2692
rect 3734 2638 3738 2642
rect 3678 2328 3682 2332
rect 3678 2248 3682 2252
rect 3574 1588 3578 1592
rect 3590 1618 3594 1622
rect 3614 1458 3618 1462
rect 3606 1368 3610 1372
rect 3582 1258 3586 1262
rect 3574 1198 3578 1202
rect 3686 2078 3690 2082
rect 3686 2028 3690 2032
rect 3630 1868 3634 1872
rect 3662 1868 3666 1872
rect 3670 1798 3674 1802
rect 3654 1778 3658 1782
rect 3654 1738 3658 1742
rect 3622 1138 3626 1142
rect 3526 838 3530 842
rect 3542 648 3546 652
rect 3542 468 3546 472
rect 3534 448 3538 452
rect 3542 348 3546 352
rect 3534 268 3538 272
rect 3430 68 3434 72
rect 3622 668 3626 672
rect 3662 1558 3666 1562
rect 3654 1458 3658 1462
rect 3638 1108 3642 1112
rect 3654 868 3658 872
rect 3638 808 3642 812
rect 3638 528 3642 532
rect 3670 1358 3674 1362
rect 3734 2468 3738 2472
rect 3734 2418 3738 2422
rect 3734 2358 3738 2362
rect 3726 2178 3730 2182
rect 3734 2138 3738 2142
rect 3718 2058 3722 2062
rect 3710 1938 3714 1942
rect 3710 1848 3714 1852
rect 3798 3848 3802 3852
rect 3814 3848 3818 3852
rect 3806 3518 3810 3522
rect 3830 3558 3834 3562
rect 3822 3488 3826 3492
rect 3822 3308 3826 3312
rect 3814 3258 3818 3262
rect 3798 2778 3802 2782
rect 3806 2708 3810 2712
rect 3790 2668 3794 2672
rect 3798 2668 3802 2672
rect 3774 2558 3778 2562
rect 3798 2548 3802 2552
rect 3766 2368 3770 2372
rect 3798 2368 3802 2372
rect 3750 1918 3754 1922
rect 3702 1538 3706 1542
rect 3734 1468 3738 1472
rect 3702 1358 3706 1362
rect 3694 1158 3698 1162
rect 3686 1048 3690 1052
rect 3678 908 3682 912
rect 3726 1168 3730 1172
rect 3742 1438 3746 1442
rect 3774 1878 3778 1882
rect 3790 1758 3794 1762
rect 3766 1638 3770 1642
rect 3742 1228 3746 1232
rect 3742 1098 3746 1102
rect 3726 858 3730 862
rect 3718 838 3722 842
rect 3838 3238 3842 3242
rect 3830 2658 3834 2662
rect 3814 2508 3818 2512
rect 3846 3158 3850 3162
rect 3922 4503 3926 4507
rect 3929 4503 3930 4507
rect 3930 4503 3933 4507
rect 3934 4368 3938 4372
rect 3886 4338 3890 4342
rect 3922 4303 3926 4307
rect 3929 4303 3930 4307
rect 3930 4303 3933 4307
rect 3910 4108 3914 4112
rect 3922 4103 3926 4107
rect 3929 4103 3930 4107
rect 3930 4103 3933 4107
rect 3886 4078 3890 4082
rect 3894 4038 3898 4042
rect 3894 3978 3898 3982
rect 3910 3948 3914 3952
rect 3922 3903 3926 3907
rect 3929 3903 3930 3907
rect 3930 3903 3933 3907
rect 3878 3848 3882 3852
rect 3902 3708 3906 3712
rect 3922 3703 3926 3707
rect 3929 3703 3930 3707
rect 3930 3703 3933 3707
rect 3894 3668 3898 3672
rect 3922 3503 3926 3507
rect 3929 3503 3930 3507
rect 3930 3503 3933 3507
rect 3922 3303 3926 3307
rect 3929 3303 3930 3307
rect 3930 3303 3933 3307
rect 3942 3188 3946 3192
rect 3922 3103 3926 3107
rect 3929 3103 3930 3107
rect 3930 3103 3933 3107
rect 3910 3098 3914 3102
rect 3838 2438 3842 2442
rect 3822 2268 3826 2272
rect 3862 2238 3866 2242
rect 3806 2058 3810 2062
rect 3806 1548 3810 1552
rect 3798 1428 3802 1432
rect 3790 1368 3794 1372
rect 3782 1298 3786 1302
rect 3798 1288 3802 1292
rect 3790 1258 3794 1262
rect 3782 1178 3786 1182
rect 3774 1158 3778 1162
rect 3766 1148 3770 1152
rect 3782 1078 3786 1082
rect 3750 968 3754 972
rect 3662 448 3666 452
rect 3662 368 3666 372
rect 3606 148 3610 152
rect 3638 98 3642 102
rect 3814 1298 3818 1302
rect 3846 2098 3850 2102
rect 3894 2928 3898 2932
rect 3922 2903 3926 2907
rect 3929 2903 3930 2907
rect 3930 2903 3933 2907
rect 3922 2703 3926 2707
rect 3929 2703 3930 2707
rect 3930 2703 3933 2707
rect 3902 2578 3906 2582
rect 3922 2503 3926 2507
rect 3929 2503 3930 2507
rect 3930 2503 3933 2507
rect 4426 5003 4430 5007
rect 4433 5003 4434 5007
rect 4434 5003 4437 5007
rect 4134 4848 4138 4852
rect 4134 4828 4138 4832
rect 3958 4548 3962 4552
rect 3966 4538 3970 4542
rect 3958 3128 3962 3132
rect 3950 2488 3954 2492
rect 3902 2448 3906 2452
rect 3990 3758 3994 3762
rect 4006 3738 4010 3742
rect 3998 3718 4002 3722
rect 3982 3648 3986 3652
rect 3990 3608 3994 3612
rect 3982 3298 3986 3302
rect 3974 3218 3978 3222
rect 3966 2858 3970 2862
rect 3958 2368 3962 2372
rect 3922 2303 3926 2307
rect 3929 2303 3930 2307
rect 3930 2303 3933 2307
rect 4038 4118 4042 4122
rect 4062 4328 4066 4332
rect 4062 4298 4066 4302
rect 4078 4548 4082 4552
rect 4102 4528 4106 4532
rect 4102 4438 4106 4442
rect 4070 4018 4074 4022
rect 4030 3608 4034 3612
rect 4030 3478 4034 3482
rect 4014 3438 4018 3442
rect 4022 3438 4026 3442
rect 4006 2498 4010 2502
rect 4006 2368 4010 2372
rect 3910 2268 3914 2272
rect 3894 2148 3898 2152
rect 3862 1918 3866 1922
rect 3830 1528 3834 1532
rect 3830 1318 3834 1322
rect 3830 1048 3834 1052
rect 3830 1028 3834 1032
rect 3822 898 3826 902
rect 3822 848 3826 852
rect 3846 1518 3850 1522
rect 3854 1488 3858 1492
rect 3870 1268 3874 1272
rect 3922 2103 3926 2107
rect 3929 2103 3930 2107
rect 3930 2103 3933 2107
rect 3886 2048 3890 2052
rect 3922 1903 3926 1907
rect 3929 1903 3930 1907
rect 3930 1903 3933 1907
rect 3942 1888 3946 1892
rect 3910 1858 3914 1862
rect 3950 1808 3954 1812
rect 3922 1703 3926 1707
rect 3929 1703 3930 1707
rect 3930 1703 3933 1707
rect 3910 1688 3914 1692
rect 3902 1578 3906 1582
rect 3902 1558 3906 1562
rect 3894 1548 3898 1552
rect 3922 1503 3926 1507
rect 3929 1503 3930 1507
rect 3930 1503 3933 1507
rect 3886 1258 3890 1262
rect 3878 1068 3882 1072
rect 3862 858 3866 862
rect 3950 1328 3954 1332
rect 3922 1303 3926 1307
rect 3929 1303 3930 1307
rect 3930 1303 3933 1307
rect 3910 1288 3914 1292
rect 3934 1138 3938 1142
rect 3922 1103 3926 1107
rect 3929 1103 3930 1107
rect 3930 1103 3933 1107
rect 3910 908 3914 912
rect 3922 903 3926 907
rect 3929 903 3930 907
rect 3930 903 3933 907
rect 3854 758 3858 762
rect 3922 703 3926 707
rect 3929 703 3930 707
rect 3930 703 3933 707
rect 3982 1858 3986 1862
rect 3974 1748 3978 1752
rect 3974 1448 3978 1452
rect 3998 1668 4002 1672
rect 3998 1558 4002 1562
rect 3990 1378 3994 1382
rect 3982 1318 3986 1322
rect 4022 3268 4026 3272
rect 4030 3088 4034 3092
rect 4070 3878 4074 3882
rect 4078 3878 4082 3882
rect 4062 3538 4066 3542
rect 4070 3538 4074 3542
rect 4062 3298 4066 3302
rect 4046 2908 4050 2912
rect 4054 2628 4058 2632
rect 4054 2588 4058 2592
rect 4046 2478 4050 2482
rect 4038 2468 4042 2472
rect 4014 1378 4018 1382
rect 4006 968 4010 972
rect 3998 858 4002 862
rect 3838 558 3842 562
rect 3830 458 3834 462
rect 3838 358 3842 362
rect 3750 258 3754 262
rect 3922 503 3926 507
rect 3929 503 3930 507
rect 3930 503 3933 507
rect 4038 2238 4042 2242
rect 4038 2128 4042 2132
rect 4142 4568 4146 4572
rect 4142 4538 4146 4542
rect 4174 4558 4178 4562
rect 4150 4368 4154 4372
rect 4142 4078 4146 4082
rect 4102 3358 4106 3362
rect 4102 3348 4106 3352
rect 4086 3278 4090 3282
rect 4142 3468 4146 3472
rect 4134 3218 4138 3222
rect 4086 3068 4090 3072
rect 4094 2988 4098 2992
rect 4078 2748 4082 2752
rect 4086 2738 4090 2742
rect 4078 2688 4082 2692
rect 4070 2408 4074 2412
rect 4110 2838 4114 2842
rect 4126 2828 4130 2832
rect 4158 4188 4162 4192
rect 4270 4848 4274 4852
rect 4222 4838 4226 4842
rect 4198 4528 4202 4532
rect 4182 4288 4186 4292
rect 4158 3518 4162 3522
rect 4150 2948 4154 2952
rect 4078 2188 4082 2192
rect 4110 2608 4114 2612
rect 4110 2498 4114 2502
rect 4046 1998 4050 2002
rect 4070 1918 4074 1922
rect 4046 1868 4050 1872
rect 4070 1768 4074 1772
rect 4054 1498 4058 1502
rect 4022 1148 4026 1152
rect 4030 778 4034 782
rect 3974 468 3978 472
rect 3922 303 3926 307
rect 3929 303 3930 307
rect 3930 303 3933 307
rect 4022 528 4026 532
rect 4110 2038 4114 2042
rect 4110 1628 4114 1632
rect 4086 1058 4090 1062
rect 4078 858 4082 862
rect 4110 1248 4114 1252
rect 4086 648 4090 652
rect 4134 2548 4138 2552
rect 4190 4128 4194 4132
rect 4214 4128 4218 4132
rect 4246 4448 4250 4452
rect 4262 4328 4266 4332
rect 4238 4118 4242 4122
rect 4230 3818 4234 3822
rect 4190 3668 4194 3672
rect 4198 3658 4202 3662
rect 4190 3628 4194 3632
rect 4182 3418 4186 3422
rect 4190 3388 4194 3392
rect 4198 3308 4202 3312
rect 4174 3088 4178 3092
rect 4174 3058 4178 3062
rect 4174 2888 4178 2892
rect 4174 2138 4178 2142
rect 4142 2108 4146 2112
rect 4174 2078 4178 2082
rect 4150 2068 4154 2072
rect 4150 2038 4154 2042
rect 4174 1818 4178 1822
rect 4190 2958 4194 2962
rect 4214 3258 4218 3262
rect 4238 3678 4242 3682
rect 4278 4548 4282 4552
rect 4426 4803 4430 4807
rect 4433 4803 4434 4807
rect 4434 4803 4437 4807
rect 4426 4603 4430 4607
rect 4433 4603 4434 4607
rect 4434 4603 4437 4607
rect 4342 4358 4346 4362
rect 4302 4338 4306 4342
rect 4270 3658 4274 3662
rect 4254 3058 4258 3062
rect 4214 2668 4218 2672
rect 4190 2618 4194 2622
rect 4190 2268 4194 2272
rect 4190 1978 4194 1982
rect 4190 1908 4194 1912
rect 4182 1758 4186 1762
rect 4174 1718 4178 1722
rect 4142 1488 4146 1492
rect 4158 1388 4162 1392
rect 4190 1648 4194 1652
rect 4198 1558 4202 1562
rect 4198 1538 4202 1542
rect 4190 1468 4194 1472
rect 4166 1188 4170 1192
rect 4174 1168 4178 1172
rect 4174 1048 4178 1052
rect 4134 1038 4138 1042
rect 4142 1028 4146 1032
rect 4174 838 4178 842
rect 4166 808 4170 812
rect 4118 658 4122 662
rect 4110 458 4114 462
rect 3998 258 4002 262
rect 3974 138 3978 142
rect 4062 138 4066 142
rect 3922 103 3926 107
rect 3929 103 3930 107
rect 3930 103 3933 107
rect 3894 88 3898 92
rect 3910 68 3914 72
rect 4166 448 4170 452
rect 4238 2488 4242 2492
rect 4230 2408 4234 2412
rect 4310 3608 4314 3612
rect 4318 3588 4322 3592
rect 4318 3248 4322 3252
rect 4286 2858 4290 2862
rect 4278 2748 4282 2752
rect 4286 2578 4290 2582
rect 4278 2538 4282 2542
rect 4302 2698 4306 2702
rect 4302 2648 4306 2652
rect 4302 2528 4306 2532
rect 4254 2448 4258 2452
rect 4238 2258 4242 2262
rect 4214 1988 4218 1992
rect 4230 1998 4234 2002
rect 4222 1788 4226 1792
rect 4246 1958 4250 1962
rect 4246 1828 4250 1832
rect 4238 1678 4242 1682
rect 4246 1638 4250 1642
rect 4214 1558 4218 1562
rect 4230 1558 4234 1562
rect 4214 1348 4218 1352
rect 4206 1128 4210 1132
rect 4238 1538 4242 1542
rect 4206 988 4210 992
rect 4278 2208 4282 2212
rect 4350 3988 4354 3992
rect 4342 3878 4346 3882
rect 4426 4403 4430 4407
rect 4433 4403 4434 4407
rect 4434 4403 4437 4407
rect 4406 4288 4410 4292
rect 4398 4238 4402 4242
rect 4374 3818 4378 3822
rect 4334 3258 4338 3262
rect 4334 3248 4338 3252
rect 4382 3318 4386 3322
rect 4342 2768 4346 2772
rect 4350 2758 4354 2762
rect 4326 2528 4330 2532
rect 4302 2098 4306 2102
rect 4366 2958 4370 2962
rect 4358 2628 4362 2632
rect 4350 2418 4354 2422
rect 4326 2148 4330 2152
rect 4342 2108 4346 2112
rect 4318 2088 4322 2092
rect 4326 2088 4330 2092
rect 4310 2028 4314 2032
rect 4318 1838 4322 1842
rect 4318 1568 4322 1572
rect 4318 1538 4322 1542
rect 4278 1318 4282 1322
rect 4278 1278 4282 1282
rect 4262 1258 4266 1262
rect 4294 1138 4298 1142
rect 4262 848 4266 852
rect 4206 648 4210 652
rect 4342 2058 4346 2062
rect 4350 2028 4354 2032
rect 4350 1938 4354 1942
rect 4334 1558 4338 1562
rect 4326 1268 4330 1272
rect 4398 3678 4402 3682
rect 4426 4203 4430 4207
rect 4433 4203 4434 4207
rect 4434 4203 4437 4207
rect 4426 4003 4430 4007
rect 4433 4003 4434 4007
rect 4434 4003 4437 4007
rect 4426 3803 4430 3807
rect 4433 3803 4434 3807
rect 4434 3803 4437 3807
rect 4462 3888 4466 3892
rect 4446 3618 4450 3622
rect 4426 3603 4430 3607
rect 4433 3603 4434 3607
rect 4434 3603 4437 3607
rect 4414 3458 4418 3462
rect 4426 3403 4430 3407
rect 4433 3403 4434 3407
rect 4434 3403 4437 3407
rect 4426 3203 4430 3207
rect 4433 3203 4434 3207
rect 4434 3203 4437 3207
rect 4414 3158 4418 3162
rect 4486 4018 4490 4022
rect 4494 3978 4498 3982
rect 4526 4368 4530 4372
rect 4518 4018 4522 4022
rect 4502 3548 4506 3552
rect 4494 3538 4498 3542
rect 4566 4748 4570 4752
rect 4558 4258 4562 4262
rect 4550 3758 4554 3762
rect 4534 3548 4538 3552
rect 4414 3118 4418 3122
rect 4426 3003 4430 3007
rect 4433 3003 4434 3007
rect 4434 3003 4437 3007
rect 4398 2938 4402 2942
rect 4398 2878 4402 2882
rect 4390 2678 4394 2682
rect 4374 2518 4378 2522
rect 4382 2138 4386 2142
rect 4374 2038 4378 2042
rect 4358 1538 4362 1542
rect 4422 2948 4426 2952
rect 4426 2803 4430 2807
rect 4433 2803 4434 2807
rect 4434 2803 4437 2807
rect 4426 2603 4430 2607
rect 4433 2603 4434 2607
rect 4434 2603 4437 2607
rect 4430 2538 4434 2542
rect 4414 2478 4418 2482
rect 4430 2458 4434 2462
rect 4406 2208 4410 2212
rect 4426 2403 4430 2407
rect 4433 2403 4434 2407
rect 4434 2403 4437 2407
rect 4502 3348 4506 3352
rect 4486 3288 4490 3292
rect 4502 3268 4506 3272
rect 4478 3258 4482 3262
rect 4494 3258 4498 3262
rect 4534 3318 4538 3322
rect 4462 2718 4466 2722
rect 4470 2548 4474 2552
rect 4426 2203 4430 2207
rect 4433 2203 4434 2207
rect 4434 2203 4437 2207
rect 4414 2108 4418 2112
rect 4426 2003 4430 2007
rect 4433 2003 4434 2007
rect 4434 2003 4437 2007
rect 4414 1808 4418 1812
rect 4426 1803 4430 1807
rect 4433 1803 4434 1807
rect 4434 1803 4437 1807
rect 4414 1798 4418 1802
rect 4406 1608 4410 1612
rect 4382 1578 4386 1582
rect 4398 1578 4402 1582
rect 4366 1528 4370 1532
rect 4358 1498 4362 1502
rect 4398 1568 4402 1572
rect 4406 1548 4410 1552
rect 4390 1538 4394 1542
rect 4374 1428 4378 1432
rect 4398 1498 4402 1502
rect 4406 1478 4410 1482
rect 4426 1603 4430 1607
rect 4433 1603 4434 1607
rect 4434 1603 4437 1607
rect 4426 1403 4430 1407
rect 4433 1403 4434 1407
rect 4434 1403 4437 1407
rect 4462 2428 4466 2432
rect 4454 1998 4458 2002
rect 4454 1488 4458 1492
rect 4446 1358 4450 1362
rect 4406 1328 4410 1332
rect 4326 1248 4330 1252
rect 4326 658 4330 662
rect 4358 1118 4362 1122
rect 4374 1058 4378 1062
rect 4390 868 4394 872
rect 4374 768 4378 772
rect 2734 58 2738 62
rect 2910 58 2914 62
rect 2966 58 2970 62
rect 3390 58 3394 62
rect 4426 1203 4430 1207
rect 4433 1203 4434 1207
rect 4434 1203 4437 1207
rect 4426 1003 4430 1007
rect 4433 1003 4434 1007
rect 4434 1003 4437 1007
rect 4454 1028 4458 1032
rect 4414 958 4418 962
rect 4426 803 4430 807
rect 4433 803 4434 807
rect 4434 803 4437 807
rect 4494 2958 4498 2962
rect 4526 2938 4530 2942
rect 4486 2578 4490 2582
rect 4478 2258 4482 2262
rect 4470 1468 4474 1472
rect 4470 1368 4474 1372
rect 4510 2908 4514 2912
rect 4566 3528 4570 3532
rect 4542 2878 4546 2882
rect 4534 2858 4538 2862
rect 4526 2848 4530 2852
rect 4502 2678 4506 2682
rect 4622 4458 4626 4462
rect 4662 4658 4666 4662
rect 4622 4328 4626 4332
rect 4638 4288 4642 4292
rect 4630 4238 4634 4242
rect 4614 3958 4618 3962
rect 4614 3938 4618 3942
rect 4574 3338 4578 3342
rect 4558 3298 4562 3302
rect 4566 3158 4570 3162
rect 4534 2648 4538 2652
rect 4494 2548 4498 2552
rect 4502 1778 4506 1782
rect 4550 2688 4554 2692
rect 4534 2088 4538 2092
rect 4526 1668 4530 1672
rect 4494 1508 4498 1512
rect 4486 948 4490 952
rect 4534 1418 4538 1422
rect 4390 478 4394 482
rect 4426 603 4430 607
rect 4433 603 4434 607
rect 4434 603 4437 607
rect 4426 403 4430 407
rect 4433 403 4434 407
rect 4434 403 4437 407
rect 4426 203 4430 207
rect 4433 203 4434 207
rect 4434 203 4437 207
rect 4430 128 4434 132
rect 4518 1358 4522 1362
rect 4566 3148 4570 3152
rect 4558 2288 4562 2292
rect 4582 2908 4586 2912
rect 4574 2678 4578 2682
rect 4638 4228 4642 4232
rect 4630 3758 4634 3762
rect 4606 3068 4610 3072
rect 4598 2858 4602 2862
rect 4582 2248 4586 2252
rect 4566 1418 4570 1422
rect 4590 1888 4594 1892
rect 4614 2688 4618 2692
rect 4614 2588 4618 2592
rect 4606 2248 4610 2252
rect 4630 3638 4634 3642
rect 4646 3638 4650 3642
rect 4630 3548 4634 3552
rect 4670 4298 4674 4302
rect 4678 3748 4682 3752
rect 4630 2718 4634 2722
rect 4622 2098 4626 2102
rect 4606 2058 4610 2062
rect 4606 2018 4610 2022
rect 4622 1998 4626 2002
rect 4582 1678 4586 1682
rect 4590 1568 4594 1572
rect 4598 1538 4602 1542
rect 4582 1378 4586 1382
rect 4638 2138 4642 2142
rect 4702 4558 4706 4562
rect 4710 4118 4714 4122
rect 4694 3838 4698 3842
rect 4686 3468 4690 3472
rect 4678 3438 4682 3442
rect 4670 2978 4674 2982
rect 4654 2738 4658 2742
rect 4686 2758 4690 2762
rect 4686 2358 4690 2362
rect 4702 2958 4706 2962
rect 4702 2738 4706 2742
rect 4694 2258 4698 2262
rect 4654 2148 4658 2152
rect 4662 2058 4666 2062
rect 4670 2048 4674 2052
rect 4662 1588 4666 1592
rect 4718 2048 4722 2052
rect 4742 3218 4746 3222
rect 4750 3168 4754 3172
rect 4766 2678 4770 2682
rect 4830 4258 4834 4262
rect 4822 4248 4826 4252
rect 4806 4238 4810 4242
rect 4782 2768 4786 2772
rect 4766 2658 4770 2662
rect 4758 2648 4762 2652
rect 4734 2438 4738 2442
rect 4750 2428 4754 2432
rect 4774 2448 4778 2452
rect 4822 2918 4826 2922
rect 4846 3728 4850 3732
rect 4854 3368 4858 3372
rect 4838 3278 4842 3282
rect 4846 3228 4850 3232
rect 4886 3928 4890 3932
rect 4878 3508 4882 3512
rect 4870 3258 4874 3262
rect 4862 3248 4866 3252
rect 4862 3228 4866 3232
rect 4862 3148 4866 3152
rect 4878 2958 4882 2962
rect 4830 2878 4834 2882
rect 4830 2868 4834 2872
rect 4822 2858 4826 2862
rect 4798 2478 4802 2482
rect 4798 2438 4802 2442
rect 4774 2418 4778 2422
rect 4766 2278 4770 2282
rect 4758 2128 4762 2132
rect 4702 1958 4706 1962
rect 4678 1818 4682 1822
rect 4694 1658 4698 1662
rect 4718 1688 4722 1692
rect 4622 1558 4626 1562
rect 4622 1508 4626 1512
rect 4622 1388 4626 1392
rect 4574 1288 4578 1292
rect 4534 1038 4538 1042
rect 4590 1188 4594 1192
rect 4598 1138 4602 1142
rect 4582 548 4586 552
rect 4542 278 4546 282
rect 4646 1168 4650 1172
rect 4622 768 4626 772
rect 4654 668 4658 672
rect 4694 1548 4698 1552
rect 4678 1258 4682 1262
rect 4670 1138 4674 1142
rect 4670 678 4674 682
rect 4718 1358 4722 1362
rect 4702 968 4706 972
rect 4742 1518 4746 1522
rect 4734 1148 4738 1152
rect 4734 1128 4738 1132
rect 4782 1928 4786 1932
rect 4750 958 4754 962
rect 4574 68 4578 72
rect 4830 2848 4834 2852
rect 4830 2698 4834 2702
rect 4886 2868 4890 2872
rect 4878 2848 4882 2852
rect 4878 2758 4882 2762
rect 4894 2718 4898 2722
rect 4886 2618 4890 2622
rect 4854 1898 4858 1902
rect 4830 1678 4834 1682
rect 4854 1678 4858 1682
rect 4814 1578 4818 1582
rect 4806 1418 4810 1422
rect 4806 1368 4810 1372
rect 4870 1658 4874 1662
rect 4894 1468 4898 1472
rect 4886 1118 4890 1122
rect 4862 748 4866 752
rect 4838 478 4842 482
rect 4830 118 4834 122
rect 4886 658 4890 662
rect 4886 558 4890 562
rect 4886 478 4890 482
rect 4926 5048 4930 5052
rect 4910 5038 4914 5042
rect 5142 5018 5146 5022
rect 5006 4918 5010 4922
rect 4938 4903 4942 4907
rect 4945 4903 4946 4907
rect 4946 4903 4949 4907
rect 4938 4703 4942 4707
rect 4945 4703 4946 4707
rect 4946 4703 4949 4707
rect 4938 4503 4942 4507
rect 4945 4503 4946 4507
rect 4946 4503 4949 4507
rect 4958 4478 4962 4482
rect 4938 4303 4942 4307
rect 4945 4303 4946 4307
rect 4946 4303 4949 4307
rect 4938 4103 4942 4107
rect 4945 4103 4946 4107
rect 4946 4103 4949 4107
rect 4938 3903 4942 3907
rect 4945 3903 4946 3907
rect 4946 3903 4949 3907
rect 4938 3703 4942 3707
rect 4945 3703 4946 3707
rect 4946 3703 4949 3707
rect 4950 3678 4954 3682
rect 4938 3503 4942 3507
rect 4945 3503 4946 3507
rect 4946 3503 4949 3507
rect 4918 3368 4922 3372
rect 4910 3268 4914 3272
rect 4910 3148 4914 3152
rect 4910 3078 4914 3082
rect 4910 2988 4914 2992
rect 4910 2758 4914 2762
rect 4918 2718 4922 2722
rect 4918 2378 4922 2382
rect 4938 3303 4942 3307
rect 4945 3303 4946 3307
rect 4946 3303 4949 3307
rect 4938 3103 4942 3107
rect 4945 3103 4946 3107
rect 4946 3103 4949 3107
rect 4966 3118 4970 3122
rect 4938 2903 4942 2907
rect 4945 2903 4946 2907
rect 4946 2903 4949 2907
rect 4958 2878 4962 2882
rect 4938 2703 4942 2707
rect 4945 2703 4946 2707
rect 4946 2703 4949 2707
rect 4938 2503 4942 2507
rect 4945 2503 4946 2507
rect 4946 2503 4949 2507
rect 4966 2738 4970 2742
rect 4938 2303 4942 2307
rect 4945 2303 4946 2307
rect 4946 2303 4949 2307
rect 4918 2108 4922 2112
rect 4938 2103 4942 2107
rect 4945 2103 4946 2107
rect 4946 2103 4949 2107
rect 4938 1903 4942 1907
rect 4945 1903 4946 1907
rect 4946 1903 4949 1907
rect 4958 1808 4962 1812
rect 4938 1703 4942 1707
rect 4945 1703 4946 1707
rect 4946 1703 4949 1707
rect 4938 1503 4942 1507
rect 4945 1503 4946 1507
rect 4946 1503 4949 1507
rect 4926 1468 4930 1472
rect 4918 1358 4922 1362
rect 4938 1303 4942 1307
rect 4945 1303 4946 1307
rect 4946 1303 4949 1307
rect 4938 1103 4942 1107
rect 4945 1103 4946 1107
rect 4946 1103 4949 1107
rect 4938 903 4942 907
rect 4945 903 4946 907
rect 4946 903 4949 907
rect 4938 703 4942 707
rect 4945 703 4946 707
rect 4946 703 4949 707
rect 4926 678 4930 682
rect 4938 503 4942 507
rect 4945 503 4946 507
rect 4946 503 4949 507
rect 4926 478 4930 482
rect 4990 4558 4994 4562
rect 4998 4528 5002 4532
rect 4990 4168 4994 4172
rect 4982 3958 4986 3962
rect 5006 4168 5010 4172
rect 4990 3948 4994 3952
rect 4982 3938 4986 3942
rect 4990 3938 4994 3942
rect 4998 3718 5002 3722
rect 5022 4828 5026 4832
rect 5062 4868 5066 4872
rect 5046 4588 5050 4592
rect 5038 4378 5042 4382
rect 5030 4288 5034 4292
rect 5022 3928 5026 3932
rect 5054 4258 5058 4262
rect 5054 3968 5058 3972
rect 5038 3948 5042 3952
rect 5022 3758 5026 3762
rect 5014 3688 5018 3692
rect 4990 3378 4994 3382
rect 5006 3368 5010 3372
rect 4990 3188 4994 3192
rect 4982 3088 4986 3092
rect 5014 3118 5018 3122
rect 4998 2918 5002 2922
rect 5022 2988 5026 2992
rect 5014 2758 5018 2762
rect 5006 2648 5010 2652
rect 4990 2628 4994 2632
rect 4998 2058 5002 2062
rect 5046 3168 5050 3172
rect 5046 3158 5050 3162
rect 5046 2688 5050 2692
rect 5046 2668 5050 2672
rect 5038 2358 5042 2362
rect 5030 2158 5034 2162
rect 5062 2818 5066 2822
rect 5062 2808 5066 2812
rect 5062 2358 5066 2362
rect 4966 1368 4970 1372
rect 4966 1358 4970 1362
rect 4998 1428 5002 1432
rect 4982 1138 4986 1142
rect 4974 948 4978 952
rect 4938 303 4942 307
rect 4945 303 4946 307
rect 4946 303 4949 307
rect 4958 278 4962 282
rect 4894 128 4898 132
rect 4938 103 4942 107
rect 4945 103 4946 107
rect 4946 103 4949 107
rect 4910 88 4914 92
rect 4822 68 4826 72
rect 4990 748 4994 752
rect 4990 478 4994 482
rect 5006 668 5010 672
rect 5038 1878 5042 1882
rect 5038 1868 5042 1872
rect 5030 1768 5034 1772
rect 5054 1888 5058 1892
rect 5078 3188 5082 3192
rect 5094 4118 5098 4122
rect 5110 3998 5114 4002
rect 5150 4628 5154 4632
rect 5142 4378 5146 4382
rect 5134 4118 5138 4122
rect 5182 4718 5186 4722
rect 5166 4548 5170 4552
rect 5182 4448 5186 4452
rect 5174 4318 5178 4322
rect 5174 4308 5178 4312
rect 5150 4108 5154 4112
rect 5102 3218 5106 3222
rect 5094 3178 5098 3182
rect 5094 2828 5098 2832
rect 5094 2818 5098 2822
rect 5086 2718 5090 2722
rect 5086 2698 5090 2702
rect 5078 2638 5082 2642
rect 5086 2248 5090 2252
rect 5070 1568 5074 1572
rect 5070 1228 5074 1232
rect 5038 658 5042 662
rect 5070 958 5074 962
rect 5022 278 5026 282
rect 4998 268 5002 272
rect 5070 658 5074 662
rect 5126 3758 5130 3762
rect 5134 3718 5138 3722
rect 5126 3708 5130 3712
rect 5118 3688 5122 3692
rect 5126 3508 5130 3512
rect 5126 3468 5130 3472
rect 5118 2978 5122 2982
rect 5110 2848 5114 2852
rect 5110 2828 5114 2832
rect 5102 2548 5106 2552
rect 5102 2428 5106 2432
rect 5118 2548 5122 2552
rect 5110 2188 5114 2192
rect 5094 1958 5098 1962
rect 5094 1928 5098 1932
rect 5102 1878 5106 1882
rect 5102 1718 5106 1722
rect 5134 3188 5138 3192
rect 5126 2188 5130 2192
rect 5118 1878 5122 1882
rect 5110 1428 5114 1432
rect 5094 1118 5098 1122
rect 5126 1728 5130 1732
rect 5102 728 5106 732
rect 5158 3998 5162 4002
rect 5166 3928 5170 3932
rect 5182 4068 5186 4072
rect 5198 4328 5202 4332
rect 5198 4318 5202 4322
rect 5158 3698 5162 3702
rect 5158 3688 5162 3692
rect 5150 2968 5154 2972
rect 5142 2848 5146 2852
rect 5142 2488 5146 2492
rect 5174 2808 5178 2812
rect 5142 2248 5146 2252
rect 5126 978 5130 982
rect 5014 258 5018 262
rect 5086 188 5090 192
rect 5038 78 5042 82
rect 5134 578 5138 582
rect 5150 1498 5154 1502
rect 5174 2318 5178 2322
rect 5190 3848 5194 3852
rect 5198 3168 5202 3172
rect 5230 4788 5234 4792
rect 5238 4698 5242 4702
rect 5214 4128 5218 4132
rect 5214 4108 5218 4112
rect 5214 3178 5218 3182
rect 5198 2898 5202 2902
rect 5190 2828 5194 2832
rect 5206 2858 5210 2862
rect 5198 2808 5202 2812
rect 5190 2568 5194 2572
rect 5190 2498 5194 2502
rect 5182 2168 5186 2172
rect 5182 2138 5186 2142
rect 5182 2108 5186 2112
rect 5158 1428 5162 1432
rect 5166 1158 5170 1162
rect 5182 1498 5186 1502
rect 5206 1698 5210 1702
rect 5190 1168 5194 1172
rect 5174 1138 5178 1142
rect 5158 1068 5162 1072
rect 5190 978 5194 982
rect 5182 858 5186 862
rect 5182 768 5186 772
rect 5182 648 5186 652
rect 5174 58 5178 62
rect 5254 4858 5258 4862
rect 5246 3868 5250 3872
rect 5238 3858 5242 3862
rect 5230 3118 5234 3122
rect 5222 2838 5226 2842
rect 5222 2098 5226 2102
rect 5222 1518 5226 1522
rect 5246 2558 5250 2562
rect 5238 2548 5242 2552
rect 5246 2328 5250 2332
rect 5278 3688 5282 3692
rect 5270 2318 5274 2322
rect 5238 2128 5242 2132
rect 5254 2138 5258 2142
rect 5246 2118 5250 2122
rect 5238 1858 5242 1862
rect 5254 1858 5258 1862
rect 5238 1518 5242 1522
rect 5214 318 5218 322
rect 5198 288 5202 292
rect 5246 1178 5250 1182
rect 5238 888 5242 892
rect 5230 438 5234 442
rect 5294 3248 5298 3252
rect 5294 2888 5298 2892
rect 5286 2568 5290 2572
rect 5286 2388 5290 2392
rect 5294 2318 5298 2322
rect 5278 2058 5282 2062
rect 5270 988 5274 992
rect 5302 2238 5306 2242
rect 5302 2228 5306 2232
rect 5294 1908 5298 1912
rect 5286 1158 5290 1162
rect 5278 978 5282 982
rect 5270 758 5274 762
rect 5270 468 5274 472
rect 5286 318 5290 322
rect 5246 158 5250 162
rect 5278 148 5282 152
rect 5262 138 5266 142
rect 5222 68 5226 72
rect 330 3 334 7
rect 337 3 338 7
rect 338 3 341 7
rect 1354 3 1358 7
rect 1361 3 1362 7
rect 1362 3 1365 7
rect 2386 3 2390 7
rect 2393 3 2394 7
rect 2394 3 2397 7
rect 3402 3 3406 7
rect 3409 3 3410 7
rect 3410 3 3413 7
rect 4426 3 4430 7
rect 4433 3 4434 7
rect 4434 3 4437 7
<< metal5 >>
rect 854 5103 857 5107
rect 853 5102 858 5103
rect 863 5102 864 5107
rect 1878 5103 1881 5107
rect 1877 5102 1882 5103
rect 1887 5102 1888 5107
rect 2894 5103 2897 5107
rect 2893 5102 2898 5103
rect 2903 5102 2904 5107
rect 3926 5103 3929 5107
rect 3925 5102 3930 5103
rect 3935 5102 3936 5107
rect 4942 5103 4945 5107
rect 4941 5102 4946 5103
rect 4951 5102 4952 5107
rect 4506 5078 4541 5081
rect 4490 5068 4509 5071
rect 170 5058 198 5061
rect 4586 5058 4621 5061
rect 4926 5052 4929 5057
rect 1786 5048 3950 5051
rect 4910 5042 4913 5047
rect 4850 5018 5142 5021
rect 334 5003 337 5007
rect 333 5002 338 5003
rect 343 5002 344 5007
rect 1358 5003 1361 5007
rect 1357 5002 1362 5003
rect 1367 5002 1368 5007
rect 2390 5003 2393 5007
rect 2389 5002 2394 5003
rect 2399 5002 2400 5007
rect 3406 5003 3409 5007
rect 3405 5002 3410 5003
rect 3415 5002 3416 5007
rect 4430 5003 4433 5007
rect 4429 5002 4434 5003
rect 4439 5002 4440 5007
rect 474 4958 742 4961
rect 194 4948 774 4951
rect 1466 4948 1726 4951
rect 202 4928 870 4931
rect 5006 4928 5069 4931
rect 5006 4922 5009 4928
rect 854 4903 857 4907
rect 853 4902 858 4903
rect 863 4902 864 4907
rect 1878 4903 1881 4907
rect 1877 4902 1882 4903
rect 1887 4902 1888 4907
rect 2894 4903 2897 4907
rect 2893 4902 2898 4903
rect 2903 4902 2904 4907
rect 3926 4903 3929 4907
rect 3925 4902 3930 4903
rect 3935 4902 3936 4907
rect 4942 4903 4945 4907
rect 4941 4902 4946 4903
rect 4951 4902 4952 4907
rect 546 4878 702 4881
rect 5010 4868 5062 4871
rect 794 4858 870 4861
rect 3266 4858 4137 4861
rect 4134 4852 4137 4858
rect 4818 4858 5254 4861
rect 250 4848 734 4851
rect 4138 4848 4270 4851
rect 3442 4838 4222 4841
rect 3586 4828 4134 4831
rect 5026 4828 5037 4831
rect 334 4803 337 4807
rect 333 4802 338 4803
rect 343 4802 344 4807
rect 1358 4803 1361 4807
rect 1357 4802 1362 4803
rect 1367 4802 1368 4807
rect 2390 4803 2393 4807
rect 2389 4802 2394 4803
rect 2399 4802 2400 4807
rect 3406 4803 3409 4807
rect 3405 4802 3410 4803
rect 3415 4802 3416 4807
rect 4430 4803 4433 4807
rect 4429 4802 4434 4803
rect 4439 4802 4440 4807
rect 5090 4788 5230 4791
rect 434 4758 638 4761
rect 734 4761 737 4768
rect 642 4758 737 4761
rect 1458 4748 1614 4751
rect 1722 4748 2478 4751
rect 3074 4748 4566 4751
rect 642 4728 910 4731
rect 2866 4728 2878 4731
rect 4834 4718 5182 4721
rect 854 4703 857 4707
rect 853 4702 858 4703
rect 863 4702 864 4707
rect 1878 4703 1881 4707
rect 1877 4702 1882 4703
rect 1887 4702 1888 4707
rect 2894 4703 2897 4707
rect 2893 4702 2898 4703
rect 2903 4702 2904 4707
rect 3926 4703 3929 4707
rect 3925 4702 3930 4703
rect 3935 4702 3936 4707
rect 4942 4703 4945 4707
rect 4941 4702 4946 4703
rect 4951 4702 4952 4707
rect 5242 4698 5245 4701
rect 2906 4668 3366 4671
rect 2874 4658 4662 4661
rect 5138 4638 5153 4641
rect 5150 4632 5153 4638
rect 582 4618 694 4621
rect 582 4612 585 4618
rect 334 4603 337 4607
rect 333 4602 338 4603
rect 343 4602 344 4607
rect 1358 4603 1361 4607
rect 1357 4602 1362 4603
rect 1367 4602 1368 4607
rect 2390 4603 2393 4607
rect 2389 4602 2394 4603
rect 2399 4602 2400 4607
rect 3406 4603 3409 4607
rect 3405 4602 3410 4603
rect 3415 4602 3416 4607
rect 4430 4603 4433 4607
rect 4429 4602 4434 4603
rect 4439 4602 4440 4607
rect 5026 4588 5046 4591
rect 450 4558 598 4561
rect 1150 4558 1358 4561
rect 4142 4561 4145 4568
rect 3946 4558 4145 4561
rect 4178 4558 4702 4561
rect 1150 4552 1153 4558
rect 4978 4558 4990 4561
rect 2794 4548 2950 4551
rect 3538 4548 3958 4551
rect 4082 4548 4278 4551
rect 5166 4542 5169 4548
rect 378 4538 438 4541
rect 2834 4538 3870 4541
rect 3970 4538 4142 4541
rect 4994 4538 5001 4541
rect 4998 4532 5001 4538
rect 2862 4528 3462 4531
rect 4106 4528 4198 4531
rect 2862 4522 2865 4528
rect 854 4503 857 4507
rect 853 4502 858 4503
rect 863 4502 864 4507
rect 1878 4503 1881 4507
rect 1877 4502 1882 4503
rect 1887 4502 1888 4507
rect 2894 4503 2897 4507
rect 2893 4502 2898 4503
rect 2903 4502 2904 4507
rect 3926 4503 3929 4507
rect 3925 4502 3930 4503
rect 3935 4502 3936 4507
rect 4942 4503 4945 4507
rect 4941 4502 4946 4503
rect 4951 4502 4952 4507
rect 4958 4472 4961 4478
rect 722 4458 1070 4461
rect 2066 4458 2070 4461
rect 2754 4458 3118 4461
rect 3530 4458 4622 4461
rect 5182 4458 5197 4461
rect 5182 4452 5185 4458
rect 890 4448 1190 4451
rect 1994 4448 2022 4451
rect 3458 4448 4246 4451
rect 3258 4438 3838 4441
rect 3842 4438 4102 4441
rect 2690 4428 3638 4431
rect 334 4403 337 4407
rect 333 4402 338 4403
rect 343 4402 344 4407
rect 1358 4403 1361 4407
rect 1357 4402 1362 4403
rect 1367 4402 1368 4407
rect 2390 4403 2393 4407
rect 2389 4402 2394 4403
rect 2399 4402 2400 4407
rect 3406 4403 3409 4407
rect 3405 4402 3410 4403
rect 3415 4402 3416 4407
rect 4430 4403 4433 4407
rect 4429 4402 4434 4403
rect 4439 4402 4440 4407
rect 5042 4378 5142 4381
rect 2562 4368 3934 4371
rect 3938 4368 4150 4371
rect 4154 4368 4526 4371
rect 1454 4362 1457 4368
rect 3130 4358 4093 4361
rect 4098 4358 4342 4361
rect 138 4348 798 4351
rect 2098 4348 3206 4351
rect 3346 4348 3398 4351
rect 490 4338 702 4341
rect 2522 4338 3886 4341
rect 3890 4338 4302 4341
rect 4866 4338 5201 4341
rect 5198 4332 5201 4338
rect 322 4328 566 4331
rect 3338 4328 4062 4331
rect 4266 4328 4622 4331
rect 5178 4318 5198 4321
rect 5178 4308 5277 4311
rect 854 4303 857 4307
rect 853 4302 858 4303
rect 863 4302 864 4307
rect 1878 4303 1881 4307
rect 1877 4302 1882 4303
rect 1887 4302 1888 4307
rect 2894 4303 2897 4307
rect 2893 4302 2898 4303
rect 2903 4302 2904 4307
rect 3926 4303 3929 4307
rect 3925 4302 3930 4303
rect 3935 4302 3936 4307
rect 4942 4303 4945 4307
rect 4941 4302 4946 4303
rect 4951 4302 4952 4307
rect 2050 4298 2838 4301
rect 4066 4298 4670 4301
rect 1466 4288 2077 4291
rect 3210 4288 4182 4291
rect 4410 4288 4638 4291
rect 5034 4288 5101 4291
rect 210 4278 614 4281
rect 2834 4278 2886 4281
rect 642 4268 734 4271
rect 1682 4268 1685 4271
rect 2474 4268 3174 4271
rect 5054 4262 5057 4267
rect 602 4258 782 4261
rect 1674 4258 2054 4261
rect 2090 4258 2573 4261
rect 2578 4258 3526 4261
rect 4562 4258 4830 4261
rect 3550 4252 3553 4258
rect 362 4248 646 4251
rect 778 4248 830 4251
rect 2950 4241 2953 4248
rect 4658 4248 4822 4251
rect 2002 4238 2953 4241
rect 2962 4238 3598 4241
rect 4402 4238 4630 4241
rect 4634 4238 4806 4241
rect 354 4228 814 4231
rect 2442 4228 4638 4231
rect 2570 4218 3486 4221
rect 334 4203 337 4207
rect 333 4202 338 4203
rect 343 4202 344 4207
rect 1358 4203 1361 4207
rect 1357 4202 1362 4203
rect 1367 4202 1368 4207
rect 2390 4203 2393 4207
rect 2389 4202 2394 4203
rect 2399 4202 2400 4207
rect 3406 4203 3409 4207
rect 3405 4202 3410 4203
rect 3415 4202 3416 4207
rect 4430 4203 4433 4207
rect 4429 4202 4434 4203
rect 4439 4202 4440 4207
rect 2858 4188 4158 4191
rect 386 4178 526 4181
rect 2458 4168 4653 4171
rect 4994 4168 5006 4171
rect 3038 4152 3041 4157
rect 1482 4148 2174 4151
rect 2202 4148 2926 4151
rect 1282 4138 1902 4141
rect 2122 4138 2254 4141
rect 2618 4138 3030 4141
rect 2770 4128 4190 4131
rect 4218 4128 4525 4131
rect 5214 4122 5217 4128
rect 1298 4118 1878 4121
rect 4042 4118 4238 4121
rect 4242 4118 4710 4121
rect 5098 4118 5134 4121
rect 1930 4108 2822 4111
rect 3042 4108 3910 4111
rect 5154 4108 5214 4111
rect 854 4103 857 4107
rect 853 4102 858 4103
rect 863 4102 864 4107
rect 1878 4103 1881 4107
rect 1877 4102 1882 4103
rect 1887 4102 1888 4107
rect 2894 4103 2897 4107
rect 2893 4102 2898 4103
rect 2903 4102 2904 4107
rect 3926 4103 3929 4107
rect 3925 4102 3930 4103
rect 3935 4102 3936 4107
rect 4942 4103 4945 4107
rect 4941 4102 4946 4103
rect 4951 4102 4952 4107
rect 1922 4088 2118 4091
rect 554 4078 3886 4081
rect 3890 4078 4142 4081
rect 5182 4078 5261 4081
rect 5182 4072 5185 4078
rect 1722 4068 1934 4071
rect 1602 4058 1694 4061
rect 1738 4058 1918 4061
rect 1966 4061 1969 4068
rect 1946 4058 1969 4061
rect 3018 4058 3510 4061
rect 1450 4038 1854 4041
rect 2546 4038 2854 4041
rect 2922 4038 3894 4041
rect 978 4028 3054 4031
rect 3058 4018 4070 4021
rect 4074 4018 4486 4021
rect 4522 4018 4589 4021
rect 2874 4008 3086 4011
rect 3210 4008 3261 4011
rect 334 4003 337 4007
rect 333 4002 338 4003
rect 343 4002 344 4007
rect 1358 4003 1361 4007
rect 1357 4002 1362 4003
rect 1367 4002 1368 4007
rect 2390 4003 2393 4007
rect 2389 4002 2394 4003
rect 2399 4002 2400 4007
rect 2686 4002 2689 4008
rect 3406 4003 3409 4007
rect 3405 4002 3410 4003
rect 3415 4002 3416 4007
rect 4430 4003 4433 4007
rect 4429 4002 4434 4003
rect 4439 4002 4440 4007
rect 1458 3998 1469 4001
rect 5114 3998 5117 4001
rect 5154 3998 5158 4001
rect 3386 3988 4350 3991
rect 578 3978 598 3981
rect 3186 3978 3638 3981
rect 3898 3978 4493 3981
rect 2858 3968 3790 3971
rect 5026 3968 5054 3971
rect 2042 3958 2134 3961
rect 3246 3958 3774 3961
rect 4618 3958 4685 3961
rect 3246 3951 3249 3958
rect 2082 3948 3249 3951
rect 3730 3948 3910 3951
rect 3486 3942 3489 3948
rect 4982 3942 4985 3958
rect 4994 3948 5038 3951
rect 1746 3938 2038 3941
rect 2194 3938 3485 3941
rect 3690 3938 4614 3941
rect 4994 3938 5037 3941
rect 2138 3928 2854 3931
rect 4890 3928 5022 3931
rect 5154 3928 5166 3931
rect 938 3918 1286 3921
rect 2018 3918 3398 3921
rect 854 3903 857 3907
rect 853 3902 858 3903
rect 863 3902 864 3907
rect 1878 3903 1881 3907
rect 1877 3902 1882 3903
rect 1887 3902 1888 3907
rect 2894 3903 2897 3907
rect 2893 3902 2898 3903
rect 2903 3902 2904 3907
rect 3926 3903 3929 3907
rect 3925 3902 3930 3903
rect 3935 3902 3936 3907
rect 4942 3903 4945 3907
rect 4941 3902 4946 3903
rect 4951 3902 4952 3907
rect 1066 3898 1865 3901
rect 1226 3888 1742 3891
rect 1862 3891 1865 3898
rect 1862 3888 3174 3891
rect 3522 3888 4462 3891
rect 1170 3878 1238 3881
rect 1786 3878 2142 3881
rect 3434 3878 4070 3881
rect 4074 3878 4078 3881
rect 4082 3878 4342 3881
rect 1090 3868 1182 3871
rect 1322 3868 1350 3871
rect 2002 3868 2006 3871
rect 2466 3868 2678 3871
rect 2682 3868 3766 3871
rect 5186 3868 5246 3871
rect 970 3858 1822 3861
rect 1930 3858 1965 3861
rect 1970 3858 2038 3861
rect 3298 3858 3718 3861
rect 5234 3858 5238 3861
rect 1898 3848 2973 3851
rect 2978 3848 3270 3851
rect 3530 3848 3798 3851
rect 3818 3848 3878 3851
rect 4994 3848 5190 3851
rect 114 3838 214 3841
rect 218 3838 462 3841
rect 1746 3838 2518 3841
rect 3074 3838 4694 3841
rect 4978 3838 4989 3841
rect 1418 3828 2878 3831
rect 3202 3828 3206 3831
rect 1002 3818 3382 3821
rect 3386 3818 4230 3821
rect 4234 3818 4374 3821
rect 334 3803 337 3807
rect 333 3802 338 3803
rect 343 3802 344 3807
rect 1358 3803 1361 3807
rect 1357 3802 1362 3803
rect 1367 3802 1368 3807
rect 2390 3803 2393 3807
rect 2389 3802 2394 3803
rect 2399 3802 2400 3807
rect 3406 3803 3409 3807
rect 3405 3802 3410 3803
rect 3415 3802 3416 3807
rect 4430 3803 4433 3807
rect 4429 3802 4434 3803
rect 4439 3802 4440 3807
rect 1946 3788 2390 3791
rect 2266 3778 2494 3781
rect 2930 3778 2934 3781
rect 2370 3768 3590 3771
rect 2090 3758 3046 3761
rect 3050 3758 3206 3761
rect 3994 3758 4550 3761
rect 4634 3758 4701 3761
rect 58 3748 86 3751
rect 1610 3748 2086 3751
rect 2786 3748 3150 3751
rect 3214 3751 3217 3758
rect 5026 3758 5126 3761
rect 3214 3748 3374 3751
rect 3602 3748 4678 3751
rect 1258 3738 1422 3741
rect 1618 3738 1622 3741
rect 1914 3738 3262 3741
rect 3538 3738 4006 3741
rect 922 3728 1278 3731
rect 1538 3728 2710 3731
rect 2882 3728 2926 3731
rect 3082 3728 3337 3731
rect 3346 3728 4846 3731
rect 1938 3718 2078 3721
rect 2162 3718 2173 3721
rect 2178 3718 2990 3721
rect 3334 3721 3337 3728
rect 3334 3718 3998 3721
rect 5002 3718 5005 3721
rect 5138 3718 5149 3721
rect 1066 3708 1069 3711
rect 2074 3708 2446 3711
rect 3362 3708 3902 3711
rect 5130 3708 5133 3711
rect 854 3703 857 3707
rect 853 3702 858 3703
rect 863 3702 864 3707
rect 1878 3703 1881 3707
rect 1877 3702 1882 3703
rect 1887 3702 1888 3707
rect 2894 3703 2897 3707
rect 2893 3702 2898 3703
rect 2903 3702 2904 3707
rect 3926 3703 3929 3707
rect 3925 3702 3930 3703
rect 3935 3702 3936 3707
rect 4942 3703 4945 3707
rect 4941 3702 4946 3703
rect 4951 3702 4952 3707
rect 1354 3688 1838 3691
rect 2654 3691 2657 3698
rect 2706 3698 2710 3701
rect 2994 3698 3542 3701
rect 5042 3698 5158 3701
rect 2654 3688 2966 3691
rect 3666 3688 3901 3691
rect 5010 3688 5014 3691
rect 5122 3688 5133 3691
rect 5162 3688 5165 3691
rect 1218 3678 1854 3681
rect 2418 3678 2662 3681
rect 2690 3678 3046 3681
rect 3354 3678 3598 3681
rect 3738 3678 4238 3681
rect 4242 3678 4398 3681
rect 4954 3678 4973 3681
rect 3310 3672 3313 3678
rect 5278 3681 5281 3688
rect 4978 3678 5281 3681
rect 634 3668 1246 3671
rect 2194 3668 2766 3671
rect 2938 3668 3030 3671
rect 3490 3668 3894 3671
rect 3906 3668 4190 3671
rect 722 3658 1118 3661
rect 3042 3658 3366 3661
rect 4202 3658 4270 3661
rect 754 3648 1741 3651
rect 1794 3648 1797 3651
rect 2442 3648 2797 3651
rect 2802 3648 2982 3651
rect 3170 3648 3174 3651
rect 3218 3648 3982 3651
rect 1058 3638 1117 3641
rect 1122 3638 2014 3641
rect 2066 3638 2662 3641
rect 2690 3638 4630 3641
rect 4650 3638 4669 3641
rect 1338 3628 1630 3631
rect 2106 3628 2109 3631
rect 2258 3628 2854 3631
rect 2858 3628 3254 3631
rect 3298 3628 4190 3631
rect 2170 3618 2566 3621
rect 2610 3618 3558 3621
rect 4162 3618 4446 3621
rect 2746 3608 2774 3611
rect 3450 3608 3990 3611
rect 4034 3608 4310 3611
rect 334 3603 337 3607
rect 333 3602 338 3603
rect 343 3602 344 3607
rect 1358 3603 1361 3607
rect 1357 3602 1362 3603
rect 1367 3602 1368 3607
rect 2390 3603 2393 3607
rect 2389 3602 2394 3603
rect 2399 3602 2400 3607
rect 3406 3603 3409 3607
rect 3405 3602 3410 3603
rect 3415 3602 3416 3607
rect 4430 3603 4433 3607
rect 4429 3602 4434 3603
rect 4439 3602 4440 3607
rect 1490 3598 2062 3601
rect 466 3588 1798 3591
rect 2258 3588 3222 3591
rect 3730 3588 4318 3591
rect 1642 3578 3030 3581
rect 3154 3578 3702 3581
rect 154 3568 1630 3571
rect 1650 3568 1662 3571
rect 1666 3568 2253 3571
rect 2266 3568 3126 3571
rect 3130 3568 3310 3571
rect 3314 3568 3702 3571
rect 1178 3558 1526 3561
rect 1746 3558 1790 3561
rect 1802 3558 2574 3561
rect 3570 3558 3830 3561
rect 5106 3558 5165 3561
rect 1850 3548 2590 3551
rect 2682 3548 3438 3551
rect 4070 3548 4502 3551
rect 4526 3548 4534 3551
rect 4538 3548 4630 3551
rect 4070 3542 4073 3548
rect 786 3538 1686 3541
rect 1698 3538 1790 3541
rect 3210 3538 3213 3541
rect 3102 3532 3105 3538
rect 3754 3538 4062 3541
rect 474 3528 566 3531
rect 866 3528 1022 3531
rect 1618 3528 2966 3531
rect 3202 3528 3446 3531
rect 4494 3531 4497 3538
rect 4494 3528 4566 3531
rect 1546 3518 1622 3521
rect 1666 3518 1678 3521
rect 3678 3521 3681 3528
rect 1690 3518 3681 3521
rect 3810 3518 4158 3521
rect 1538 3508 1822 3511
rect 2482 3508 2502 3511
rect 3106 3508 3470 3511
rect 854 3503 857 3507
rect 853 3502 858 3503
rect 863 3502 864 3507
rect 1878 3503 1881 3507
rect 1877 3502 1882 3503
rect 1887 3502 1888 3507
rect 2894 3503 2897 3507
rect 2893 3502 2898 3503
rect 2903 3502 2904 3507
rect 3926 3503 3929 3507
rect 3925 3502 3930 3503
rect 3935 3502 3936 3507
rect 4878 3502 4881 3508
rect 5026 3508 5126 3511
rect 4942 3503 4945 3507
rect 4941 3502 4946 3503
rect 4951 3502 4952 3507
rect 1810 3498 1822 3501
rect 1906 3498 1982 3501
rect 1986 3498 2670 3501
rect 3242 3498 3574 3501
rect 1178 3488 2246 3491
rect 2250 3488 2301 3491
rect 2306 3488 3566 3491
rect 3578 3488 3822 3491
rect 2714 3478 3206 3481
rect 3370 3478 4030 3481
rect 650 3468 897 3471
rect 1794 3468 3150 3471
rect 3178 3468 3646 3471
rect 4146 3468 4173 3471
rect 894 3462 897 3468
rect 1274 3458 1806 3461
rect 3174 3461 3177 3468
rect 4690 3468 4765 3471
rect 1858 3458 3177 3461
rect 5126 3461 5129 3468
rect 4418 3458 5129 3461
rect 402 3448 1198 3451
rect 1330 3448 1710 3451
rect 2602 3448 3206 3451
rect 3314 3448 4681 3451
rect 4678 3442 4681 3448
rect 1458 3438 1510 3441
rect 1786 3438 3110 3441
rect 3146 3438 4014 3441
rect 4018 3438 4022 3441
rect 658 3428 2022 3431
rect 2026 3428 3230 3431
rect 514 3418 2054 3421
rect 3018 3418 4182 3421
rect 4186 3418 4205 3421
rect 2246 3411 2249 3418
rect 1554 3408 2249 3411
rect 2410 3408 3038 3411
rect 334 3403 337 3407
rect 333 3402 338 3403
rect 343 3402 344 3407
rect 1358 3403 1361 3407
rect 1357 3402 1362 3403
rect 1367 3402 1368 3407
rect 2390 3403 2393 3407
rect 2389 3402 2394 3403
rect 2399 3402 2400 3407
rect 3406 3403 3409 3407
rect 3405 3402 3410 3403
rect 3415 3402 3416 3407
rect 4430 3403 4433 3407
rect 4429 3402 4434 3403
rect 4439 3402 4440 3407
rect 2794 3398 2806 3401
rect 3114 3398 3230 3401
rect 2642 3388 4190 3391
rect 4990 3382 4993 3387
rect 1946 3378 2246 3381
rect 2250 3378 2406 3381
rect 2506 3378 2910 3381
rect 2986 3378 3726 3381
rect 3730 3378 3997 3381
rect 1250 3368 2126 3371
rect 3386 3368 3718 3371
rect 4858 3368 4918 3371
rect 4994 3368 5006 3371
rect 570 3358 766 3361
rect 1578 3358 1902 3361
rect 2066 3358 2238 3361
rect 2242 3358 2438 3361
rect 2946 3358 4102 3361
rect 802 3348 886 3351
rect 2138 3348 2925 3351
rect 3042 3348 3574 3351
rect 4106 3348 4502 3351
rect 434 3338 1150 3341
rect 1330 3338 1774 3341
rect 2082 3338 2126 3341
rect 2626 3338 3446 3341
rect 4574 3332 4577 3338
rect 450 3328 1014 3331
rect 1018 3328 1645 3331
rect 2322 3328 2758 3331
rect 3098 3328 3606 3331
rect 738 3318 1574 3321
rect 2258 3318 2710 3321
rect 2738 3318 3014 3321
rect 3522 3318 4382 3321
rect 4386 3318 4534 3321
rect 1146 3308 1534 3311
rect 2330 3308 2333 3311
rect 3266 3308 3822 3311
rect 3982 3308 4198 3311
rect 854 3303 857 3307
rect 853 3302 858 3303
rect 863 3302 864 3307
rect 1878 3303 1881 3307
rect 1877 3302 1882 3303
rect 1887 3302 1888 3307
rect 2894 3303 2897 3307
rect 2893 3302 2898 3303
rect 2903 3302 2904 3307
rect 3926 3303 3929 3307
rect 3925 3302 3930 3303
rect 3935 3302 3936 3307
rect 3982 3302 3985 3308
rect 4942 3303 4945 3307
rect 4941 3302 4946 3303
rect 4951 3302 4952 3307
rect 2066 3298 2270 3301
rect 2274 3298 2854 3301
rect 4066 3298 4558 3301
rect 1746 3288 2486 3291
rect 2882 3288 4477 3291
rect 4482 3288 4486 3291
rect 1586 3278 2438 3281
rect 3298 3278 3302 3281
rect 4090 3278 4838 3281
rect 594 3268 750 3271
rect 1794 3268 2413 3271
rect 2418 3268 2550 3271
rect 2746 3268 2838 3271
rect 3306 3268 3350 3271
rect 3714 3268 4022 3271
rect 4506 3268 4910 3271
rect 730 3258 1430 3261
rect 2058 3258 2781 3261
rect 3818 3258 4214 3261
rect 4338 3258 4478 3261
rect 4498 3258 4870 3261
rect 5294 3252 5297 3257
rect 1466 3248 1534 3251
rect 2842 3248 4318 3251
rect 4338 3248 4862 3251
rect 1498 3238 1614 3241
rect 2042 3238 2086 3241
rect 3842 3238 4865 3241
rect 4862 3232 4865 3238
rect 474 3228 2014 3231
rect 2026 3228 2902 3231
rect 3658 3228 4605 3231
rect 4610 3228 4846 3231
rect 410 3218 1470 3221
rect 1474 3218 3462 3221
rect 3890 3218 3974 3221
rect 4138 3218 4742 3221
rect 5102 3212 5105 3218
rect 2410 3208 3142 3211
rect 334 3203 337 3207
rect 333 3202 338 3203
rect 343 3202 344 3207
rect 1358 3203 1361 3207
rect 1357 3202 1362 3203
rect 1367 3202 1368 3207
rect 2390 3203 2393 3207
rect 2389 3202 2394 3203
rect 2399 3202 2400 3207
rect 3406 3203 3409 3207
rect 3405 3202 3410 3203
rect 3415 3202 3416 3207
rect 4430 3203 4433 3207
rect 4429 3202 4434 3203
rect 4439 3202 4440 3207
rect 2474 3198 2542 3201
rect 2658 3198 2798 3201
rect 2802 3198 3374 3201
rect 2210 3188 2782 3191
rect 2946 3188 3942 3191
rect 4962 3188 4990 3191
rect 5082 3188 5134 3191
rect 5214 3182 5217 3187
rect 1722 3178 2150 3181
rect 2154 3178 2678 3181
rect 2914 3178 3102 3181
rect 5042 3178 5094 3181
rect 1410 3168 2822 3171
rect 3202 3168 4750 3171
rect 5042 3168 5046 3171
rect 5202 3168 5213 3171
rect 930 3158 1630 3161
rect 2010 3158 2406 3161
rect 2450 3158 2870 3161
rect 3458 3158 3846 3161
rect 4418 3158 4566 3161
rect 5050 3158 5277 3161
rect 1670 3151 1673 3158
rect 1186 3148 1673 3151
rect 2010 3148 2030 3151
rect 2114 3148 2118 3151
rect 2242 3148 2278 3151
rect 3030 3151 3033 3158
rect 2842 3148 3033 3151
rect 3042 3148 3046 3151
rect 4546 3148 4566 3151
rect 4866 3148 4910 3151
rect 946 3138 1462 3141
rect 1634 3138 1694 3141
rect 1786 3138 2622 3141
rect 594 3128 838 3131
rect 1138 3128 1406 3131
rect 1498 3128 1918 3131
rect 2274 3128 2654 3131
rect 3042 3128 3958 3131
rect 5230 3128 5277 3131
rect 4414 3122 4417 3127
rect 5230 3122 5233 3128
rect 1666 3118 2493 3121
rect 2858 3118 3182 3121
rect 4970 3118 5014 3121
rect 1522 3108 1702 3111
rect 2130 3108 2598 3111
rect 2602 3108 2838 3111
rect 854 3103 857 3107
rect 853 3102 858 3103
rect 863 3102 864 3107
rect 1878 3103 1881 3107
rect 1877 3102 1882 3103
rect 1887 3102 1888 3107
rect 2894 3103 2897 3107
rect 2893 3102 2898 3103
rect 2903 3102 2904 3107
rect 3926 3103 3929 3107
rect 3925 3102 3930 3103
rect 3935 3102 3936 3107
rect 4942 3103 4945 3107
rect 4941 3102 4946 3103
rect 4951 3102 4952 3107
rect 2226 3098 2622 3101
rect 2938 3098 3910 3101
rect 914 3088 1438 3091
rect 1570 3088 1726 3091
rect 2202 3088 2702 3091
rect 2706 3088 2990 3091
rect 3262 3088 3678 3091
rect 4034 3088 4174 3091
rect 1314 3078 1654 3081
rect 1658 3078 2349 3081
rect 3262 3081 3265 3088
rect 4898 3088 4982 3091
rect 2490 3078 3265 3081
rect 4910 3082 4913 3088
rect 1898 3068 2486 3071
rect 2530 3068 2734 3071
rect 2882 3068 3262 3071
rect 3666 3068 4086 3071
rect 1222 3061 1225 3068
rect 1222 3058 1334 3061
rect 1602 3058 1854 3061
rect 1954 3058 2022 3061
rect 2026 3058 2669 3061
rect 2830 3061 2833 3068
rect 2830 3058 3086 3061
rect 3634 3058 4174 3061
rect 4606 3061 4609 3068
rect 4258 3058 4609 3061
rect 1458 3048 1870 3051
rect 1922 3048 2790 3051
rect 2938 3048 3742 3051
rect 3746 3048 4061 3051
rect 1922 3038 3334 3041
rect 1690 3028 2125 3031
rect 2130 3028 2134 3031
rect 2498 3028 3054 3031
rect 3066 3028 3430 3031
rect 1098 3018 2646 3021
rect 2674 3018 3382 3021
rect 1522 3008 1854 3011
rect 1858 3008 2278 3011
rect 3306 3008 3341 3011
rect 334 3003 337 3007
rect 333 3002 338 3003
rect 343 3002 344 3007
rect 1358 3003 1361 3007
rect 1357 3002 1362 3003
rect 1367 3002 1368 3007
rect 2390 3003 2393 3007
rect 2389 3002 2394 3003
rect 2399 3002 2400 3007
rect 2558 3002 2561 3008
rect 3406 3003 3409 3007
rect 3405 3002 3410 3003
rect 3415 3002 3416 3007
rect 4430 3003 4433 3007
rect 4429 3002 4434 3003
rect 4439 3002 4440 3007
rect 5022 2992 5025 2997
rect 1298 2988 1558 2991
rect 1786 2988 2358 2991
rect 2370 2988 2685 2991
rect 2690 2988 3206 2991
rect 4098 2988 4910 2991
rect 1634 2978 1734 2981
rect 1770 2978 1958 2981
rect 2146 2978 2502 2981
rect 2586 2978 3030 2981
rect 3146 2978 4670 2981
rect 5122 2978 5149 2981
rect 1466 2968 1597 2971
rect 1650 2968 2302 2971
rect 2314 2968 2845 2971
rect 2850 2968 2910 2971
rect 3050 2968 3053 2971
rect 3178 2968 3558 2971
rect 5150 2962 5153 2968
rect 1658 2958 1950 2961
rect 1962 2958 2486 2961
rect 2674 2958 3254 2961
rect 4498 2958 4702 2961
rect 4882 2958 4957 2961
rect 4190 2952 4193 2958
rect 678 2948 790 2951
rect 794 2948 1038 2951
rect 1178 2948 1453 2951
rect 678 2942 681 2948
rect 1458 2948 1966 2951
rect 1978 2948 2174 2951
rect 2578 2948 2733 2951
rect 2770 2948 2877 2951
rect 3042 2948 4150 2951
rect 4366 2951 4369 2958
rect 4366 2948 4422 2951
rect 1818 2938 2670 2941
rect 2994 2938 3390 2941
rect 4402 2938 4526 2941
rect 1642 2928 2637 2931
rect 2690 2928 2694 2931
rect 2738 2928 3030 2931
rect 3898 2928 4813 2931
rect 970 2918 1374 2921
rect 1378 2918 2157 2921
rect 2306 2918 3006 2921
rect 3426 2918 3462 2921
rect 4826 2918 4998 2921
rect 1090 2908 1773 2911
rect 1922 2908 2121 2911
rect 2418 2908 2654 2911
rect 4050 2908 4510 2911
rect 4514 2908 4582 2911
rect 854 2903 857 2907
rect 853 2902 858 2903
rect 863 2902 864 2907
rect 1878 2903 1881 2907
rect 1877 2902 1882 2903
rect 1887 2902 1888 2907
rect 1282 2898 1453 2901
rect 1594 2898 1798 2901
rect 2118 2901 2121 2908
rect 2894 2903 2897 2907
rect 2893 2902 2898 2903
rect 2903 2902 2904 2907
rect 3926 2903 3929 2907
rect 3925 2902 3930 2903
rect 3935 2902 3936 2907
rect 4942 2903 4945 2907
rect 4941 2902 4946 2903
rect 4951 2902 4952 2907
rect 5198 2902 5201 2907
rect 2118 2898 2750 2901
rect 458 2888 814 2891
rect 1170 2888 2910 2891
rect 4178 2888 5294 2891
rect 602 2878 1254 2881
rect 1610 2878 1806 2881
rect 2162 2878 3565 2881
rect 4402 2878 4542 2881
rect 4834 2878 4958 2881
rect 714 2868 718 2871
rect 754 2868 806 2871
rect 810 2868 1373 2871
rect 1482 2868 2150 2871
rect 2162 2868 2998 2871
rect 3010 2868 3629 2871
rect 4498 2868 4830 2871
rect 50 2858 262 2861
rect 1290 2858 1558 2861
rect 1634 2858 1741 2861
rect 1778 2858 2317 2861
rect 2610 2858 2662 2861
rect 2946 2858 3966 2861
rect 4290 2858 4534 2861
rect 4602 2858 4822 2861
rect 4886 2861 4889 2868
rect 4826 2858 4889 2861
rect 5202 2858 5206 2861
rect 514 2848 1302 2851
rect 1322 2848 1325 2851
rect 1546 2848 1965 2851
rect 1986 2848 3246 2851
rect 4834 2848 4878 2851
rect 5114 2848 5142 2851
rect 4526 2842 4529 2848
rect 706 2838 1309 2841
rect 1314 2838 1646 2841
rect 1762 2838 2046 2841
rect 2354 2838 2990 2841
rect 3194 2838 4110 2841
rect 5226 2838 5229 2841
rect 1586 2828 2678 2831
rect 2762 2828 2813 2831
rect 2874 2828 2910 2831
rect 2914 2828 3542 2831
rect 3570 2828 4126 2831
rect 5098 2828 5110 2831
rect 5194 2828 5229 2831
rect 362 2818 734 2821
rect 738 2818 2270 2821
rect 2282 2818 3062 2821
rect 3466 2818 3734 2821
rect 5066 2818 5094 2821
rect 1562 2808 2094 2811
rect 2466 2808 2502 2811
rect 2666 2808 2669 2811
rect 2682 2808 3070 2811
rect 5066 2808 5085 2811
rect 5178 2808 5198 2811
rect 334 2803 337 2807
rect 333 2802 338 2803
rect 343 2802 344 2807
rect 1358 2803 1361 2807
rect 1357 2802 1362 2803
rect 1367 2802 1368 2807
rect 2390 2803 2393 2807
rect 2389 2802 2394 2803
rect 2399 2802 2400 2807
rect 3406 2803 3409 2807
rect 3405 2802 3410 2803
rect 3415 2802 3416 2807
rect 4430 2803 4433 2807
rect 4429 2802 4434 2803
rect 4439 2802 4440 2807
rect 786 2798 1102 2801
rect 1378 2798 2334 2801
rect 2406 2798 3110 2801
rect 1042 2788 2198 2791
rect 2406 2791 2409 2798
rect 2322 2788 2409 2791
rect 2302 2782 2305 2787
rect 834 2778 1558 2781
rect 1826 2778 2206 2781
rect 2370 2778 2462 2781
rect 2466 2778 2958 2781
rect 2962 2778 3798 2781
rect 3802 2778 3805 2781
rect 1050 2768 1758 2771
rect 1922 2768 2702 2771
rect 2770 2768 2925 2771
rect 2930 2768 3453 2771
rect 3458 2768 3558 2771
rect 3570 2768 4342 2771
rect 4786 2768 4813 2771
rect 738 2758 942 2761
rect 1682 2758 1990 2761
rect 2186 2758 2301 2761
rect 266 2748 606 2751
rect 718 2751 721 2758
rect 3330 2758 4350 2761
rect 4690 2758 4878 2761
rect 5018 2758 5021 2761
rect 2798 2752 2801 2757
rect 3166 2752 3169 2757
rect 718 2748 974 2751
rect 1714 2748 1725 2751
rect 1762 2748 1902 2751
rect 2026 2748 2798 2751
rect 3290 2748 3494 2751
rect 3498 2748 4078 2751
rect 4910 2751 4913 2758
rect 4282 2748 4913 2751
rect 890 2738 1990 2741
rect 2002 2738 2278 2741
rect 2290 2738 2542 2741
rect 2962 2738 3565 2741
rect 4090 2738 4654 2741
rect 4658 2738 4702 2741
rect 4930 2738 4966 2741
rect 1506 2728 1798 2731
rect 1802 2728 1830 2731
rect 2586 2728 2589 2731
rect 3058 2728 3222 2731
rect 1186 2718 1710 2721
rect 1786 2718 1862 2721
rect 1866 2718 3462 2721
rect 3594 2718 4462 2721
rect 4634 2718 4894 2721
rect 4898 2718 4918 2721
rect 5086 2712 5089 2718
rect 1426 2708 1430 2711
rect 1570 2708 1590 2711
rect 1938 2708 2614 2711
rect 2618 2708 2749 2711
rect 3362 2708 3806 2711
rect 854 2703 857 2707
rect 853 2702 858 2703
rect 863 2702 864 2707
rect 1878 2703 1881 2707
rect 1877 2702 1882 2703
rect 1887 2702 1888 2707
rect 2894 2703 2897 2707
rect 2893 2702 2898 2703
rect 2903 2702 2904 2707
rect 3926 2703 3929 2707
rect 3925 2702 3930 2703
rect 3935 2702 3936 2707
rect 4942 2703 4945 2707
rect 4941 2702 4946 2703
rect 4951 2702 4952 2707
rect 218 2698 310 2701
rect 2050 2698 2073 2701
rect 2186 2698 2189 2701
rect 498 2688 638 2691
rect 1154 2688 2062 2691
rect 2070 2691 2073 2698
rect 2290 2698 2478 2701
rect 2514 2698 2590 2701
rect 3146 2698 3149 2701
rect 4306 2698 4830 2701
rect 5042 2698 5086 2701
rect 2070 2688 2222 2691
rect 2610 2688 2710 2691
rect 2714 2688 3309 2691
rect 3314 2688 3502 2691
rect 3642 2688 3645 2691
rect 3730 2688 4078 2691
rect 4554 2688 4614 2691
rect 5042 2688 5046 2691
rect 530 2678 710 2681
rect 714 2678 1102 2681
rect 1562 2678 1917 2681
rect 2066 2678 2078 2681
rect 2146 2678 2150 2681
rect 2178 2678 2185 2681
rect 2202 2678 2878 2681
rect 3498 2678 3606 2681
rect 4394 2678 4397 2681
rect 2182 2672 2185 2678
rect 4506 2678 4574 2681
rect 4770 2678 4797 2681
rect 90 2668 118 2671
rect 402 2668 550 2671
rect 554 2668 1485 2671
rect 2050 2668 2054 2671
rect 2274 2668 2806 2671
rect 2118 2661 2121 2668
rect 2834 2668 3486 2671
rect 3802 2668 4214 2671
rect 1858 2658 2121 2661
rect 2146 2658 2310 2661
rect 2338 2658 2798 2661
rect 3546 2658 3646 2661
rect 3790 2661 3793 2668
rect 4514 2668 5046 2671
rect 3658 2658 3793 2661
rect 3834 2658 4733 2661
rect 4738 2658 4766 2661
rect 5006 2652 5009 2657
rect 2082 2648 2150 2651
rect 2962 2648 3318 2651
rect 3610 2648 4302 2651
rect 4538 2648 4758 2651
rect 2158 2642 2161 2647
rect 1330 2638 1678 2641
rect 2218 2638 2334 2641
rect 2382 2638 2790 2641
rect 3458 2638 3533 2641
rect 1346 2628 1726 2631
rect 2382 2631 2385 2638
rect 2990 2632 2993 2638
rect 3022 2632 3025 2638
rect 3538 2638 3734 2641
rect 4914 2638 5078 2641
rect 1730 2628 2385 2631
rect 3106 2628 3229 2631
rect 3234 2628 4054 2631
rect 4362 2628 4381 2631
rect 4994 2628 5005 2631
rect 2162 2618 3238 2621
rect 3306 2618 4190 2621
rect 4890 2618 4893 2621
rect 626 2608 1110 2611
rect 2066 2608 2246 2611
rect 2514 2608 3086 2611
rect 3090 2608 3246 2611
rect 3490 2608 3534 2611
rect 3538 2608 4110 2611
rect 334 2603 337 2607
rect 333 2602 338 2603
rect 343 2602 344 2607
rect 1358 2603 1361 2607
rect 1357 2602 1362 2603
rect 1367 2602 1368 2607
rect 2390 2603 2393 2607
rect 2389 2602 2394 2603
rect 2399 2602 2400 2607
rect 3406 2603 3409 2607
rect 3405 2602 3410 2603
rect 3415 2602 3416 2607
rect 4430 2603 4433 2607
rect 4429 2602 4434 2603
rect 4439 2602 4440 2607
rect 762 2598 1341 2601
rect 1450 2598 1934 2601
rect 1970 2598 2198 2601
rect 2626 2598 3094 2601
rect 1330 2588 1686 2591
rect 2186 2588 2534 2591
rect 3074 2588 3558 2591
rect 4058 2588 4614 2591
rect 1266 2578 1526 2581
rect 1586 2578 1758 2581
rect 2642 2578 3062 2581
rect 3906 2578 4286 2581
rect 4490 2578 4493 2581
rect 1122 2568 1462 2571
rect 2106 2568 2118 2571
rect 2250 2568 2422 2571
rect 2570 2568 2637 2571
rect 2762 2568 2990 2571
rect 3650 2568 5190 2571
rect 5250 2568 5286 2571
rect 1906 2558 2086 2561
rect 2178 2558 2398 2561
rect 2906 2558 2982 2561
rect 3082 2558 3406 2561
rect 3410 2558 3417 2561
rect 3778 2558 5246 2561
rect 1242 2548 1830 2551
rect 1842 2548 1918 2551
rect 1946 2548 2438 2551
rect 2570 2548 2573 2551
rect 2826 2548 2950 2551
rect 3010 2548 3030 2551
rect 3802 2548 4134 2551
rect 4474 2548 4494 2551
rect 5106 2548 5118 2551
rect 5242 2548 5245 2551
rect 3102 2542 3105 2548
rect 1346 2538 2206 2541
rect 2218 2538 2558 2541
rect 2866 2538 3086 2541
rect 4282 2538 4430 2541
rect 658 2528 2109 2531
rect 2130 2528 2718 2531
rect 2890 2528 2925 2531
rect 3298 2528 3309 2531
rect 3338 2528 3373 2531
rect 4306 2528 4326 2531
rect 1418 2518 1949 2521
rect 2106 2518 2253 2521
rect 2258 2518 2726 2521
rect 2730 2518 2774 2521
rect 2786 2518 3174 2521
rect 3354 2518 3357 2521
rect 3394 2518 4374 2521
rect 898 2508 934 2511
rect 938 2508 1534 2511
rect 1946 2508 2302 2511
rect 2698 2508 2798 2511
rect 3010 2508 3022 2511
rect 3138 2508 3310 2511
rect 3330 2508 3549 2511
rect 3554 2508 3814 2511
rect 854 2503 857 2507
rect 853 2502 858 2503
rect 863 2502 864 2507
rect 1878 2503 1881 2507
rect 1877 2502 1882 2503
rect 1887 2502 1888 2507
rect 2894 2503 2897 2507
rect 2893 2502 2898 2503
rect 2903 2502 2904 2507
rect 3926 2503 3929 2507
rect 3925 2502 3930 2503
rect 3935 2502 3936 2507
rect 4942 2503 4945 2507
rect 4941 2502 4946 2503
rect 4951 2502 4952 2507
rect 1442 2498 1518 2501
rect 2090 2498 2790 2501
rect 3018 2498 3630 2501
rect 4010 2498 4110 2501
rect 5170 2498 5190 2501
rect 586 2488 813 2491
rect 818 2488 2174 2491
rect 2202 2488 2918 2491
rect 2922 2488 2982 2491
rect 3034 2488 3037 2491
rect 3202 2488 3213 2491
rect 3282 2488 3950 2491
rect 3954 2488 4238 2491
rect 5146 2488 5165 2491
rect 1562 2478 2045 2481
rect 2162 2478 2861 2481
rect 2882 2478 3005 2481
rect 3010 2478 3197 2481
rect 3242 2478 3574 2481
rect 3602 2478 4046 2481
rect 4418 2478 4798 2481
rect 706 2468 854 2471
rect 1506 2468 1878 2471
rect 1906 2468 2054 2471
rect 2450 2468 2662 2471
rect 2762 2468 3046 2471
rect 3186 2468 3326 2471
rect 3346 2468 3470 2471
rect 3738 2468 4038 2471
rect 1570 2458 1574 2461
rect 1634 2458 1926 2461
rect 2018 2458 2022 2461
rect 2126 2461 2129 2468
rect 2114 2458 2129 2461
rect 2146 2458 2366 2461
rect 2378 2458 2477 2461
rect 2522 2458 2525 2461
rect 2562 2458 2766 2461
rect 2786 2458 2929 2461
rect 2938 2458 2974 2461
rect 882 2448 1918 2451
rect 1938 2448 2094 2451
rect 2330 2448 2462 2451
rect 2498 2448 2862 2451
rect 2926 2451 2929 2458
rect 3042 2458 3222 2461
rect 3618 2458 4430 2461
rect 2926 2448 3238 2451
rect 3522 2448 3902 2451
rect 4258 2448 4261 2451
rect 4734 2448 4774 2451
rect 2142 2442 2145 2447
rect 4734 2442 4737 2448
rect 1010 2438 1230 2441
rect 1234 2438 1958 2441
rect 2018 2438 2093 2441
rect 2346 2438 3150 2441
rect 3346 2438 3838 2441
rect 4802 2438 4845 2441
rect 434 2428 974 2431
rect 978 2428 2198 2431
rect 2210 2428 2621 2431
rect 2746 2428 2894 2431
rect 2898 2428 3006 2431
rect 3154 2428 4462 2431
rect 4754 2428 5102 2431
rect 898 2418 1470 2421
rect 1474 2418 1629 2421
rect 2050 2418 2438 2421
rect 2514 2418 2542 2421
rect 2666 2418 3734 2421
rect 4354 2418 4774 2421
rect 906 2408 1342 2411
rect 1842 2408 2205 2411
rect 334 2403 337 2407
rect 333 2402 338 2403
rect 343 2402 344 2407
rect 1358 2403 1361 2407
rect 1357 2402 1362 2403
rect 1367 2402 1368 2407
rect 2390 2403 2393 2407
rect 2389 2402 2394 2403
rect 2399 2402 2400 2407
rect 2558 2402 2561 2417
rect 2706 2408 2726 2411
rect 2842 2408 3037 2411
rect 3066 2408 3334 2411
rect 3490 2408 4070 2411
rect 4074 2408 4230 2411
rect 3406 2403 3409 2407
rect 3405 2402 3410 2403
rect 3415 2402 3416 2407
rect 4430 2403 4433 2407
rect 4429 2402 4434 2403
rect 4439 2402 4440 2407
rect 1394 2398 2054 2401
rect 2698 2398 2966 2401
rect 3106 2398 3190 2401
rect 3202 2398 3393 2401
rect 1458 2388 1670 2391
rect 1834 2388 2361 2391
rect 2370 2388 2829 2391
rect 1586 2378 1846 2381
rect 2074 2378 2262 2381
rect 2358 2381 2361 2388
rect 2978 2388 3078 2391
rect 3390 2391 3393 2398
rect 3390 2388 3582 2391
rect 3618 2388 5286 2391
rect 2358 2378 2654 2381
rect 2674 2378 2694 2381
rect 2802 2378 3197 2381
rect 3330 2378 3446 2381
rect 4922 2378 4925 2381
rect 538 2368 662 2371
rect 746 2368 1638 2371
rect 2058 2368 2521 2371
rect 2530 2368 2790 2371
rect 2818 2368 3037 2371
rect 522 2358 934 2361
rect 1434 2358 1670 2361
rect 1802 2358 2102 2361
rect 2122 2358 2125 2361
rect 2518 2361 2521 2368
rect 3050 2368 3318 2371
rect 3338 2368 3510 2371
rect 3770 2368 3798 2371
rect 3962 2368 4006 2371
rect 2518 2358 2614 2361
rect 2866 2358 3062 2361
rect 3226 2358 3446 2361
rect 3738 2358 4686 2361
rect 5042 2358 5062 2361
rect 554 2348 694 2351
rect 922 2348 1166 2351
rect 1282 2348 1702 2351
rect 1706 2348 1958 2351
rect 1970 2348 2174 2351
rect 2954 2348 3030 2351
rect 3170 2348 3502 2351
rect 3506 2348 3638 2351
rect 458 2338 718 2341
rect 938 2338 1134 2341
rect 1138 2338 1214 2341
rect 1218 2338 1398 2341
rect 1458 2338 1638 2341
rect 1642 2338 1838 2341
rect 1858 2338 1878 2341
rect 2362 2338 2797 2341
rect 2810 2338 2886 2341
rect 3114 2338 3198 2341
rect 3346 2338 3414 2341
rect 3490 2338 3961 2341
rect 1422 2332 1425 2337
rect 1522 2328 1830 2331
rect 1850 2328 2145 2331
rect 2330 2328 3022 2331
rect 1274 2318 1550 2321
rect 1602 2318 1757 2321
rect 1762 2318 1910 2321
rect 2142 2321 2145 2328
rect 3042 2328 3326 2331
rect 3390 2328 3398 2331
rect 3402 2328 3486 2331
rect 3562 2328 3678 2331
rect 3958 2331 3961 2338
rect 3958 2328 5246 2331
rect 2142 2318 2278 2321
rect 2722 2318 3089 2321
rect 3138 2318 3406 2321
rect 3522 2318 5174 2321
rect 5274 2318 5294 2321
rect 1106 2308 1190 2311
rect 2050 2308 2062 2311
rect 2098 2308 2173 2311
rect 2194 2308 2222 2311
rect 2346 2308 2670 2311
rect 3086 2311 3089 2318
rect 3086 2308 3390 2311
rect 854 2303 857 2307
rect 853 2302 858 2303
rect 863 2302 864 2307
rect 1878 2303 1881 2307
rect 1877 2302 1882 2303
rect 1887 2302 1888 2307
rect 2894 2303 2897 2307
rect 2893 2302 2898 2303
rect 2903 2302 2904 2307
rect 3926 2303 3929 2307
rect 3925 2302 3930 2303
rect 3935 2302 3936 2307
rect 4942 2303 4945 2307
rect 4941 2302 4946 2303
rect 4951 2302 4952 2307
rect 1962 2298 2542 2301
rect 2690 2298 2765 2301
rect 2994 2298 3470 2301
rect 818 2288 1374 2291
rect 1490 2288 1606 2291
rect 1866 2288 3214 2291
rect 3226 2288 3438 2291
rect 3442 2288 3550 2291
rect 3554 2288 3614 2291
rect 314 2278 1014 2281
rect 1242 2278 2022 2281
rect 2058 2278 2358 2281
rect 2450 2278 2486 2281
rect 2850 2278 2990 2281
rect 3002 2278 3030 2281
rect 3282 2278 3534 2281
rect 4558 2281 4561 2288
rect 4558 2278 4766 2281
rect 298 2268 374 2271
rect 378 2268 758 2271
rect 802 2268 974 2271
rect 1970 2268 2350 2271
rect 2474 2268 2477 2271
rect 2674 2268 2918 2271
rect 3470 2268 3518 2271
rect 3642 2268 3822 2271
rect 3914 2268 4190 2271
rect 3470 2262 3473 2268
rect 322 2258 990 2261
rect 1186 2258 1246 2261
rect 1818 2258 2126 2261
rect 2258 2258 2406 2261
rect 2458 2258 2646 2261
rect 2658 2258 3134 2261
rect 3234 2258 3382 2261
rect 3554 2258 4238 2261
rect 4242 2258 4478 2261
rect 4698 2258 4717 2261
rect 1302 2251 1305 2258
rect 1058 2248 1305 2251
rect 1638 2248 2669 2251
rect 1638 2241 1641 2248
rect 2690 2248 2710 2251
rect 2730 2248 2742 2251
rect 2746 2248 2822 2251
rect 3210 2248 3678 2251
rect 3846 2248 4449 2251
rect 4586 2248 4606 2251
rect 5090 2248 5142 2251
rect 842 2238 1641 2241
rect 1650 2238 2070 2241
rect 2466 2238 2574 2241
rect 3846 2241 3849 2248
rect 3378 2238 3849 2241
rect 3858 2238 3862 2241
rect 4042 2238 4045 2241
rect 4446 2241 4449 2248
rect 4446 2238 5302 2241
rect 562 2228 1694 2231
rect 1698 2228 1926 2231
rect 1930 2228 1942 2231
rect 2010 2228 2246 2231
rect 2290 2228 2558 2231
rect 3266 2228 3454 2231
rect 5282 2228 5302 2231
rect 1370 2218 1478 2221
rect 1482 2218 1718 2221
rect 1722 2218 1789 2221
rect 2162 2218 2534 2221
rect 1490 2208 1729 2211
rect 2026 2208 2110 2211
rect 2210 2208 2269 2211
rect 334 2203 337 2207
rect 333 2202 338 2203
rect 343 2202 344 2207
rect 1358 2203 1361 2207
rect 1357 2202 1362 2203
rect 1367 2202 1368 2207
rect 1726 2202 1729 2208
rect 2746 2208 3278 2211
rect 4282 2208 4406 2211
rect 2390 2203 2393 2207
rect 2389 2202 2394 2203
rect 2399 2202 2400 2207
rect 3326 2202 3329 2207
rect 3406 2203 3409 2207
rect 3405 2202 3410 2203
rect 3415 2202 3416 2207
rect 4430 2203 4433 2207
rect 4429 2202 4434 2203
rect 4439 2202 4440 2207
rect 1746 2198 2209 2201
rect 2242 2198 2262 2201
rect 2282 2198 2333 2201
rect 2206 2192 2209 2198
rect 2842 2198 3302 2201
rect 666 2188 1462 2191
rect 1590 2181 1593 2188
rect 2306 2188 2374 2191
rect 2514 2188 2550 2191
rect 2578 2188 3277 2191
rect 3306 2188 3342 2191
rect 3346 2188 4078 2191
rect 5114 2188 5126 2191
rect 1338 2178 1593 2181
rect 1602 2178 2342 2181
rect 2490 2178 3726 2181
rect 738 2168 2070 2171
rect 2090 2168 2526 2171
rect 2594 2168 2606 2171
rect 2610 2168 3606 2171
rect 5186 2168 5197 2171
rect 1306 2158 1997 2161
rect 2002 2158 2230 2161
rect 2234 2158 2622 2161
rect 4162 2158 5030 2161
rect 162 2148 950 2151
rect 1170 2148 1542 2151
rect 2298 2148 2317 2151
rect 1226 2138 1534 2141
rect 1934 2141 1937 2148
rect 2774 2148 3286 2151
rect 3370 2148 3894 2151
rect 4330 2148 4654 2151
rect 1650 2138 1937 2141
rect 2774 2141 2777 2148
rect 2298 2138 2777 2141
rect 2786 2138 3334 2141
rect 3738 2138 4174 2141
rect 4178 2138 4382 2141
rect 4386 2138 4638 2141
rect 5182 2132 5185 2138
rect 5218 2138 5254 2141
rect 1010 2128 1486 2131
rect 1706 2128 2374 2131
rect 4042 2128 4758 2131
rect 5218 2128 5238 2131
rect 1042 2118 1686 2121
rect 1714 2118 1718 2121
rect 1862 2118 2270 2121
rect 2366 2118 2478 2121
rect 2530 2118 2758 2121
rect 2914 2118 5246 2121
rect 1862 2111 1865 2118
rect 1194 2108 1865 2111
rect 2366 2111 2369 2118
rect 2074 2108 2369 2111
rect 2378 2108 2670 2111
rect 3010 2108 3078 2111
rect 4146 2108 4342 2111
rect 4418 2108 4918 2111
rect 5186 2108 5229 2111
rect 854 2103 857 2107
rect 853 2102 858 2103
rect 863 2102 864 2107
rect 1878 2103 1881 2107
rect 1877 2102 1882 2103
rect 1887 2102 1888 2107
rect 2894 2103 2897 2107
rect 2893 2102 2898 2103
rect 2903 2102 2904 2107
rect 3926 2103 3929 2107
rect 3925 2102 3930 2103
rect 3935 2102 3936 2107
rect 4942 2103 4945 2107
rect 4941 2102 4946 2103
rect 4951 2102 4952 2107
rect 2194 2098 2230 2101
rect 2930 2098 3846 2101
rect 3850 2098 3885 2101
rect 4306 2098 4622 2101
rect 5226 2098 5245 2101
rect 1770 2088 2589 2091
rect 2594 2088 4318 2091
rect 4330 2088 4534 2091
rect 546 2078 1174 2081
rect 1930 2078 2462 2081
rect 2798 2078 2806 2081
rect 2962 2078 3617 2081
rect 3690 2078 4174 2081
rect 1330 2068 1566 2071
rect 1762 2068 1878 2071
rect 902 2061 905 2068
rect 2146 2068 2166 2071
rect 2798 2071 2801 2078
rect 3614 2072 3617 2078
rect 2226 2068 2801 2071
rect 2810 2068 2973 2071
rect 2986 2068 3414 2071
rect 3418 2068 3518 2071
rect 3562 2068 3598 2071
rect 4154 2068 4157 2071
rect 5234 2068 5281 2071
rect 5278 2062 5281 2068
rect 786 2058 905 2061
rect 1346 2058 1382 2061
rect 1410 2058 1846 2061
rect 1850 2058 1934 2061
rect 2106 2058 2518 2061
rect 3722 2058 3806 2061
rect 4346 2058 4606 2061
rect 4666 2058 4701 2061
rect 4706 2058 4998 2061
rect 3598 2052 3601 2057
rect 514 2048 622 2051
rect 1610 2048 2054 2051
rect 2298 2048 2710 2051
rect 3026 2048 3286 2051
rect 4674 2048 4718 2051
rect 1426 2038 1934 2041
rect 2362 2038 3038 2041
rect 3290 2038 3310 2041
rect 3886 2041 3889 2048
rect 3886 2038 4110 2041
rect 4154 2038 4374 2041
rect 1834 2028 2014 2031
rect 2042 2028 2630 2031
rect 3690 2028 4310 2031
rect 4354 2028 4357 2031
rect 4606 2022 4609 2027
rect 1178 2018 1990 2021
rect 2034 2018 2734 2021
rect 1506 2008 1750 2011
rect 2162 2008 2318 2011
rect 334 2003 337 2007
rect 333 2002 338 2003
rect 343 2002 344 2007
rect 1358 2003 1361 2007
rect 1357 2002 1362 2003
rect 1367 2002 1368 2007
rect 2390 2003 2393 2007
rect 2389 2002 2394 2003
rect 2399 2002 2400 2007
rect 3406 2003 3409 2007
rect 3405 2002 3410 2003
rect 3415 2002 3416 2007
rect 4430 2003 4433 2007
rect 4429 2002 4434 2003
rect 4439 2002 4440 2007
rect 954 1998 957 2001
rect 1786 1998 2214 2001
rect 2650 1998 2678 2001
rect 4050 1998 4230 2001
rect 4458 1998 4622 2001
rect 1234 1988 1726 1991
rect 1842 1988 1854 1991
rect 3282 1988 4214 1991
rect 1866 1978 2118 1981
rect 2266 1978 2478 1981
rect 2482 1978 2806 1981
rect 2810 1978 3078 1981
rect 3210 1978 4190 1981
rect 1782 1971 1785 1978
rect 1466 1968 1785 1971
rect 2162 1968 2798 1971
rect 3010 1968 3430 1971
rect 2846 1962 2849 1967
rect 1426 1958 1702 1961
rect 1730 1958 2254 1961
rect 2266 1958 2742 1961
rect 2962 1958 3414 1961
rect 3418 1958 4246 1961
rect 826 1948 1446 1951
rect 1842 1948 1853 1951
rect 1914 1948 1974 1951
rect 2546 1948 2550 1951
rect 2774 1951 2777 1958
rect 4482 1958 4702 1961
rect 5098 1958 5245 1961
rect 2682 1948 2777 1951
rect 3266 1948 3270 1951
rect 3506 1948 3542 1951
rect 594 1938 654 1941
rect 666 1938 1582 1941
rect 1610 1938 1886 1941
rect 1922 1938 2078 1941
rect 2110 1938 2125 1941
rect 1590 1931 1593 1938
rect 2110 1932 2113 1938
rect 2362 1938 2662 1941
rect 3274 1938 3293 1941
rect 3714 1938 4350 1941
rect 4354 1938 4653 1941
rect 1590 1928 1646 1931
rect 1650 1928 1750 1931
rect 2770 1928 2781 1931
rect 3202 1928 4782 1931
rect 1586 1918 1726 1921
rect 2770 1918 3750 1921
rect 3866 1918 4070 1921
rect 5094 1921 5097 1928
rect 4770 1918 5097 1921
rect 5294 1912 5297 1917
rect 1122 1908 1374 1911
rect 1898 1908 2630 1911
rect 3298 1908 3302 1911
rect 854 1903 857 1907
rect 853 1902 858 1903
rect 863 1902 864 1907
rect 1878 1903 1881 1907
rect 1877 1902 1882 1903
rect 1887 1902 1888 1907
rect 2894 1903 2897 1907
rect 2893 1902 2898 1903
rect 2903 1902 2904 1907
rect 3926 1903 3929 1907
rect 3925 1902 3930 1903
rect 3935 1902 3936 1907
rect 1106 1898 1630 1901
rect 2058 1898 2061 1901
rect 2338 1898 2502 1901
rect 4190 1901 4193 1908
rect 4942 1903 4945 1907
rect 4941 1902 4946 1903
rect 4951 1902 4952 1907
rect 4190 1898 4854 1901
rect 5054 1892 5057 1897
rect 1130 1888 1566 1891
rect 1754 1888 2822 1891
rect 3546 1888 3942 1891
rect 650 1878 1517 1881
rect 1626 1878 2094 1881
rect 2098 1878 2110 1881
rect 2330 1878 2462 1881
rect 2506 1878 2509 1881
rect 2658 1878 3182 1881
rect 3354 1878 3774 1881
rect 4590 1881 4593 1888
rect 4590 1878 5038 1881
rect 5106 1878 5118 1881
rect 850 1868 1142 1871
rect 1150 1868 2038 1871
rect 2082 1868 2454 1871
rect 2522 1868 3150 1871
rect 3546 1868 3630 1871
rect 3666 1868 4046 1871
rect 1150 1861 1153 1868
rect 2062 1862 2065 1868
rect 714 1858 1153 1861
rect 2490 1858 2590 1861
rect 2754 1858 2822 1861
rect 3498 1858 3910 1861
rect 3914 1858 3982 1861
rect 5038 1861 5041 1868
rect 5038 1858 5117 1861
rect 5122 1858 5238 1861
rect 5258 1858 5261 1861
rect 1474 1848 1574 1851
rect 1618 1848 2230 1851
rect 2522 1848 2670 1851
rect 2866 1848 3710 1851
rect 1162 1838 2870 1841
rect 2922 1838 4318 1841
rect 698 1828 2206 1831
rect 2426 1828 3190 1831
rect 3554 1828 4246 1831
rect 34 1818 318 1821
rect 322 1818 782 1821
rect 1530 1818 1950 1821
rect 2570 1818 3110 1821
rect 4178 1818 4557 1821
rect 4562 1818 4678 1821
rect 1378 1808 2070 1811
rect 2634 1808 3030 1811
rect 3858 1808 3950 1811
rect 3954 1808 4414 1811
rect 4594 1808 4958 1811
rect 334 1803 337 1807
rect 333 1802 338 1803
rect 343 1802 344 1807
rect 1358 1803 1361 1807
rect 1357 1802 1362 1803
rect 1367 1802 1368 1807
rect 2390 1803 2393 1807
rect 2389 1802 2394 1803
rect 2399 1802 2400 1807
rect 3406 1803 3409 1807
rect 3405 1802 3410 1803
rect 3415 1802 3416 1807
rect 4430 1803 4433 1807
rect 4429 1802 4434 1803
rect 4439 1802 4440 1807
rect 1386 1798 1814 1801
rect 1970 1798 2174 1801
rect 2666 1798 3382 1801
rect 3674 1798 4414 1801
rect 1918 1792 1921 1797
rect 2074 1788 3166 1791
rect 3170 1788 4222 1791
rect 2034 1778 2038 1781
rect 2122 1778 2566 1781
rect 2714 1778 3654 1781
rect 4498 1778 4502 1781
rect 714 1768 2238 1771
rect 2754 1768 3302 1771
rect 4074 1768 5030 1771
rect 610 1758 758 1761
rect 762 1758 1790 1761
rect 1850 1758 2813 1761
rect 2818 1758 3790 1761
rect 2934 1752 2937 1758
rect 4066 1758 4182 1761
rect 1418 1748 1485 1751
rect 1674 1748 2102 1751
rect 2954 1748 3542 1751
rect 3634 1748 3974 1751
rect 1226 1738 2270 1741
rect 3026 1738 3566 1741
rect 3570 1738 3654 1741
rect 1106 1728 2141 1731
rect 2874 1728 3198 1731
rect 5130 1728 5181 1731
rect 1466 1718 2646 1721
rect 4178 1718 5102 1721
rect 2282 1708 2285 1711
rect 854 1703 857 1707
rect 853 1702 858 1703
rect 863 1702 864 1707
rect 1878 1703 1881 1707
rect 1877 1702 1882 1703
rect 1887 1702 1888 1707
rect 2894 1703 2897 1707
rect 2893 1702 2898 1703
rect 2903 1702 2904 1707
rect 3926 1703 3929 1707
rect 3925 1702 3930 1703
rect 3935 1702 3936 1707
rect 4942 1703 4945 1707
rect 4941 1702 4946 1703
rect 4951 1702 4952 1707
rect 2034 1698 2605 1701
rect 3230 1692 3233 1697
rect 1482 1688 1677 1691
rect 1682 1688 2758 1691
rect 2922 1688 3150 1691
rect 3914 1688 4718 1691
rect 5206 1691 5209 1698
rect 5090 1688 5209 1691
rect 1866 1678 2174 1681
rect 4242 1678 4582 1681
rect 4834 1678 4854 1681
rect 930 1668 1142 1671
rect 1426 1668 1645 1671
rect 2682 1668 3142 1671
rect 3238 1671 3241 1678
rect 3154 1668 3241 1671
rect 4002 1668 4526 1671
rect 2486 1661 2489 1668
rect 2486 1658 2534 1661
rect 2538 1658 2710 1661
rect 3226 1658 3398 1661
rect 4698 1658 4870 1661
rect 1402 1648 1678 1651
rect 2014 1651 2017 1658
rect 2014 1648 2350 1651
rect 2490 1648 2958 1651
rect 3110 1651 3113 1658
rect 3002 1648 3113 1651
rect 3478 1648 4190 1651
rect 1234 1638 1470 1641
rect 1474 1638 2406 1641
rect 3478 1641 3481 1648
rect 2418 1638 3481 1641
rect 3770 1638 4246 1641
rect 5138 1638 5261 1641
rect 1210 1628 1565 1631
rect 1770 1628 2046 1631
rect 2698 1628 4110 1631
rect 1826 1618 2077 1621
rect 2626 1618 3590 1621
rect 2410 1608 2918 1611
rect 3458 1608 4406 1611
rect 334 1603 337 1607
rect 333 1602 338 1603
rect 343 1602 344 1607
rect 1358 1603 1361 1607
rect 1357 1602 1362 1603
rect 1367 1602 1368 1607
rect 2390 1603 2393 1607
rect 2389 1602 2394 1603
rect 2399 1602 2400 1607
rect 3406 1603 3409 1607
rect 3405 1602 3410 1603
rect 3415 1602 3416 1607
rect 4430 1603 4433 1607
rect 4429 1602 4434 1603
rect 4439 1602 4440 1607
rect 1434 1598 2262 1601
rect 2434 1598 3021 1601
rect 3026 1598 3070 1601
rect 1242 1588 2070 1591
rect 2106 1588 2798 1591
rect 2922 1588 3454 1591
rect 3578 1588 4662 1591
rect 458 1578 1062 1581
rect 1418 1578 2157 1581
rect 2170 1578 3278 1581
rect 3538 1578 3542 1581
rect 3906 1578 4382 1581
rect 4402 1578 4814 1581
rect 978 1568 2477 1571
rect 2514 1568 3094 1571
rect 3362 1568 4318 1571
rect 4386 1568 4398 1571
rect 4578 1568 4590 1571
rect 4594 1568 5070 1571
rect 418 1558 1510 1561
rect 1514 1558 1846 1561
rect 2002 1558 2173 1561
rect 2178 1558 3118 1561
rect 3338 1558 3662 1561
rect 3666 1558 3902 1561
rect 4002 1558 4198 1561
rect 4218 1558 4230 1561
rect 4338 1558 4622 1561
rect 634 1548 662 1551
rect 722 1548 1230 1551
rect 1730 1548 1742 1551
rect 2458 1548 2461 1551
rect 2466 1548 3342 1551
rect 3434 1548 3806 1551
rect 3898 1548 4406 1551
rect 4598 1548 4694 1551
rect 3806 1542 3809 1548
rect 4598 1542 4601 1548
rect 410 1538 638 1541
rect 1114 1538 2253 1541
rect 3086 1538 3110 1541
rect 3266 1538 3470 1541
rect 3474 1538 3702 1541
rect 3086 1532 3089 1538
rect 4202 1538 4238 1541
rect 4258 1538 4318 1541
rect 4362 1538 4390 1541
rect 214 1528 598 1531
rect 706 1528 717 1531
rect 214 1522 217 1528
rect 1122 1528 1230 1531
rect 1234 1528 1526 1531
rect 1994 1528 2014 1531
rect 2018 1528 2989 1531
rect 3146 1528 3830 1531
rect 4366 1522 4369 1528
rect 1266 1518 1470 1521
rect 1578 1518 1774 1521
rect 1778 1518 2838 1521
rect 3026 1518 3846 1521
rect 4738 1518 4742 1521
rect 5226 1518 5238 1521
rect 1994 1508 2558 1511
rect 4498 1508 4622 1511
rect 854 1503 857 1507
rect 853 1502 858 1503
rect 863 1502 864 1507
rect 1878 1503 1881 1507
rect 1877 1502 1882 1503
rect 1887 1502 1888 1507
rect 2894 1503 2897 1507
rect 2893 1502 2898 1503
rect 2903 1502 2904 1507
rect 3926 1503 3929 1507
rect 3925 1502 3930 1503
rect 3935 1502 3936 1507
rect 4398 1502 4401 1507
rect 4942 1503 4945 1507
rect 4941 1502 4946 1503
rect 4951 1502 4952 1507
rect 1834 1498 1837 1501
rect 1938 1498 2038 1501
rect 4058 1498 4358 1501
rect 5154 1498 5182 1501
rect 1002 1488 1373 1491
rect 1378 1488 1542 1491
rect 1714 1488 1758 1491
rect 2186 1488 3854 1491
rect 4146 1488 4454 1491
rect 1418 1478 2013 1481
rect 2298 1478 2622 1481
rect 4410 1478 4413 1481
rect 794 1468 1278 1471
rect 1450 1468 1470 1471
rect 1578 1468 1581 1471
rect 1634 1468 1750 1471
rect 1938 1468 2166 1471
rect 2458 1468 3494 1471
rect 410 1458 614 1461
rect 1166 1458 1270 1461
rect 1514 1458 1517 1461
rect 1166 1452 1169 1458
rect 1886 1461 1889 1468
rect 3650 1468 3734 1471
rect 4194 1468 4470 1471
rect 4474 1468 4861 1471
rect 4866 1468 4894 1471
rect 4898 1468 4926 1471
rect 1810 1458 1901 1461
rect 1702 1451 1705 1458
rect 2554 1458 2646 1461
rect 2650 1458 2910 1461
rect 3298 1458 3302 1461
rect 3618 1458 3654 1461
rect 1702 1448 1902 1451
rect 1914 1448 1934 1451
rect 346 1438 686 1441
rect 1730 1438 1894 1441
rect 2006 1441 2009 1448
rect 2322 1448 2998 1451
rect 3106 1448 3118 1451
rect 3258 1448 3974 1451
rect 2006 1438 2270 1441
rect 2410 1438 3053 1441
rect 3290 1438 3742 1441
rect 1522 1428 3438 1431
rect 3802 1428 4374 1431
rect 4994 1428 4998 1431
rect 5042 1428 5110 1431
rect 5138 1428 5158 1431
rect 2274 1418 2550 1421
rect 3066 1418 4525 1421
rect 4530 1418 4534 1421
rect 4570 1418 4806 1421
rect 1834 1408 2310 1411
rect 334 1403 337 1407
rect 333 1402 338 1403
rect 343 1402 344 1407
rect 1358 1403 1361 1407
rect 1357 1402 1362 1403
rect 1367 1402 1368 1407
rect 2390 1403 2393 1407
rect 2389 1402 2394 1403
rect 2399 1402 2400 1407
rect 3406 1403 3409 1407
rect 3405 1402 3410 1403
rect 3415 1402 3416 1407
rect 4430 1403 4433 1407
rect 4429 1402 4434 1403
rect 4439 1402 4440 1407
rect 986 1388 1462 1391
rect 2266 1388 2638 1391
rect 3010 1388 3462 1391
rect 3466 1388 3502 1391
rect 4162 1388 4622 1391
rect 2098 1378 2230 1381
rect 3986 1378 3990 1381
rect 4018 1378 4582 1381
rect 2514 1368 3006 1371
rect 3354 1368 3357 1371
rect 3602 1368 3606 1371
rect 3794 1368 4470 1371
rect 4810 1368 4966 1371
rect 4718 1362 4721 1367
rect 1218 1358 1790 1361
rect 1898 1358 2414 1361
rect 2530 1358 2542 1361
rect 3346 1358 3670 1361
rect 3706 1358 4446 1361
rect 4450 1358 4518 1361
rect 4922 1358 4966 1361
rect 402 1348 422 1351
rect 1610 1348 1710 1351
rect 1762 1348 1782 1351
rect 2234 1348 2509 1351
rect 2522 1348 2798 1351
rect 4210 1348 4214 1351
rect 1498 1338 1766 1341
rect 2074 1338 2401 1341
rect 874 1328 1222 1331
rect 2398 1331 2401 1338
rect 2546 1338 2550 1341
rect 2858 1338 2982 1341
rect 3026 1338 3294 1341
rect 2398 1328 3950 1331
rect 4050 1328 4406 1331
rect 2778 1318 3006 1321
rect 3834 1318 3982 1321
rect 3986 1318 4278 1321
rect 2914 1308 3526 1311
rect 854 1303 857 1307
rect 853 1302 858 1303
rect 863 1302 864 1307
rect 1878 1303 1881 1307
rect 1877 1302 1882 1303
rect 1887 1302 1888 1307
rect 2894 1303 2897 1307
rect 2893 1302 2898 1303
rect 2903 1302 2904 1307
rect 3926 1303 3929 1307
rect 3925 1302 3930 1303
rect 3935 1302 3936 1307
rect 4942 1303 4945 1307
rect 4941 1302 4946 1303
rect 4951 1302 4952 1307
rect 2962 1298 3782 1301
rect 3810 1298 3814 1301
rect 682 1288 798 1291
rect 802 1288 1430 1291
rect 2578 1288 3166 1291
rect 3170 1288 3798 1291
rect 3914 1288 4574 1291
rect 1442 1278 2094 1281
rect 2522 1278 2909 1281
rect 3130 1278 3222 1281
rect 3282 1278 4278 1281
rect 410 1268 854 1271
rect 970 1268 1069 1271
rect 1074 1268 1278 1271
rect 1330 1268 1406 1271
rect 2322 1268 3134 1271
rect 3874 1268 4326 1271
rect 2062 1262 2065 1267
rect 242 1258 958 1261
rect 1674 1258 1870 1261
rect 2490 1258 2534 1261
rect 2962 1258 2990 1261
rect 3302 1258 3582 1261
rect 3586 1258 3790 1261
rect 442 1248 1486 1251
rect 1658 1248 1961 1251
rect 2098 1248 2445 1251
rect 1958 1242 1961 1248
rect 3302 1251 3305 1258
rect 3810 1258 3886 1261
rect 4266 1258 4678 1261
rect 2450 1248 3305 1251
rect 3310 1248 4110 1251
rect 4330 1248 4349 1251
rect 3310 1241 3313 1248
rect 2146 1238 3313 1241
rect 1194 1228 3038 1231
rect 3314 1228 3742 1231
rect 5042 1228 5070 1231
rect 2706 1218 3558 1221
rect 2426 1208 3318 1211
rect 3322 1208 3390 1211
rect 334 1203 337 1207
rect 333 1202 338 1203
rect 343 1202 344 1207
rect 1310 1202 1313 1208
rect 1358 1203 1361 1207
rect 1357 1202 1362 1203
rect 1367 1202 1368 1207
rect 2390 1203 2393 1207
rect 2389 1202 2394 1203
rect 2399 1202 2400 1207
rect 3406 1203 3409 1207
rect 3405 1202 3410 1203
rect 3415 1202 3416 1207
rect 4430 1203 4433 1207
rect 4429 1202 4434 1203
rect 4439 1202 4440 1207
rect 2642 1198 3358 1201
rect 3530 1198 3574 1201
rect 922 1188 1341 1191
rect 1346 1188 2166 1191
rect 2258 1188 2278 1191
rect 3378 1188 4166 1191
rect 4170 1188 4590 1191
rect 2850 1178 3782 1181
rect 5218 1178 5246 1181
rect 4174 1172 4177 1177
rect 570 1168 1014 1171
rect 1018 1168 2686 1171
rect 2730 1168 3014 1171
rect 3170 1168 3726 1171
rect 4650 1168 5190 1171
rect 842 1158 1326 1161
rect 1530 1158 2086 1161
rect 2170 1158 3030 1161
rect 3042 1158 3310 1161
rect 3698 1158 3774 1161
rect 3310 1152 3313 1158
rect 1626 1148 2118 1151
rect 2482 1148 3110 1151
rect 3266 1148 3270 1151
rect 3770 1148 4022 1151
rect 5166 1151 5169 1158
rect 5282 1158 5286 1161
rect 4738 1148 5169 1151
rect 2786 1138 3014 1141
rect 3362 1138 3622 1141
rect 3938 1138 4294 1141
rect 4298 1138 4598 1141
rect 4674 1138 4982 1141
rect 2602 1128 3030 1131
rect 3334 1131 3337 1138
rect 5170 1138 5174 1141
rect 3334 1128 4206 1131
rect 4738 1128 4829 1131
rect 1482 1118 1709 1121
rect 1714 1118 3358 1121
rect 4362 1118 4886 1121
rect 5090 1118 5094 1121
rect 2130 1108 2166 1111
rect 2946 1108 3638 1111
rect 854 1103 857 1107
rect 853 1102 858 1103
rect 863 1102 864 1107
rect 1878 1103 1881 1107
rect 1877 1102 1882 1103
rect 1887 1102 1888 1107
rect 2894 1103 2897 1107
rect 2893 1102 2898 1103
rect 2903 1102 2904 1107
rect 3926 1103 3929 1107
rect 3925 1102 3930 1103
rect 3935 1102 3936 1107
rect 4942 1103 4945 1107
rect 4941 1102 4946 1103
rect 4951 1102 4952 1107
rect 3298 1098 3742 1101
rect 2634 1088 3230 1091
rect 998 1081 1001 1088
rect 998 1078 1134 1081
rect 1138 1078 1638 1081
rect 3154 1078 3782 1081
rect 2674 1068 2726 1071
rect 2994 1068 3878 1071
rect 4930 1068 5158 1071
rect 474 1058 2918 1061
rect 4090 1058 4374 1061
rect 1938 1048 2942 1051
rect 3226 1048 3686 1051
rect 3834 1048 4174 1051
rect 4178 1048 4189 1051
rect 1258 1038 1966 1041
rect 4138 1038 4365 1041
rect 4370 1038 4534 1041
rect 2146 1028 3830 1031
rect 4146 1028 4454 1031
rect 1170 1018 2702 1021
rect 334 1003 337 1007
rect 333 1002 338 1003
rect 343 1002 344 1007
rect 1358 1003 1361 1007
rect 1357 1002 1362 1003
rect 1367 1002 1368 1007
rect 2390 1003 2393 1007
rect 2389 1002 2394 1003
rect 2399 1002 2400 1007
rect 2414 1002 2417 1007
rect 3406 1003 3409 1007
rect 3405 1002 3410 1003
rect 3415 1002 3416 1007
rect 4430 1003 4433 1007
rect 4429 1002 4434 1003
rect 4439 1002 4440 1007
rect 482 988 982 991
rect 1922 988 2790 991
rect 2882 988 4206 991
rect 5274 988 5277 991
rect 594 978 846 981
rect 850 978 1910 981
rect 5130 978 5190 981
rect 5282 978 5293 981
rect 954 968 1662 971
rect 2714 968 3750 971
rect 4010 968 4702 971
rect 814 962 817 967
rect 5070 962 5073 967
rect 1674 958 1821 961
rect 1118 952 1121 958
rect 706 948 1094 951
rect 1174 951 1177 958
rect 1130 948 1177 951
rect 1414 951 1417 958
rect 2266 958 2317 961
rect 2426 958 3222 961
rect 4418 958 4750 961
rect 1414 948 1437 951
rect 1970 948 2294 951
rect 3178 948 4486 951
rect 4490 948 4974 951
rect 322 938 910 941
rect 2710 941 2713 948
rect 1026 938 2713 941
rect 2782 932 2785 938
rect 1098 928 1678 931
rect 1970 918 3142 921
rect 2978 908 3678 911
rect 3682 908 3910 911
rect 854 903 857 907
rect 853 902 858 903
rect 863 902 864 907
rect 1878 903 1881 907
rect 1877 902 1882 903
rect 1887 902 1888 907
rect 2894 903 2897 907
rect 2893 902 2898 903
rect 2903 902 2904 907
rect 3926 903 3929 907
rect 3925 902 3930 903
rect 3935 902 3936 907
rect 4942 903 4945 907
rect 4941 902 4946 903
rect 4951 902 4952 907
rect 2930 898 3822 901
rect 2930 888 3030 891
rect 4626 888 5238 891
rect 946 878 2414 881
rect 618 868 934 871
rect 2322 868 2990 871
rect 3362 868 3414 871
rect 3658 868 4390 871
rect 5182 862 5185 867
rect 586 858 1022 861
rect 1250 858 1613 861
rect 1618 858 1710 861
rect 1714 858 2486 861
rect 3730 858 3862 861
rect 4002 858 4078 861
rect 2990 852 2993 857
rect 1490 848 2478 851
rect 3826 848 4262 851
rect 2378 838 3526 841
rect 3722 838 4174 841
rect 922 818 1246 821
rect 2498 818 3054 821
rect 3642 808 4166 811
rect 334 803 337 807
rect 333 802 338 803
rect 343 802 344 807
rect 1358 803 1361 807
rect 1357 802 1362 803
rect 1367 802 1368 807
rect 2390 803 2393 807
rect 2389 802 2394 803
rect 2399 802 2400 807
rect 3406 803 3409 807
rect 3405 802 3410 803
rect 3415 802 3416 807
rect 4430 803 4433 807
rect 4429 802 4434 803
rect 4439 802 4440 807
rect 1066 788 2310 791
rect 1826 778 4030 781
rect 2322 768 3022 771
rect 4378 768 4622 771
rect 4962 768 5182 771
rect 1226 758 1229 761
rect 998 751 1001 758
rect 3034 758 3149 761
rect 3498 758 3854 761
rect 4690 758 5270 761
rect 998 748 2238 751
rect 4866 748 4990 751
rect 5102 732 5105 737
rect 418 728 934 731
rect 1786 728 1958 731
rect 2978 728 3294 731
rect 58 718 574 721
rect 854 703 857 707
rect 853 702 858 703
rect 863 702 864 707
rect 1878 703 1881 707
rect 1877 702 1882 703
rect 1887 702 1888 707
rect 2894 703 2897 707
rect 2893 702 2898 703
rect 2903 702 2904 707
rect 3926 703 3929 707
rect 3925 702 3930 703
rect 3935 702 3936 707
rect 4942 703 4945 707
rect 4941 702 4946 703
rect 4951 702 4952 707
rect 882 698 1382 701
rect 1962 698 2190 701
rect 874 688 1494 691
rect 3454 682 3457 688
rect 4674 678 4926 681
rect 1374 672 1377 677
rect 5006 672 5009 677
rect 1122 668 1374 671
rect 3626 668 4654 671
rect 1458 658 2358 661
rect 3322 658 4118 661
rect 4122 658 4209 661
rect 4330 658 4886 661
rect 5042 658 5070 661
rect 4206 652 4209 658
rect 2338 648 3062 651
rect 3066 648 3542 651
rect 4090 648 4093 651
rect 4818 648 5182 651
rect 1818 628 3038 631
rect 498 618 1422 621
rect 334 603 337 607
rect 333 602 338 603
rect 343 602 344 607
rect 1358 603 1361 607
rect 1357 602 1362 603
rect 1367 602 1368 607
rect 2390 603 2393 607
rect 2389 602 2394 603
rect 2399 602 2400 607
rect 3406 603 3409 607
rect 3405 602 3410 603
rect 3415 602 3416 607
rect 4430 603 4433 607
rect 4429 602 4434 603
rect 4439 602 4440 607
rect 538 588 1342 591
rect 962 568 1022 571
rect 1026 568 2254 571
rect 2482 568 4205 571
rect 5134 571 5137 578
rect 5026 568 5137 571
rect 346 558 1262 561
rect 1282 558 1798 561
rect 2034 558 2046 561
rect 2050 558 2886 561
rect 3842 558 4886 561
rect 674 548 2093 551
rect 2162 548 2238 551
rect 4562 548 4582 551
rect 210 538 1294 541
rect 1298 538 1782 541
rect 1794 538 2174 541
rect 954 528 3158 531
rect 3642 528 4022 531
rect 854 503 857 507
rect 853 502 858 503
rect 863 502 864 507
rect 1878 503 1881 507
rect 1877 502 1882 503
rect 1887 502 1888 507
rect 2894 503 2897 507
rect 2893 502 2898 503
rect 2903 502 2904 507
rect 3926 503 3929 507
rect 3925 502 3930 503
rect 3935 502 3936 507
rect 4942 503 4945 507
rect 4941 502 4946 503
rect 4951 502 4952 507
rect 1578 488 1934 491
rect 806 478 902 481
rect 906 478 1694 481
rect 1778 478 1894 481
rect 2530 478 4390 481
rect 4842 478 4886 481
rect 4930 478 4990 481
rect 806 472 809 478
rect 3546 468 3974 471
rect 2782 461 2785 468
rect 5202 468 5270 471
rect 2782 458 2870 461
rect 3834 458 4110 461
rect 2706 448 3006 451
rect 3474 448 3534 451
rect 3666 448 4166 451
rect 5230 442 5233 447
rect 1298 438 1965 441
rect 334 403 337 407
rect 333 402 338 403
rect 343 402 344 407
rect 1358 403 1361 407
rect 1357 402 1362 403
rect 1367 402 1368 407
rect 2390 403 2393 407
rect 2389 402 2394 403
rect 2399 402 2400 407
rect 3406 403 3409 407
rect 3405 402 3410 403
rect 3415 402 3416 407
rect 4430 403 4433 407
rect 4429 402 4434 403
rect 4439 402 4440 407
rect 1986 388 3054 391
rect 682 378 1590 381
rect 1594 378 2637 381
rect 818 368 1534 371
rect 1538 368 3662 371
rect 3282 358 3838 361
rect 3842 358 3981 361
rect 338 348 798 351
rect 3202 348 3542 351
rect 994 338 1758 341
rect 5218 318 5286 321
rect 854 303 857 307
rect 853 302 858 303
rect 863 302 864 307
rect 1878 303 1881 307
rect 1877 302 1882 303
rect 1887 302 1888 307
rect 2894 303 2897 307
rect 2893 302 2898 303
rect 2903 302 2904 307
rect 3926 303 3929 307
rect 3925 302 3930 303
rect 3935 302 3936 307
rect 4942 303 4945 307
rect 4941 302 4946 303
rect 4951 302 4952 307
rect 4802 288 5198 291
rect 4002 278 4542 281
rect 4962 278 5022 281
rect 1970 268 1973 271
rect 3490 268 3534 271
rect 5002 268 5037 271
rect 154 258 262 261
rect 3754 258 3998 261
rect 4882 258 5014 261
rect 2034 248 2326 251
rect 334 203 337 207
rect 333 202 338 203
rect 343 202 344 207
rect 1358 203 1361 207
rect 1357 202 1362 203
rect 1367 202 1368 207
rect 2390 203 2393 207
rect 2389 202 2394 203
rect 2399 202 2400 207
rect 3406 203 3409 207
rect 3405 202 3410 203
rect 3415 202 3416 207
rect 4430 203 4433 207
rect 4429 202 4434 203
rect 4439 202 4440 207
rect 5086 192 5089 197
rect 5246 152 5249 158
rect 1786 148 1838 151
rect 2994 148 3078 151
rect 3106 148 3606 151
rect 5282 148 5293 151
rect 3978 138 4062 141
rect 5262 132 5265 138
rect 4434 128 4894 131
rect 4834 118 4973 121
rect 854 103 857 107
rect 853 102 858 103
rect 863 102 864 107
rect 1878 103 1881 107
rect 1877 102 1882 103
rect 1887 102 1888 107
rect 2894 103 2897 107
rect 2893 102 2898 103
rect 2903 102 2904 107
rect 3926 103 3929 107
rect 3925 102 3930 103
rect 3935 102 3936 107
rect 4942 103 4945 107
rect 4941 102 4946 103
rect 4951 102 4952 107
rect 3474 98 3638 101
rect 3490 88 3894 91
rect 4914 88 5149 91
rect 2546 78 3094 81
rect 4674 78 5038 81
rect 2826 68 3430 71
rect 3914 68 4574 71
rect 4826 68 5222 71
rect 2738 58 2910 61
rect 2970 58 3390 61
rect 5138 58 5174 61
rect 334 3 337 7
rect 333 2 338 3
rect 343 2 344 7
rect 1358 3 1361 7
rect 1357 2 1362 3
rect 1367 2 1368 7
rect 2390 3 2393 7
rect 2389 2 2394 3
rect 2399 2 2400 7
rect 3406 3 3409 7
rect 3405 2 3410 3
rect 3415 2 3416 7
rect 4430 3 4433 7
rect 4429 2 4434 3
rect 4439 2 4440 7
<< m6contact >>
rect 848 5103 850 5107
rect 850 5103 853 5107
rect 858 5103 861 5107
rect 861 5103 863 5107
rect 848 5102 853 5103
rect 858 5102 863 5103
rect 1872 5103 1874 5107
rect 1874 5103 1877 5107
rect 1882 5103 1885 5107
rect 1885 5103 1887 5107
rect 1872 5102 1877 5103
rect 1882 5102 1887 5103
rect 2888 5103 2890 5107
rect 2890 5103 2893 5107
rect 2898 5103 2901 5107
rect 2901 5103 2903 5107
rect 2888 5102 2893 5103
rect 2898 5102 2903 5103
rect 3920 5103 3922 5107
rect 3922 5103 3925 5107
rect 3930 5103 3933 5107
rect 3933 5103 3935 5107
rect 3920 5102 3925 5103
rect 3930 5102 3935 5103
rect 4936 5103 4938 5107
rect 4938 5103 4941 5107
rect 4946 5103 4949 5107
rect 4949 5103 4951 5107
rect 4936 5102 4941 5103
rect 4946 5102 4951 5103
rect 4541 5077 4546 5082
rect 4509 5067 4514 5072
rect 4621 5057 4626 5062
rect 4925 5057 4930 5062
rect 4909 5047 4914 5052
rect 4845 5017 4850 5022
rect 328 5003 330 5007
rect 330 5003 333 5007
rect 338 5003 341 5007
rect 341 5003 343 5007
rect 328 5002 333 5003
rect 338 5002 343 5003
rect 1352 5003 1354 5007
rect 1354 5003 1357 5007
rect 1362 5003 1365 5007
rect 1365 5003 1367 5007
rect 1352 5002 1357 5003
rect 1362 5002 1367 5003
rect 2384 5003 2386 5007
rect 2386 5003 2389 5007
rect 2394 5003 2397 5007
rect 2397 5003 2399 5007
rect 2384 5002 2389 5003
rect 2394 5002 2399 5003
rect 3400 5003 3402 5007
rect 3402 5003 3405 5007
rect 3410 5003 3413 5007
rect 3413 5003 3415 5007
rect 3400 5002 3405 5003
rect 3410 5002 3415 5003
rect 4424 5003 4426 5007
rect 4426 5003 4429 5007
rect 4434 5003 4437 5007
rect 4437 5003 4439 5007
rect 4424 5002 4429 5003
rect 4434 5002 4439 5003
rect 5069 4927 5074 4932
rect 848 4903 850 4907
rect 850 4903 853 4907
rect 858 4903 861 4907
rect 861 4903 863 4907
rect 848 4902 853 4903
rect 858 4902 863 4903
rect 1872 4903 1874 4907
rect 1874 4903 1877 4907
rect 1882 4903 1885 4907
rect 1885 4903 1887 4907
rect 1872 4902 1877 4903
rect 1882 4902 1887 4903
rect 2888 4903 2890 4907
rect 2890 4903 2893 4907
rect 2898 4903 2901 4907
rect 2901 4903 2903 4907
rect 2888 4902 2893 4903
rect 2898 4902 2903 4903
rect 3920 4903 3922 4907
rect 3922 4903 3925 4907
rect 3930 4903 3933 4907
rect 3933 4903 3935 4907
rect 3920 4902 3925 4903
rect 3930 4902 3935 4903
rect 4936 4903 4938 4907
rect 4938 4903 4941 4907
rect 4946 4903 4949 4907
rect 4949 4903 4951 4907
rect 4936 4902 4941 4903
rect 4946 4902 4951 4903
rect 5005 4867 5010 4872
rect 4813 4857 4818 4862
rect 5037 4827 5042 4832
rect 328 4803 330 4807
rect 330 4803 333 4807
rect 338 4803 341 4807
rect 341 4803 343 4807
rect 328 4802 333 4803
rect 338 4802 343 4803
rect 1352 4803 1354 4807
rect 1354 4803 1357 4807
rect 1362 4803 1365 4807
rect 1365 4803 1367 4807
rect 1352 4802 1357 4803
rect 1362 4802 1367 4803
rect 2384 4803 2386 4807
rect 2386 4803 2389 4807
rect 2394 4803 2397 4807
rect 2397 4803 2399 4807
rect 2384 4802 2389 4803
rect 2394 4802 2399 4803
rect 3400 4803 3402 4807
rect 3402 4803 3405 4807
rect 3410 4803 3413 4807
rect 3413 4803 3415 4807
rect 3400 4802 3405 4803
rect 3410 4802 3415 4803
rect 4424 4803 4426 4807
rect 4426 4803 4429 4807
rect 4434 4803 4437 4807
rect 4437 4803 4439 4807
rect 4424 4802 4429 4803
rect 4434 4802 4439 4803
rect 5085 4787 5090 4792
rect 4829 4717 4834 4722
rect 848 4703 850 4707
rect 850 4703 853 4707
rect 858 4703 861 4707
rect 861 4703 863 4707
rect 848 4702 853 4703
rect 858 4702 863 4703
rect 1872 4703 1874 4707
rect 1874 4703 1877 4707
rect 1882 4703 1885 4707
rect 1885 4703 1887 4707
rect 1872 4702 1877 4703
rect 1882 4702 1887 4703
rect 2888 4703 2890 4707
rect 2890 4703 2893 4707
rect 2898 4703 2901 4707
rect 2901 4703 2903 4707
rect 2888 4702 2893 4703
rect 2898 4702 2903 4703
rect 3920 4703 3922 4707
rect 3922 4703 3925 4707
rect 3930 4703 3933 4707
rect 3933 4703 3935 4707
rect 3920 4702 3925 4703
rect 3930 4702 3935 4703
rect 4936 4703 4938 4707
rect 4938 4703 4941 4707
rect 4946 4703 4949 4707
rect 4949 4703 4951 4707
rect 4936 4702 4941 4703
rect 4946 4702 4951 4703
rect 5245 4697 5250 4702
rect 5133 4637 5138 4642
rect 328 4603 330 4607
rect 330 4603 333 4607
rect 338 4603 341 4607
rect 341 4603 343 4607
rect 328 4602 333 4603
rect 338 4602 343 4603
rect 1352 4603 1354 4607
rect 1354 4603 1357 4607
rect 1362 4603 1365 4607
rect 1365 4603 1367 4607
rect 1352 4602 1357 4603
rect 1362 4602 1367 4603
rect 2384 4603 2386 4607
rect 2386 4603 2389 4607
rect 2394 4603 2397 4607
rect 2397 4603 2399 4607
rect 2384 4602 2389 4603
rect 2394 4602 2399 4603
rect 3400 4603 3402 4607
rect 3402 4603 3405 4607
rect 3410 4603 3413 4607
rect 3413 4603 3415 4607
rect 3400 4602 3405 4603
rect 3410 4602 3415 4603
rect 4424 4603 4426 4607
rect 4426 4603 4429 4607
rect 4434 4603 4437 4607
rect 4437 4603 4439 4607
rect 4424 4602 4429 4603
rect 4434 4602 4439 4603
rect 5021 4587 5026 4592
rect 4973 4557 4978 4562
rect 4989 4537 4994 4542
rect 5165 4537 5170 4542
rect 848 4503 850 4507
rect 850 4503 853 4507
rect 858 4503 861 4507
rect 861 4503 863 4507
rect 848 4502 853 4503
rect 858 4502 863 4503
rect 1872 4503 1874 4507
rect 1874 4503 1877 4507
rect 1882 4503 1885 4507
rect 1885 4503 1887 4507
rect 1872 4502 1877 4503
rect 1882 4502 1887 4503
rect 2888 4503 2890 4507
rect 2890 4503 2893 4507
rect 2898 4503 2901 4507
rect 2901 4503 2903 4507
rect 2888 4502 2893 4503
rect 2898 4502 2903 4503
rect 3920 4503 3922 4507
rect 3922 4503 3925 4507
rect 3930 4503 3933 4507
rect 3933 4503 3935 4507
rect 3920 4502 3925 4503
rect 3930 4502 3935 4503
rect 4936 4503 4938 4507
rect 4938 4503 4941 4507
rect 4946 4503 4949 4507
rect 4949 4503 4951 4507
rect 4936 4502 4941 4503
rect 4946 4502 4951 4503
rect 4957 4467 4962 4472
rect 2061 4457 2066 4462
rect 2749 4457 2754 4462
rect 5197 4457 5202 4462
rect 328 4403 330 4407
rect 330 4403 333 4407
rect 338 4403 341 4407
rect 341 4403 343 4407
rect 328 4402 333 4403
rect 338 4402 343 4403
rect 1352 4403 1354 4407
rect 1354 4403 1357 4407
rect 1362 4403 1365 4407
rect 1365 4403 1367 4407
rect 1352 4402 1357 4403
rect 1362 4402 1367 4403
rect 2384 4403 2386 4407
rect 2386 4403 2389 4407
rect 2394 4403 2397 4407
rect 2397 4403 2399 4407
rect 2384 4402 2389 4403
rect 2394 4402 2399 4403
rect 3400 4403 3402 4407
rect 3402 4403 3405 4407
rect 3410 4403 3413 4407
rect 3413 4403 3415 4407
rect 3400 4402 3405 4403
rect 3410 4402 3415 4403
rect 4424 4403 4426 4407
rect 4426 4403 4429 4407
rect 4434 4403 4437 4407
rect 4437 4403 4439 4407
rect 4424 4402 4429 4403
rect 4434 4402 4439 4403
rect 1453 4357 1458 4362
rect 4093 4357 4098 4362
rect 4861 4337 4866 4342
rect 5277 4307 5282 4312
rect 848 4303 850 4307
rect 850 4303 853 4307
rect 858 4303 861 4307
rect 861 4303 863 4307
rect 848 4302 853 4303
rect 858 4302 863 4303
rect 1872 4303 1874 4307
rect 1874 4303 1877 4307
rect 1882 4303 1885 4307
rect 1885 4303 1887 4307
rect 1872 4302 1877 4303
rect 1882 4302 1887 4303
rect 2888 4303 2890 4307
rect 2890 4303 2893 4307
rect 2898 4303 2901 4307
rect 2901 4303 2903 4307
rect 2888 4302 2893 4303
rect 2898 4302 2903 4303
rect 3920 4303 3922 4307
rect 3922 4303 3925 4307
rect 3930 4303 3933 4307
rect 3933 4303 3935 4307
rect 3920 4302 3925 4303
rect 3930 4302 3935 4303
rect 4936 4303 4938 4307
rect 4938 4303 4941 4307
rect 4946 4303 4949 4307
rect 4949 4303 4951 4307
rect 4936 4302 4941 4303
rect 4946 4302 4951 4303
rect 2077 4287 2082 4292
rect 5101 4287 5106 4292
rect 1685 4267 1690 4272
rect 5053 4267 5058 4272
rect 2573 4257 2578 4262
rect 3549 4247 3554 4252
rect 4653 4247 4658 4252
rect 328 4203 330 4207
rect 330 4203 333 4207
rect 338 4203 341 4207
rect 341 4203 343 4207
rect 328 4202 333 4203
rect 338 4202 343 4203
rect 1352 4203 1354 4207
rect 1354 4203 1357 4207
rect 1362 4203 1365 4207
rect 1365 4203 1367 4207
rect 1352 4202 1357 4203
rect 1362 4202 1367 4203
rect 2384 4203 2386 4207
rect 2386 4203 2389 4207
rect 2394 4203 2397 4207
rect 2397 4203 2399 4207
rect 2384 4202 2389 4203
rect 2394 4202 2399 4203
rect 3400 4203 3402 4207
rect 3402 4203 3405 4207
rect 3410 4203 3413 4207
rect 3413 4203 3415 4207
rect 3400 4202 3405 4203
rect 3410 4202 3415 4203
rect 4424 4203 4426 4207
rect 4426 4203 4429 4207
rect 4434 4203 4437 4207
rect 4437 4203 4439 4207
rect 4424 4202 4429 4203
rect 4434 4202 4439 4203
rect 4653 4167 4658 4172
rect 3037 4157 3042 4162
rect 4525 4127 4530 4132
rect 5213 4117 5218 4122
rect 3037 4107 3042 4112
rect 848 4103 850 4107
rect 850 4103 853 4107
rect 858 4103 861 4107
rect 861 4103 863 4107
rect 848 4102 853 4103
rect 858 4102 863 4103
rect 1872 4103 1874 4107
rect 1874 4103 1877 4107
rect 1882 4103 1885 4107
rect 1885 4103 1887 4107
rect 1872 4102 1877 4103
rect 1882 4102 1887 4103
rect 2888 4103 2890 4107
rect 2890 4103 2893 4107
rect 2898 4103 2901 4107
rect 2901 4103 2903 4107
rect 2888 4102 2893 4103
rect 2898 4102 2903 4103
rect 3920 4103 3922 4107
rect 3922 4103 3925 4107
rect 3930 4103 3933 4107
rect 3933 4103 3935 4107
rect 3920 4102 3925 4103
rect 3930 4102 3935 4103
rect 4936 4103 4938 4107
rect 4938 4103 4941 4107
rect 4946 4103 4949 4107
rect 4949 4103 4951 4107
rect 4936 4102 4941 4103
rect 4946 4102 4951 4103
rect 5261 4077 5266 4082
rect 1597 4057 1602 4062
rect 4589 4017 4594 4022
rect 328 4003 330 4007
rect 330 4003 333 4007
rect 338 4003 341 4007
rect 341 4003 343 4007
rect 328 4002 333 4003
rect 338 4002 343 4003
rect 1352 4003 1354 4007
rect 1354 4003 1357 4007
rect 1362 4003 1365 4007
rect 1365 4003 1367 4007
rect 1352 4002 1357 4003
rect 1362 4002 1367 4003
rect 2384 4003 2386 4007
rect 2386 4003 2389 4007
rect 2394 4003 2397 4007
rect 2397 4003 2399 4007
rect 2384 4002 2389 4003
rect 2394 4002 2399 4003
rect 3261 4007 3266 4012
rect 3400 4003 3402 4007
rect 3402 4003 3405 4007
rect 3410 4003 3413 4007
rect 3413 4003 3415 4007
rect 3400 4002 3405 4003
rect 3410 4002 3415 4003
rect 4424 4003 4426 4007
rect 4426 4003 4429 4007
rect 4434 4003 4437 4007
rect 4437 4003 4439 4007
rect 4424 4002 4429 4003
rect 4434 4002 4439 4003
rect 1469 3997 1474 4002
rect 2685 3997 2690 4002
rect 5117 3997 5122 4002
rect 5149 3997 5154 4002
rect 4493 3978 4494 3982
rect 4494 3978 4498 3982
rect 4493 3977 4498 3978
rect 5021 3967 5026 3972
rect 4685 3957 4690 3962
rect 3485 3937 3490 3942
rect 5037 3937 5042 3942
rect 5149 3927 5154 3932
rect 848 3903 850 3907
rect 850 3903 853 3907
rect 858 3903 861 3907
rect 861 3903 863 3907
rect 848 3902 853 3903
rect 858 3902 863 3903
rect 1872 3903 1874 3907
rect 1874 3903 1877 3907
rect 1882 3903 1885 3907
rect 1885 3903 1887 3907
rect 1872 3902 1877 3903
rect 1882 3902 1887 3903
rect 2888 3903 2890 3907
rect 2890 3903 2893 3907
rect 2898 3903 2901 3907
rect 2901 3903 2903 3907
rect 2888 3902 2893 3903
rect 2898 3902 2903 3903
rect 3920 3903 3922 3907
rect 3922 3903 3925 3907
rect 3930 3903 3933 3907
rect 3933 3903 3935 3907
rect 3920 3902 3925 3903
rect 3930 3902 3935 3903
rect 4936 3903 4938 3907
rect 4938 3903 4941 3907
rect 4946 3903 4949 3907
rect 4949 3903 4951 3907
rect 4936 3902 4941 3903
rect 4946 3902 4951 3903
rect 1997 3867 2002 3872
rect 5181 3867 5186 3872
rect 1965 3857 1970 3862
rect 5229 3857 5234 3862
rect 2973 3847 2978 3852
rect 4989 3847 4994 3852
rect 4973 3837 4978 3842
rect 4989 3837 4994 3842
rect 3197 3827 3202 3832
rect 328 3803 330 3807
rect 330 3803 333 3807
rect 338 3803 341 3807
rect 341 3803 343 3807
rect 328 3802 333 3803
rect 338 3802 343 3803
rect 1352 3803 1354 3807
rect 1354 3803 1357 3807
rect 1362 3803 1365 3807
rect 1365 3803 1367 3807
rect 1352 3802 1357 3803
rect 1362 3802 1367 3803
rect 2384 3803 2386 3807
rect 2386 3803 2389 3807
rect 2394 3803 2397 3807
rect 2397 3803 2399 3807
rect 2384 3802 2389 3803
rect 2394 3802 2399 3803
rect 3400 3803 3402 3807
rect 3402 3803 3405 3807
rect 3410 3803 3413 3807
rect 3413 3803 3415 3807
rect 3400 3802 3405 3803
rect 3410 3802 3415 3803
rect 4424 3803 4426 3807
rect 4426 3803 4429 3807
rect 4434 3803 4437 3807
rect 4437 3803 4439 3807
rect 4424 3802 4429 3803
rect 4434 3802 4439 3803
rect 2925 3777 2930 3782
rect 4701 3757 4706 3762
rect 1613 3737 1618 3742
rect 2877 3727 2882 3732
rect 2173 3717 2178 3722
rect 5005 3717 5010 3722
rect 5149 3717 5154 3722
rect 1069 3707 1074 3712
rect 5133 3707 5138 3712
rect 848 3703 850 3707
rect 850 3703 853 3707
rect 858 3703 861 3707
rect 861 3703 863 3707
rect 848 3702 853 3703
rect 858 3702 863 3703
rect 1872 3703 1874 3707
rect 1874 3703 1877 3707
rect 1882 3703 1885 3707
rect 1885 3703 1887 3707
rect 1872 3702 1877 3703
rect 1882 3702 1887 3703
rect 2888 3703 2890 3707
rect 2890 3703 2893 3707
rect 2898 3703 2901 3707
rect 2901 3703 2903 3707
rect 2888 3702 2893 3703
rect 2898 3702 2903 3703
rect 3920 3703 3922 3707
rect 3922 3703 3925 3707
rect 3930 3703 3933 3707
rect 3933 3703 3935 3707
rect 3920 3702 3925 3703
rect 3930 3702 3935 3703
rect 4936 3703 4938 3707
rect 4938 3703 4941 3707
rect 4946 3703 4949 3707
rect 4949 3703 4951 3707
rect 4936 3702 4941 3703
rect 4946 3702 4951 3703
rect 2701 3697 2706 3702
rect 5037 3697 5042 3702
rect 3901 3687 3906 3692
rect 5005 3687 5010 3692
rect 5133 3687 5138 3692
rect 5165 3687 5170 3692
rect 4973 3677 4978 3682
rect 3309 3667 3314 3672
rect 3901 3667 3906 3672
rect 1741 3647 1746 3652
rect 1797 3647 1802 3652
rect 2797 3647 2802 3652
rect 3165 3647 3170 3652
rect 1117 3637 1122 3642
rect 4669 3637 4674 3642
rect 2109 3627 2114 3632
rect 4157 3617 4162 3622
rect 328 3603 330 3607
rect 330 3603 333 3607
rect 338 3603 341 3607
rect 341 3603 343 3607
rect 328 3602 333 3603
rect 338 3602 343 3603
rect 1352 3603 1354 3607
rect 1354 3603 1357 3607
rect 1362 3603 1365 3607
rect 1365 3603 1367 3607
rect 1352 3602 1357 3603
rect 1362 3602 1367 3603
rect 2384 3603 2386 3607
rect 2386 3603 2389 3607
rect 2394 3603 2397 3607
rect 2397 3603 2399 3607
rect 2384 3602 2389 3603
rect 2394 3602 2399 3603
rect 3400 3603 3402 3607
rect 3402 3603 3405 3607
rect 3410 3603 3413 3607
rect 3413 3603 3415 3607
rect 3400 3602 3405 3603
rect 3410 3602 3415 3603
rect 4424 3603 4426 3607
rect 4426 3603 4429 3607
rect 4434 3603 4437 3607
rect 4437 3603 4439 3607
rect 4424 3602 4429 3603
rect 4434 3602 4439 3603
rect 1485 3597 1490 3602
rect 2253 3587 2258 3592
rect 1645 3567 1650 3572
rect 2253 3567 2258 3572
rect 1741 3557 1746 3562
rect 5101 3557 5106 3562
rect 5165 3557 5170 3562
rect 3213 3537 3218 3542
rect 3101 3527 3106 3532
rect 2477 3507 2482 3512
rect 848 3503 850 3507
rect 850 3503 853 3507
rect 858 3503 861 3507
rect 861 3503 863 3507
rect 848 3502 853 3503
rect 858 3502 863 3503
rect 1872 3503 1874 3507
rect 1874 3503 1877 3507
rect 1882 3503 1885 3507
rect 1885 3503 1887 3507
rect 1872 3502 1877 3503
rect 1882 3502 1887 3503
rect 2888 3503 2890 3507
rect 2890 3503 2893 3507
rect 2898 3503 2901 3507
rect 2901 3503 2903 3507
rect 2888 3502 2893 3503
rect 2898 3502 2903 3503
rect 3920 3503 3922 3507
rect 3922 3503 3925 3507
rect 3930 3503 3933 3507
rect 3933 3503 3935 3507
rect 3920 3502 3925 3503
rect 3930 3502 3935 3503
rect 5021 3507 5026 3512
rect 4936 3503 4938 3507
rect 4938 3503 4941 3507
rect 4946 3503 4949 3507
rect 4949 3503 4951 3507
rect 4936 3502 4941 3503
rect 4946 3502 4951 3503
rect 1901 3497 1906 3502
rect 4877 3497 4882 3502
rect 2301 3487 2306 3492
rect 4173 3467 4178 3472
rect 4765 3467 4770 3472
rect 1325 3447 1330 3452
rect 3309 3447 3314 3452
rect 4205 3417 4210 3422
rect 328 3403 330 3407
rect 330 3403 333 3407
rect 338 3403 341 3407
rect 341 3403 343 3407
rect 328 3402 333 3403
rect 338 3402 343 3403
rect 1352 3403 1354 3407
rect 1354 3403 1357 3407
rect 1362 3403 1365 3407
rect 1365 3403 1367 3407
rect 1352 3402 1357 3403
rect 1362 3402 1367 3403
rect 2384 3403 2386 3407
rect 2386 3403 2389 3407
rect 2394 3403 2397 3407
rect 2397 3403 2399 3407
rect 2384 3402 2389 3403
rect 2394 3402 2399 3403
rect 3400 3403 3402 3407
rect 3402 3403 3405 3407
rect 3410 3403 3413 3407
rect 3413 3403 3415 3407
rect 3400 3402 3405 3403
rect 3410 3402 3415 3403
rect 4424 3403 4426 3407
rect 4426 3403 4429 3407
rect 4434 3403 4437 3407
rect 4437 3403 4439 3407
rect 4424 3402 4429 3403
rect 4434 3402 4439 3403
rect 4989 3387 4994 3392
rect 3997 3377 4002 3382
rect 4989 3367 4994 3372
rect 2925 3347 2930 3352
rect 1645 3327 1650 3332
rect 4573 3327 4578 3332
rect 2333 3307 2338 3312
rect 848 3303 850 3307
rect 850 3303 853 3307
rect 858 3303 861 3307
rect 861 3303 863 3307
rect 848 3302 853 3303
rect 858 3302 863 3303
rect 1872 3303 1874 3307
rect 1874 3303 1877 3307
rect 1882 3303 1885 3307
rect 1885 3303 1887 3307
rect 1872 3302 1877 3303
rect 1882 3302 1887 3303
rect 2888 3303 2890 3307
rect 2890 3303 2893 3307
rect 2898 3303 2901 3307
rect 2901 3303 2903 3307
rect 2888 3302 2893 3303
rect 2898 3302 2903 3303
rect 3920 3303 3922 3307
rect 3922 3303 3925 3307
rect 3930 3303 3933 3307
rect 3933 3303 3935 3307
rect 3920 3302 3925 3303
rect 3930 3302 3935 3303
rect 4936 3303 4938 3307
rect 4938 3303 4941 3307
rect 4946 3303 4949 3307
rect 4949 3303 4951 3307
rect 4936 3302 4941 3303
rect 4946 3302 4951 3303
rect 2877 3287 2882 3292
rect 4477 3287 4482 3292
rect 3293 3277 3298 3282
rect 2413 3267 2418 3272
rect 2781 3257 2786 3262
rect 5293 3257 5298 3262
rect 4605 3227 4610 3232
rect 3885 3217 3890 3222
rect 5101 3207 5106 3212
rect 328 3203 330 3207
rect 330 3203 333 3207
rect 338 3203 341 3207
rect 341 3203 343 3207
rect 328 3202 333 3203
rect 338 3202 343 3203
rect 1352 3203 1354 3207
rect 1354 3203 1357 3207
rect 1362 3203 1365 3207
rect 1365 3203 1367 3207
rect 1352 3202 1357 3203
rect 1362 3202 1367 3203
rect 2384 3203 2386 3207
rect 2386 3203 2389 3207
rect 2394 3203 2397 3207
rect 2397 3203 2399 3207
rect 2384 3202 2389 3203
rect 2394 3202 2399 3203
rect 3400 3203 3402 3207
rect 3402 3203 3405 3207
rect 3410 3203 3413 3207
rect 3413 3203 3415 3207
rect 3400 3202 3405 3203
rect 3410 3202 3415 3203
rect 4424 3203 4426 3207
rect 4426 3203 4429 3207
rect 4434 3203 4437 3207
rect 4437 3203 4439 3207
rect 4424 3202 4429 3203
rect 4434 3202 4439 3203
rect 4957 3187 4962 3192
rect 5213 3187 5218 3192
rect 5037 3177 5042 3182
rect 5037 3167 5042 3172
rect 5213 3167 5218 3172
rect 2109 3147 2114 3152
rect 5277 3157 5282 3162
rect 3037 3147 3042 3152
rect 4541 3147 4546 3152
rect 3037 3127 3042 3132
rect 4413 3127 4418 3132
rect 5277 3127 5282 3132
rect 2493 3117 2498 3122
rect 848 3103 850 3107
rect 850 3103 853 3107
rect 858 3103 861 3107
rect 861 3103 863 3107
rect 848 3102 853 3103
rect 858 3102 863 3103
rect 1872 3103 1874 3107
rect 1874 3103 1877 3107
rect 1882 3103 1885 3107
rect 1885 3103 1887 3107
rect 1872 3102 1877 3103
rect 1882 3102 1887 3103
rect 2888 3103 2890 3107
rect 2890 3103 2893 3107
rect 2898 3103 2901 3107
rect 2901 3103 2903 3107
rect 2888 3102 2893 3103
rect 2898 3102 2903 3103
rect 3920 3103 3922 3107
rect 3922 3103 3925 3107
rect 3930 3103 3933 3107
rect 3933 3103 3935 3107
rect 3920 3102 3925 3103
rect 3930 3102 3935 3103
rect 4936 3103 4938 3107
rect 4938 3103 4941 3107
rect 4946 3103 4949 3107
rect 4949 3103 4951 3107
rect 4936 3102 4941 3103
rect 4946 3102 4951 3103
rect 2349 3077 2354 3082
rect 4893 3087 4898 3092
rect 1949 3057 1954 3062
rect 2669 3057 2674 3062
rect 1917 3047 1922 3052
rect 4061 3047 4066 3052
rect 2125 3027 2130 3032
rect 2493 3027 2498 3032
rect 2669 3017 2674 3022
rect 1517 3007 1522 3012
rect 328 3003 330 3007
rect 330 3003 333 3007
rect 338 3003 341 3007
rect 341 3003 343 3007
rect 328 3002 333 3003
rect 338 3002 343 3003
rect 1352 3003 1354 3007
rect 1354 3003 1357 3007
rect 1362 3003 1365 3007
rect 1365 3003 1367 3007
rect 1352 3002 1357 3003
rect 1362 3002 1367 3003
rect 2384 3003 2386 3007
rect 2386 3003 2389 3007
rect 2394 3003 2397 3007
rect 2397 3003 2399 3007
rect 2384 3002 2389 3003
rect 2394 3002 2399 3003
rect 3341 3007 3346 3012
rect 3400 3003 3402 3007
rect 3402 3003 3405 3007
rect 3410 3003 3413 3007
rect 3413 3003 3415 3007
rect 3400 3002 3405 3003
rect 3410 3002 3415 3003
rect 4424 3003 4426 3007
rect 4426 3003 4429 3007
rect 4434 3003 4437 3007
rect 4437 3003 4439 3007
rect 4424 3002 4429 3003
rect 4434 3002 4439 3003
rect 2557 2997 2562 3002
rect 5021 2997 5026 3002
rect 2685 2987 2690 2992
rect 5149 2977 5154 2982
rect 1597 2967 1602 2972
rect 2845 2967 2850 2972
rect 3053 2967 3058 2972
rect 1453 2947 1458 2952
rect 2733 2947 2738 2952
rect 2877 2947 2882 2952
rect 4189 2947 4194 2952
rect 4957 2957 4962 2962
rect 5149 2957 5154 2962
rect 2637 2927 2642 2932
rect 2685 2927 2690 2932
rect 2733 2927 2738 2932
rect 4813 2927 4818 2932
rect 2157 2917 2162 2922
rect 1773 2907 1778 2912
rect 848 2903 850 2907
rect 850 2903 853 2907
rect 858 2903 861 2907
rect 861 2903 863 2907
rect 848 2902 853 2903
rect 858 2902 863 2903
rect 1872 2903 1874 2907
rect 1874 2903 1877 2907
rect 1882 2903 1885 2907
rect 1885 2903 1887 2907
rect 1872 2902 1877 2903
rect 1882 2902 1887 2903
rect 1453 2897 1458 2902
rect 5197 2907 5202 2912
rect 2888 2903 2890 2907
rect 2890 2903 2893 2907
rect 2898 2903 2901 2907
rect 2901 2903 2903 2907
rect 2888 2902 2893 2903
rect 2898 2902 2903 2903
rect 3920 2903 3922 2907
rect 3922 2903 3925 2907
rect 3930 2903 3933 2907
rect 3933 2903 3935 2907
rect 3920 2902 3925 2903
rect 3930 2902 3935 2903
rect 4936 2903 4938 2907
rect 4938 2903 4941 2907
rect 4946 2903 4949 2907
rect 4949 2903 4951 2907
rect 4936 2902 4941 2903
rect 4946 2902 4951 2903
rect 3565 2877 3570 2882
rect 709 2867 714 2872
rect 1373 2867 1378 2872
rect 2157 2867 2162 2872
rect 3629 2867 3634 2872
rect 4493 2867 4498 2872
rect 1741 2857 1746 2862
rect 1773 2857 1778 2862
rect 2317 2857 2322 2862
rect 5197 2857 5202 2862
rect 1325 2847 1330 2852
rect 1965 2847 1970 2852
rect 1309 2837 1314 2842
rect 2349 2837 2354 2842
rect 4525 2837 4530 2842
rect 5229 2837 5234 2842
rect 2813 2827 2818 2832
rect 3565 2828 3566 2832
rect 3566 2828 3570 2832
rect 3565 2827 3570 2828
rect 5229 2827 5234 2832
rect 2461 2807 2466 2812
rect 2669 2807 2674 2812
rect 5085 2807 5090 2812
rect 328 2803 330 2807
rect 330 2803 333 2807
rect 338 2803 341 2807
rect 341 2803 343 2807
rect 328 2802 333 2803
rect 338 2802 343 2803
rect 1352 2803 1354 2807
rect 1354 2803 1357 2807
rect 1362 2803 1365 2807
rect 1365 2803 1367 2807
rect 1352 2802 1357 2803
rect 1362 2802 1367 2803
rect 2384 2803 2386 2807
rect 2386 2803 2389 2807
rect 2394 2803 2397 2807
rect 2397 2803 2399 2807
rect 2384 2802 2389 2803
rect 2394 2802 2399 2803
rect 3400 2803 3402 2807
rect 3402 2803 3405 2807
rect 3410 2803 3413 2807
rect 3413 2803 3415 2807
rect 3400 2802 3405 2803
rect 3410 2802 3415 2803
rect 4424 2803 4426 2807
rect 4426 2803 4429 2807
rect 4434 2803 4437 2807
rect 4437 2803 4439 2807
rect 4424 2802 4429 2803
rect 4434 2802 4439 2803
rect 1373 2797 1378 2802
rect 2301 2787 2306 2792
rect 2317 2787 2322 2792
rect 1821 2777 1826 2782
rect 3805 2777 3810 2782
rect 2765 2767 2770 2772
rect 2925 2767 2930 2772
rect 3453 2767 3458 2772
rect 3565 2767 3570 2772
rect 4813 2767 4818 2772
rect 2301 2757 2306 2762
rect 2797 2757 2802 2762
rect 3165 2757 3170 2762
rect 1725 2747 1730 2752
rect 5021 2757 5026 2762
rect 2285 2737 2290 2742
rect 3565 2737 3570 2742
rect 4925 2737 4930 2742
rect 2589 2727 2594 2732
rect 1421 2707 1426 2712
rect 2749 2707 2754 2712
rect 5085 2707 5090 2712
rect 848 2703 850 2707
rect 850 2703 853 2707
rect 858 2703 861 2707
rect 861 2703 863 2707
rect 848 2702 853 2703
rect 858 2702 863 2703
rect 1872 2703 1874 2707
rect 1874 2703 1877 2707
rect 1882 2703 1885 2707
rect 1885 2703 1887 2707
rect 1872 2702 1877 2703
rect 1882 2702 1887 2703
rect 2888 2703 2890 2707
rect 2890 2703 2893 2707
rect 2898 2703 2901 2707
rect 2901 2703 2903 2707
rect 2888 2702 2893 2703
rect 2898 2702 2903 2703
rect 3920 2703 3922 2707
rect 3922 2703 3925 2707
rect 3930 2703 3933 2707
rect 3933 2703 3935 2707
rect 3920 2702 3925 2703
rect 3930 2702 3935 2703
rect 4936 2703 4938 2707
rect 4938 2703 4941 2707
rect 4946 2703 4949 2707
rect 4949 2703 4951 2707
rect 4936 2702 4941 2703
rect 4946 2702 4951 2703
rect 2189 2697 2194 2702
rect 3149 2697 3154 2702
rect 5037 2697 5042 2702
rect 2605 2687 2610 2692
rect 3309 2687 3314 2692
rect 3645 2687 3650 2692
rect 5037 2687 5042 2692
rect 1917 2677 1922 2682
rect 2061 2677 2066 2682
rect 2141 2677 2146 2682
rect 2173 2677 2178 2682
rect 4397 2677 4402 2682
rect 4797 2677 4802 2682
rect 1485 2667 1490 2672
rect 2045 2667 2050 2672
rect 2829 2667 2834 2672
rect 4509 2667 4514 2672
rect 4733 2657 4738 2662
rect 5005 2657 5010 2662
rect 2077 2647 2082 2652
rect 2157 2647 2162 2652
rect 3533 2637 3538 2642
rect 4909 2637 4914 2642
rect 2989 2627 2994 2632
rect 3021 2627 3026 2632
rect 3229 2627 3234 2632
rect 4381 2627 4386 2632
rect 5005 2627 5010 2632
rect 2157 2617 2162 2622
rect 4893 2617 4898 2622
rect 2061 2607 2066 2612
rect 3485 2607 3490 2612
rect 328 2603 330 2607
rect 330 2603 333 2607
rect 338 2603 341 2607
rect 341 2603 343 2607
rect 328 2602 333 2603
rect 338 2602 343 2603
rect 1352 2603 1354 2607
rect 1354 2603 1357 2607
rect 1362 2603 1365 2607
rect 1365 2603 1367 2607
rect 1352 2602 1357 2603
rect 1362 2602 1367 2603
rect 2384 2603 2386 2607
rect 2386 2603 2389 2607
rect 2394 2603 2397 2607
rect 2397 2603 2399 2607
rect 2384 2602 2389 2603
rect 2394 2602 2399 2603
rect 3400 2603 3402 2607
rect 3402 2603 3405 2607
rect 3410 2603 3413 2607
rect 3413 2603 3415 2607
rect 3400 2602 3405 2603
rect 3410 2602 3415 2603
rect 4424 2603 4426 2607
rect 4426 2603 4429 2607
rect 4434 2603 4437 2607
rect 4437 2603 4439 2607
rect 4424 2602 4429 2603
rect 4434 2602 4439 2603
rect 1341 2597 1346 2602
rect 2621 2597 2626 2602
rect 1581 2577 1586 2582
rect 2637 2577 2642 2582
rect 4493 2577 4498 2582
rect 2637 2567 2642 2572
rect 5245 2567 5250 2572
rect 1837 2547 1842 2552
rect 2573 2547 2578 2552
rect 5245 2547 5250 2552
rect 1341 2537 1346 2542
rect 2861 2537 2866 2542
rect 3101 2537 3106 2542
rect 2109 2527 2114 2532
rect 2925 2527 2930 2532
rect 3309 2527 3314 2532
rect 3373 2527 3378 2532
rect 1949 2517 1954 2522
rect 2253 2517 2258 2522
rect 3357 2517 3362 2522
rect 3549 2507 3554 2512
rect 848 2503 850 2507
rect 850 2503 853 2507
rect 858 2503 861 2507
rect 861 2503 863 2507
rect 848 2502 853 2503
rect 858 2502 863 2503
rect 1872 2503 1874 2507
rect 1874 2503 1877 2507
rect 1882 2503 1885 2507
rect 1885 2503 1887 2507
rect 1872 2502 1877 2503
rect 1882 2502 1887 2503
rect 2888 2503 2890 2507
rect 2890 2503 2893 2507
rect 2898 2503 2901 2507
rect 2901 2503 2903 2507
rect 2888 2502 2893 2503
rect 2898 2502 2903 2503
rect 3920 2503 3922 2507
rect 3922 2503 3925 2507
rect 3930 2503 3933 2507
rect 3933 2503 3935 2507
rect 3920 2502 3925 2503
rect 3930 2502 3935 2503
rect 4936 2503 4938 2507
rect 4938 2503 4941 2507
rect 4946 2503 4949 2507
rect 4949 2503 4951 2507
rect 4936 2502 4941 2503
rect 4946 2502 4951 2503
rect 1437 2497 1442 2502
rect 5165 2497 5170 2502
rect 813 2487 818 2492
rect 3037 2487 3042 2492
rect 3213 2487 3218 2492
rect 5165 2487 5170 2492
rect 2045 2477 2050 2482
rect 2861 2477 2866 2482
rect 3005 2477 3010 2482
rect 3197 2477 3202 2482
rect 1565 2457 1570 2462
rect 1629 2457 1634 2462
rect 2013 2457 2018 2462
rect 2109 2457 2114 2462
rect 2477 2457 2482 2462
rect 2525 2457 2530 2462
rect 2141 2447 2146 2452
rect 3037 2457 3042 2462
rect 4261 2447 4266 2452
rect 2093 2437 2098 2442
rect 4845 2437 4850 2442
rect 2205 2427 2210 2432
rect 2621 2427 2626 2432
rect 1629 2417 1634 2422
rect 2509 2417 2514 2422
rect 2557 2417 2562 2422
rect 2205 2407 2210 2412
rect 328 2403 330 2407
rect 330 2403 333 2407
rect 338 2403 341 2407
rect 341 2403 343 2407
rect 328 2402 333 2403
rect 338 2402 343 2403
rect 1352 2403 1354 2407
rect 1354 2403 1357 2407
rect 1362 2403 1365 2407
rect 1365 2403 1367 2407
rect 1352 2402 1357 2403
rect 1362 2402 1367 2403
rect 2384 2403 2386 2407
rect 2386 2403 2389 2407
rect 2394 2403 2397 2407
rect 2397 2403 2399 2407
rect 2384 2402 2389 2403
rect 2394 2402 2399 2403
rect 2701 2407 2706 2412
rect 3037 2407 3042 2412
rect 3400 2403 3402 2407
rect 3402 2403 3405 2407
rect 3410 2403 3413 2407
rect 3413 2403 3415 2407
rect 3400 2402 3405 2403
rect 3410 2402 3415 2403
rect 4424 2403 4426 2407
rect 4426 2403 4429 2407
rect 4434 2403 4437 2407
rect 4437 2403 4439 2407
rect 4424 2402 4429 2403
rect 4434 2402 4439 2403
rect 3197 2397 3202 2402
rect 2829 2387 2834 2392
rect 2669 2377 2674 2382
rect 2797 2377 2802 2382
rect 3197 2377 3202 2382
rect 3325 2377 3330 2382
rect 4925 2377 4930 2382
rect 2125 2357 2130 2362
rect 3037 2367 3042 2372
rect 1421 2337 1426 2342
rect 1453 2337 1458 2342
rect 1853 2337 1858 2342
rect 2797 2337 2802 2342
rect 1757 2317 1762 2322
rect 3037 2327 3042 2332
rect 2045 2307 2050 2312
rect 2173 2307 2178 2312
rect 848 2303 850 2307
rect 850 2303 853 2307
rect 858 2303 861 2307
rect 861 2303 863 2307
rect 848 2302 853 2303
rect 858 2302 863 2303
rect 1872 2303 1874 2307
rect 1874 2303 1877 2307
rect 1882 2303 1885 2307
rect 1885 2303 1887 2307
rect 1872 2302 1877 2303
rect 1882 2302 1887 2303
rect 2888 2303 2890 2307
rect 2890 2303 2893 2307
rect 2898 2303 2901 2307
rect 2901 2303 2903 2307
rect 2888 2302 2893 2303
rect 2898 2302 2903 2303
rect 3920 2303 3922 2307
rect 3922 2303 3925 2307
rect 3930 2303 3933 2307
rect 3933 2303 3935 2307
rect 3920 2302 3925 2303
rect 3930 2302 3935 2303
rect 4936 2303 4938 2307
rect 4938 2303 4941 2307
rect 4946 2303 4949 2307
rect 4949 2303 4951 2307
rect 4936 2302 4941 2303
rect 4946 2302 4951 2303
rect 2765 2297 2770 2302
rect 2445 2277 2450 2282
rect 3277 2277 3282 2282
rect 1965 2267 1970 2272
rect 2477 2267 2482 2272
rect 2669 2267 2674 2272
rect 4717 2257 4722 2262
rect 2669 2247 2674 2252
rect 2685 2247 2690 2252
rect 1645 2237 1650 2242
rect 3853 2237 3858 2242
rect 4045 2237 4050 2242
rect 3261 2227 3266 2232
rect 5277 2227 5282 2232
rect 1789 2217 1794 2222
rect 328 2203 330 2207
rect 330 2203 333 2207
rect 338 2203 341 2207
rect 341 2203 343 2207
rect 328 2202 333 2203
rect 338 2202 343 2203
rect 1352 2203 1354 2207
rect 1354 2203 1357 2207
rect 1362 2203 1365 2207
rect 1365 2203 1367 2207
rect 1352 2202 1357 2203
rect 1362 2202 1367 2203
rect 2269 2207 2274 2212
rect 3325 2207 3330 2212
rect 2384 2203 2386 2207
rect 2386 2203 2389 2207
rect 2394 2203 2397 2207
rect 2397 2203 2399 2207
rect 2384 2202 2389 2203
rect 2394 2202 2399 2203
rect 3400 2203 3402 2207
rect 3402 2203 3405 2207
rect 3410 2203 3413 2207
rect 3413 2203 3415 2207
rect 3400 2202 3405 2203
rect 3410 2202 3415 2203
rect 4424 2203 4426 2207
rect 4426 2203 4429 2207
rect 4434 2203 4437 2207
rect 4437 2203 4439 2207
rect 4424 2202 4429 2203
rect 4434 2202 4439 2203
rect 2333 2197 2338 2202
rect 2301 2187 2306 2192
rect 3277 2187 3282 2192
rect 1597 2177 1602 2182
rect 5197 2167 5202 2172
rect 1997 2157 2002 2162
rect 4157 2157 4162 2162
rect 2317 2147 2322 2152
rect 2781 2137 2786 2142
rect 5213 2137 5218 2142
rect 5181 2127 5186 2132
rect 5213 2127 5218 2132
rect 1709 2117 1714 2122
rect 5229 2107 5234 2112
rect 848 2103 850 2107
rect 850 2103 853 2107
rect 858 2103 861 2107
rect 861 2103 863 2107
rect 848 2102 853 2103
rect 858 2102 863 2103
rect 1872 2103 1874 2107
rect 1874 2103 1877 2107
rect 1882 2103 1885 2107
rect 1885 2103 1887 2107
rect 1872 2102 1877 2103
rect 1882 2102 1887 2103
rect 2888 2103 2890 2107
rect 2890 2103 2893 2107
rect 2898 2103 2901 2107
rect 2901 2103 2903 2107
rect 2888 2102 2893 2103
rect 2898 2102 2903 2103
rect 3920 2103 3922 2107
rect 3922 2103 3925 2107
rect 3930 2103 3933 2107
rect 3933 2103 3935 2107
rect 3920 2102 3925 2103
rect 3930 2102 3935 2103
rect 4936 2103 4938 2107
rect 4938 2103 4941 2107
rect 4946 2103 4949 2107
rect 4949 2103 4951 2107
rect 4936 2102 4941 2103
rect 4946 2102 4951 2103
rect 2189 2097 2194 2102
rect 3885 2097 3890 2102
rect 5245 2097 5250 2102
rect 2589 2087 2594 2092
rect 2141 2067 2146 2072
rect 2973 2067 2978 2072
rect 4157 2067 4162 2072
rect 5229 2067 5234 2072
rect 1341 2057 1346 2062
rect 3597 2057 3602 2062
rect 4701 2057 4706 2062
rect 4357 2027 4362 2032
rect 4605 2027 4610 2032
rect 2157 2007 2162 2012
rect 328 2003 330 2007
rect 330 2003 333 2007
rect 338 2003 341 2007
rect 341 2003 343 2007
rect 328 2002 333 2003
rect 338 2002 343 2003
rect 1352 2003 1354 2007
rect 1354 2003 1357 2007
rect 1362 2003 1365 2007
rect 1365 2003 1367 2007
rect 1352 2002 1357 2003
rect 1362 2002 1367 2003
rect 2384 2003 2386 2007
rect 2386 2003 2389 2007
rect 2394 2003 2397 2007
rect 2397 2003 2399 2007
rect 2384 2002 2389 2003
rect 2394 2002 2399 2003
rect 3400 2003 3402 2007
rect 3402 2003 3405 2007
rect 3410 2003 3413 2007
rect 3413 2003 3415 2007
rect 3400 2002 3405 2003
rect 3410 2002 3415 2003
rect 4424 2003 4426 2007
rect 4426 2003 4429 2007
rect 4434 2003 4437 2007
rect 4437 2003 4439 2007
rect 4424 2002 4429 2003
rect 4434 2002 4439 2003
rect 957 1997 962 2002
rect 1837 1987 1842 1992
rect 2845 1967 2850 1972
rect 3005 1967 3010 1972
rect 1837 1947 1842 1952
rect 1853 1947 1858 1952
rect 2541 1947 2546 1952
rect 4477 1957 4482 1962
rect 5245 1957 5250 1962
rect 3261 1947 3266 1952
rect 2125 1937 2130 1942
rect 3293 1937 3298 1942
rect 4653 1937 4658 1942
rect 2781 1927 2786 1932
rect 4765 1917 4770 1922
rect 5293 1917 5298 1922
rect 3293 1907 3298 1912
rect 848 1903 850 1907
rect 850 1903 853 1907
rect 858 1903 861 1907
rect 861 1903 863 1907
rect 848 1902 853 1903
rect 858 1902 863 1903
rect 1872 1903 1874 1907
rect 1874 1903 1877 1907
rect 1882 1903 1885 1907
rect 1885 1903 1887 1907
rect 1872 1902 1877 1903
rect 1882 1902 1887 1903
rect 2888 1903 2890 1907
rect 2890 1903 2893 1907
rect 2898 1903 2901 1907
rect 2901 1903 2903 1907
rect 2888 1902 2893 1903
rect 2898 1902 2903 1903
rect 3920 1903 3922 1907
rect 3922 1903 3925 1907
rect 3930 1903 3933 1907
rect 3933 1903 3935 1907
rect 3920 1902 3925 1903
rect 3930 1902 3935 1903
rect 2061 1897 2066 1902
rect 4936 1903 4938 1907
rect 4938 1903 4941 1907
rect 4946 1903 4949 1907
rect 4949 1903 4951 1907
rect 4936 1902 4941 1903
rect 4946 1902 4951 1903
rect 5053 1897 5058 1902
rect 1517 1877 1522 1882
rect 2509 1877 2514 1882
rect 2061 1857 2066 1862
rect 5117 1857 5122 1862
rect 5261 1857 5266 1862
rect 1469 1847 1474 1852
rect 4557 1817 4562 1822
rect 3853 1807 3858 1812
rect 4589 1807 4594 1812
rect 328 1803 330 1807
rect 330 1803 333 1807
rect 338 1803 341 1807
rect 341 1803 343 1807
rect 328 1802 333 1803
rect 338 1802 343 1803
rect 1352 1803 1354 1807
rect 1354 1803 1357 1807
rect 1362 1803 1365 1807
rect 1365 1803 1367 1807
rect 1352 1802 1357 1803
rect 1362 1802 1367 1803
rect 2384 1803 2386 1807
rect 2386 1803 2389 1807
rect 2394 1803 2397 1807
rect 2397 1803 2399 1807
rect 2384 1802 2389 1803
rect 2394 1802 2399 1803
rect 3400 1803 3402 1807
rect 3402 1803 3405 1807
rect 3410 1803 3413 1807
rect 3413 1803 3415 1807
rect 3400 1802 3405 1803
rect 3410 1802 3415 1803
rect 4424 1803 4426 1807
rect 4426 1803 4429 1807
rect 4434 1803 4437 1807
rect 4437 1803 4439 1807
rect 4424 1802 4429 1803
rect 4434 1802 4439 1803
rect 1917 1797 1922 1802
rect 1965 1797 1970 1802
rect 2029 1777 2034 1782
rect 4493 1777 4498 1782
rect 2813 1757 2818 1762
rect 4061 1757 4066 1762
rect 1485 1747 1490 1752
rect 3629 1747 3634 1752
rect 2141 1727 2146 1732
rect 5181 1727 5186 1732
rect 2285 1707 2290 1712
rect 848 1703 850 1707
rect 850 1703 853 1707
rect 858 1703 861 1707
rect 861 1703 863 1707
rect 848 1702 853 1703
rect 858 1702 863 1703
rect 1872 1703 1874 1707
rect 1874 1703 1877 1707
rect 1882 1703 1885 1707
rect 1885 1703 1887 1707
rect 1872 1702 1877 1703
rect 1882 1702 1887 1703
rect 2888 1703 2890 1707
rect 2890 1703 2893 1707
rect 2898 1703 2901 1707
rect 2901 1703 2903 1707
rect 2888 1702 2893 1703
rect 2898 1702 2903 1703
rect 3920 1703 3922 1707
rect 3922 1703 3925 1707
rect 3930 1703 3933 1707
rect 3933 1703 3935 1707
rect 3920 1702 3925 1703
rect 3930 1702 3935 1703
rect 4936 1703 4938 1707
rect 4938 1703 4941 1707
rect 4946 1703 4949 1707
rect 4949 1703 4951 1707
rect 4936 1702 4941 1703
rect 4946 1702 4951 1703
rect 2605 1697 2610 1702
rect 3229 1697 3234 1702
rect 1677 1687 1682 1692
rect 5085 1687 5090 1692
rect 1645 1667 1650 1672
rect 1229 1637 1234 1642
rect 5133 1637 5138 1642
rect 5261 1637 5266 1642
rect 1565 1627 1570 1632
rect 2077 1617 2082 1622
rect 328 1603 330 1607
rect 330 1603 333 1607
rect 338 1603 341 1607
rect 341 1603 343 1607
rect 328 1602 333 1603
rect 338 1602 343 1603
rect 1352 1603 1354 1607
rect 1354 1603 1357 1607
rect 1362 1603 1365 1607
rect 1365 1603 1367 1607
rect 1352 1602 1357 1603
rect 1362 1602 1367 1603
rect 2384 1603 2386 1607
rect 2386 1603 2389 1607
rect 2394 1603 2397 1607
rect 2397 1603 2399 1607
rect 2384 1602 2389 1603
rect 2394 1602 2399 1603
rect 3400 1603 3402 1607
rect 3402 1603 3405 1607
rect 3410 1603 3413 1607
rect 3413 1603 3415 1607
rect 3400 1602 3405 1603
rect 3410 1602 3415 1603
rect 4424 1603 4426 1607
rect 4426 1603 4429 1607
rect 4434 1603 4437 1607
rect 4437 1603 4439 1607
rect 4424 1602 4429 1603
rect 4434 1602 4439 1603
rect 3021 1597 3026 1602
rect 2157 1577 2162 1582
rect 3533 1577 3538 1582
rect 2477 1567 2482 1572
rect 3357 1567 3362 1572
rect 4381 1567 4386 1572
rect 4573 1567 4578 1572
rect 2173 1557 2178 1562
rect 1725 1547 1730 1552
rect 2461 1547 2466 1552
rect 2253 1537 2258 1542
rect 3805 1537 3810 1542
rect 4253 1537 4258 1542
rect 717 1527 722 1532
rect 2989 1527 2994 1532
rect 4365 1517 4370 1522
rect 4733 1517 4738 1522
rect 4397 1507 4402 1512
rect 848 1503 850 1507
rect 850 1503 853 1507
rect 858 1503 861 1507
rect 861 1503 863 1507
rect 848 1502 853 1503
rect 858 1502 863 1503
rect 1872 1503 1874 1507
rect 1874 1503 1877 1507
rect 1882 1503 1885 1507
rect 1885 1503 1887 1507
rect 1872 1502 1877 1503
rect 1882 1502 1887 1503
rect 2888 1503 2890 1507
rect 2890 1503 2893 1507
rect 2898 1503 2901 1507
rect 2901 1503 2903 1507
rect 2888 1502 2893 1503
rect 2898 1502 2903 1503
rect 3920 1503 3922 1507
rect 3922 1503 3925 1507
rect 3930 1503 3933 1507
rect 3933 1503 3935 1507
rect 3920 1502 3925 1503
rect 3930 1502 3935 1503
rect 4936 1503 4938 1507
rect 4938 1503 4941 1507
rect 4946 1503 4949 1507
rect 4949 1503 4951 1507
rect 4936 1502 4941 1503
rect 4946 1502 4951 1503
rect 1837 1497 1842 1502
rect 1373 1487 1378 1492
rect 2013 1477 2018 1482
rect 4413 1477 4418 1482
rect 1581 1467 1586 1472
rect 1517 1457 1522 1462
rect 3645 1467 3650 1472
rect 4861 1467 4866 1472
rect 1901 1457 1906 1462
rect 3293 1457 3298 1462
rect 2317 1447 2322 1452
rect 3053 1437 3058 1442
rect 4989 1427 4994 1432
rect 5037 1427 5042 1432
rect 5133 1427 5138 1432
rect 2269 1417 2274 1422
rect 4525 1417 4530 1422
rect 328 1403 330 1407
rect 330 1403 333 1407
rect 338 1403 341 1407
rect 341 1403 343 1407
rect 328 1402 333 1403
rect 338 1402 343 1403
rect 1352 1403 1354 1407
rect 1354 1403 1357 1407
rect 1362 1403 1365 1407
rect 1365 1403 1367 1407
rect 1352 1402 1357 1403
rect 1362 1402 1367 1403
rect 2384 1403 2386 1407
rect 2386 1403 2389 1407
rect 2394 1403 2397 1407
rect 2397 1403 2399 1407
rect 2384 1402 2389 1403
rect 2394 1402 2399 1403
rect 3400 1403 3402 1407
rect 3402 1403 3405 1407
rect 3410 1403 3413 1407
rect 3413 1403 3415 1407
rect 3400 1402 3405 1403
rect 3410 1402 3415 1403
rect 4424 1403 4426 1407
rect 4426 1403 4429 1407
rect 4434 1403 4437 1407
rect 4437 1403 4439 1407
rect 4424 1402 4429 1403
rect 4434 1402 4439 1403
rect 2093 1377 2098 1382
rect 3981 1377 3986 1382
rect 2509 1367 2514 1372
rect 3357 1367 3362 1372
rect 3597 1367 3602 1372
rect 4717 1367 4722 1372
rect 2525 1357 2530 1362
rect 3341 1357 3346 1362
rect 1757 1347 1762 1352
rect 2509 1347 2514 1352
rect 4205 1347 4210 1352
rect 2541 1337 2546 1342
rect 4045 1327 4050 1332
rect 2909 1307 2914 1312
rect 848 1303 850 1307
rect 850 1303 853 1307
rect 858 1303 861 1307
rect 861 1303 863 1307
rect 848 1302 853 1303
rect 858 1302 863 1303
rect 1872 1303 1874 1307
rect 1874 1303 1877 1307
rect 1882 1303 1885 1307
rect 1885 1303 1887 1307
rect 1872 1302 1877 1303
rect 1882 1302 1887 1303
rect 2888 1303 2890 1307
rect 2890 1303 2893 1307
rect 2898 1303 2901 1307
rect 2901 1303 2903 1307
rect 2888 1302 2893 1303
rect 2898 1302 2903 1303
rect 3920 1303 3922 1307
rect 3922 1303 3925 1307
rect 3930 1303 3933 1307
rect 3933 1303 3935 1307
rect 3920 1302 3925 1303
rect 3930 1302 3935 1303
rect 4936 1303 4938 1307
rect 4938 1303 4941 1307
rect 4946 1303 4949 1307
rect 4949 1303 4951 1307
rect 4936 1302 4941 1303
rect 4946 1302 4951 1303
rect 3805 1297 3810 1302
rect 1437 1277 1442 1282
rect 2909 1277 2914 1282
rect 1069 1267 1074 1272
rect 1325 1267 1330 1272
rect 2061 1267 2066 1272
rect 2445 1247 2450 1252
rect 3805 1257 3810 1262
rect 4349 1247 4354 1252
rect 3309 1227 3314 1232
rect 5037 1227 5042 1232
rect 328 1203 330 1207
rect 330 1203 333 1207
rect 338 1203 341 1207
rect 341 1203 343 1207
rect 328 1202 333 1203
rect 338 1202 343 1203
rect 1352 1203 1354 1207
rect 1354 1203 1357 1207
rect 1362 1203 1365 1207
rect 1365 1203 1367 1207
rect 1352 1202 1357 1203
rect 1362 1202 1367 1203
rect 2384 1203 2386 1207
rect 2386 1203 2389 1207
rect 2394 1203 2397 1207
rect 2397 1203 2399 1207
rect 2384 1202 2389 1203
rect 2394 1202 2399 1203
rect 3400 1203 3402 1207
rect 3402 1203 3405 1207
rect 3410 1203 3413 1207
rect 3413 1203 3415 1207
rect 3400 1202 3405 1203
rect 3410 1202 3415 1203
rect 4424 1203 4426 1207
rect 4426 1203 4429 1207
rect 4434 1203 4437 1207
rect 4437 1203 4439 1207
rect 4424 1202 4429 1203
rect 4434 1202 4439 1203
rect 1309 1197 1314 1202
rect 2637 1197 2642 1202
rect 1341 1187 1346 1192
rect 2253 1187 2258 1192
rect 3373 1187 3378 1192
rect 4173 1177 4178 1182
rect 5213 1177 5218 1182
rect 3261 1147 3266 1152
rect 3309 1147 3314 1152
rect 5277 1157 5282 1162
rect 2781 1137 2786 1142
rect 5165 1137 5170 1142
rect 4829 1127 4834 1132
rect 1709 1117 1714 1122
rect 5085 1117 5090 1122
rect 2125 1107 2130 1112
rect 848 1103 850 1107
rect 850 1103 853 1107
rect 858 1103 861 1107
rect 861 1103 863 1107
rect 848 1102 853 1103
rect 858 1102 863 1103
rect 1872 1103 1874 1107
rect 1874 1103 1877 1107
rect 1882 1103 1885 1107
rect 1885 1103 1887 1107
rect 1872 1102 1877 1103
rect 1882 1102 1887 1103
rect 2888 1103 2890 1107
rect 2890 1103 2893 1107
rect 2898 1103 2901 1107
rect 2901 1103 2903 1107
rect 2888 1102 2893 1103
rect 2898 1102 2903 1103
rect 3920 1103 3922 1107
rect 3922 1103 3925 1107
rect 3930 1103 3933 1107
rect 3933 1103 3935 1107
rect 3920 1102 3925 1103
rect 3930 1102 3935 1103
rect 4936 1103 4938 1107
rect 4938 1103 4941 1107
rect 4946 1103 4949 1107
rect 4949 1103 4951 1107
rect 4936 1102 4941 1103
rect 4946 1102 4951 1103
rect 4925 1067 4930 1072
rect 4189 1047 4194 1052
rect 4365 1037 4370 1042
rect 2413 1007 2418 1012
rect 328 1003 330 1007
rect 330 1003 333 1007
rect 338 1003 341 1007
rect 341 1003 343 1007
rect 328 1002 333 1003
rect 338 1002 343 1003
rect 1352 1003 1354 1007
rect 1354 1003 1357 1007
rect 1362 1003 1365 1007
rect 1365 1003 1367 1007
rect 1352 1002 1357 1003
rect 1362 1002 1367 1003
rect 2384 1003 2386 1007
rect 2386 1003 2389 1007
rect 2394 1003 2397 1007
rect 2397 1003 2399 1007
rect 2384 1002 2389 1003
rect 2394 1002 2399 1003
rect 3400 1003 3402 1007
rect 3402 1003 3405 1007
rect 3410 1003 3413 1007
rect 3413 1003 3415 1007
rect 3400 1002 3405 1003
rect 3410 1002 3415 1003
rect 4424 1003 4426 1007
rect 4426 1003 4429 1007
rect 4434 1003 4437 1007
rect 4437 1003 4439 1007
rect 4424 1002 4429 1003
rect 4434 1002 4439 1003
rect 5277 987 5282 992
rect 5293 977 5298 982
rect 813 967 818 972
rect 5069 967 5074 972
rect 1117 947 1122 952
rect 1821 957 1826 962
rect 2317 957 2322 962
rect 1437 947 1442 952
rect 2781 927 2786 932
rect 1965 917 1970 922
rect 2973 907 2978 912
rect 848 903 850 907
rect 850 903 853 907
rect 858 903 861 907
rect 861 903 863 907
rect 848 902 853 903
rect 858 902 863 903
rect 1872 903 1874 907
rect 1874 903 1877 907
rect 1882 903 1885 907
rect 1885 903 1887 907
rect 1872 902 1877 903
rect 1882 902 1887 903
rect 2888 903 2890 907
rect 2890 903 2893 907
rect 2898 903 2901 907
rect 2901 903 2903 907
rect 2888 902 2893 903
rect 2898 902 2903 903
rect 3920 903 3922 907
rect 3922 903 3925 907
rect 3930 903 3933 907
rect 3933 903 3935 907
rect 3920 902 3925 903
rect 3930 902 3935 903
rect 4936 903 4938 907
rect 4938 903 4941 907
rect 4946 903 4949 907
rect 4949 903 4951 907
rect 4936 902 4941 903
rect 4946 902 4951 903
rect 2925 887 2930 892
rect 4621 887 4626 892
rect 5181 867 5186 872
rect 1613 857 1618 862
rect 2989 857 2994 862
rect 328 803 330 807
rect 330 803 333 807
rect 338 803 341 807
rect 341 803 343 807
rect 328 802 333 803
rect 338 802 343 803
rect 1352 803 1354 807
rect 1354 803 1357 807
rect 1362 803 1365 807
rect 1365 803 1367 807
rect 1352 802 1357 803
rect 1362 802 1367 803
rect 2384 803 2386 807
rect 2386 803 2389 807
rect 2394 803 2397 807
rect 2397 803 2399 807
rect 2384 802 2389 803
rect 2394 802 2399 803
rect 3400 803 3402 807
rect 3402 803 3405 807
rect 3410 803 3413 807
rect 3413 803 3415 807
rect 3400 802 3405 803
rect 3410 802 3415 803
rect 4424 803 4426 807
rect 4426 803 4429 807
rect 4434 803 4437 807
rect 4437 803 4439 807
rect 4424 802 4429 803
rect 4434 802 4439 803
rect 1821 777 1826 782
rect 4957 767 4962 772
rect 1229 757 1234 762
rect 3149 757 3154 762
rect 4685 757 4690 762
rect 5101 737 5106 742
rect 848 703 850 707
rect 850 703 853 707
rect 858 703 861 707
rect 861 703 863 707
rect 848 702 853 703
rect 858 702 863 703
rect 1872 703 1874 707
rect 1874 703 1877 707
rect 1882 703 1885 707
rect 1885 703 1887 707
rect 1872 702 1877 703
rect 1882 702 1887 703
rect 2888 703 2890 707
rect 2890 703 2893 707
rect 2898 703 2901 707
rect 2901 703 2903 707
rect 2888 702 2893 703
rect 2898 702 2903 703
rect 3920 703 3922 707
rect 3922 703 3925 707
rect 3930 703 3933 707
rect 3933 703 3935 707
rect 3920 702 3925 703
rect 3930 702 3935 703
rect 4936 703 4938 707
rect 4938 703 4941 707
rect 4946 703 4949 707
rect 4949 703 4951 707
rect 4936 702 4941 703
rect 4946 702 4951 703
rect 1373 677 1378 682
rect 3453 677 3458 682
rect 5005 677 5010 682
rect 4093 647 4098 652
rect 4813 647 4818 652
rect 328 603 330 607
rect 330 603 333 607
rect 338 603 341 607
rect 341 603 343 607
rect 328 602 333 603
rect 338 602 343 603
rect 1352 603 1354 607
rect 1354 603 1357 607
rect 1362 603 1365 607
rect 1365 603 1367 607
rect 1352 602 1357 603
rect 1362 602 1367 603
rect 2384 603 2386 607
rect 2386 603 2389 607
rect 2394 603 2397 607
rect 2397 603 2399 607
rect 2384 602 2389 603
rect 2394 602 2399 603
rect 3400 603 3402 607
rect 3402 603 3405 607
rect 3410 603 3413 607
rect 3413 603 3415 607
rect 3400 602 3405 603
rect 3410 602 3415 603
rect 4424 603 4426 607
rect 4426 603 4429 607
rect 4434 603 4437 607
rect 4437 603 4439 607
rect 4424 602 4429 603
rect 4434 602 4439 603
rect 957 567 962 572
rect 4205 567 4210 572
rect 5021 567 5026 572
rect 2029 557 2034 562
rect 2093 547 2098 552
rect 4557 547 4562 552
rect 848 503 850 507
rect 850 503 853 507
rect 858 503 861 507
rect 861 503 863 507
rect 848 502 853 503
rect 858 502 863 503
rect 1872 503 1874 507
rect 1874 503 1877 507
rect 1882 503 1885 507
rect 1885 503 1887 507
rect 1872 502 1877 503
rect 1882 502 1887 503
rect 2888 503 2890 507
rect 2890 503 2893 507
rect 2898 503 2901 507
rect 2901 503 2903 507
rect 2888 502 2893 503
rect 2898 502 2903 503
rect 3920 503 3922 507
rect 3922 503 3925 507
rect 3930 503 3933 507
rect 3933 503 3935 507
rect 3920 502 3925 503
rect 3930 502 3935 503
rect 4936 503 4938 507
rect 4938 503 4941 507
rect 4946 503 4949 507
rect 4949 503 4951 507
rect 4936 502 4941 503
rect 4946 502 4951 503
rect 5197 467 5202 472
rect 5229 447 5234 452
rect 1965 437 1970 442
rect 328 403 330 407
rect 330 403 333 407
rect 338 403 341 407
rect 341 403 343 407
rect 328 402 333 403
rect 338 402 343 403
rect 1352 403 1354 407
rect 1354 403 1357 407
rect 1362 403 1365 407
rect 1365 403 1367 407
rect 1352 402 1357 403
rect 1362 402 1367 403
rect 2384 403 2386 407
rect 2386 403 2389 407
rect 2394 403 2397 407
rect 2397 403 2399 407
rect 2384 402 2389 403
rect 2394 402 2399 403
rect 3400 403 3402 407
rect 3402 403 3405 407
rect 3410 403 3413 407
rect 3413 403 3415 407
rect 3400 402 3405 403
rect 3410 402 3415 403
rect 4424 403 4426 407
rect 4426 403 4429 407
rect 4434 403 4437 407
rect 4437 403 4439 407
rect 4424 402 4429 403
rect 4434 402 4439 403
rect 2637 377 2642 382
rect 3981 357 3986 362
rect 848 303 850 307
rect 850 303 853 307
rect 858 303 861 307
rect 861 303 863 307
rect 848 302 853 303
rect 858 302 863 303
rect 1872 303 1874 307
rect 1874 303 1877 307
rect 1882 303 1885 307
rect 1885 303 1887 307
rect 1872 302 1877 303
rect 1882 302 1887 303
rect 2888 303 2890 307
rect 2890 303 2893 307
rect 2898 303 2901 307
rect 2901 303 2903 307
rect 2888 302 2893 303
rect 2898 302 2903 303
rect 3920 303 3922 307
rect 3922 303 3925 307
rect 3930 303 3933 307
rect 3933 303 3935 307
rect 3920 302 3925 303
rect 3930 302 3935 303
rect 4936 303 4938 307
rect 4938 303 4941 307
rect 4946 303 4949 307
rect 4949 303 4951 307
rect 4936 302 4941 303
rect 4946 302 4951 303
rect 4797 287 4802 292
rect 3997 277 4002 282
rect 1973 267 1978 272
rect 5037 267 5042 272
rect 4877 257 4882 262
rect 328 203 330 207
rect 330 203 333 207
rect 338 203 341 207
rect 341 203 343 207
rect 328 202 333 203
rect 338 202 343 203
rect 1352 203 1354 207
rect 1354 203 1357 207
rect 1362 203 1365 207
rect 1365 203 1367 207
rect 1352 202 1357 203
rect 1362 202 1367 203
rect 2384 203 2386 207
rect 2386 203 2389 207
rect 2394 203 2397 207
rect 2397 203 2399 207
rect 2384 202 2389 203
rect 2394 202 2399 203
rect 3400 203 3402 207
rect 3402 203 3405 207
rect 3410 203 3413 207
rect 3413 203 3415 207
rect 3400 202 3405 203
rect 3410 202 3415 203
rect 4424 203 4426 207
rect 4426 203 4429 207
rect 4434 203 4437 207
rect 4437 203 4439 207
rect 4424 202 4429 203
rect 4434 202 4439 203
rect 5085 197 5090 202
rect 5245 147 5250 152
rect 5293 147 5298 152
rect 5261 127 5266 132
rect 4973 117 4978 122
rect 848 103 850 107
rect 850 103 853 107
rect 858 103 861 107
rect 861 103 863 107
rect 848 102 853 103
rect 858 102 863 103
rect 1872 103 1874 107
rect 1874 103 1877 107
rect 1882 103 1885 107
rect 1885 103 1887 107
rect 1872 102 1877 103
rect 1882 102 1887 103
rect 2888 103 2890 107
rect 2890 103 2893 107
rect 2898 103 2901 107
rect 2901 103 2903 107
rect 2888 102 2893 103
rect 2898 102 2903 103
rect 3920 103 3922 107
rect 3922 103 3925 107
rect 3930 103 3933 107
rect 3933 103 3935 107
rect 3920 102 3925 103
rect 3930 102 3935 103
rect 4936 103 4938 107
rect 4938 103 4941 107
rect 4946 103 4949 107
rect 4949 103 4951 107
rect 4936 102 4941 103
rect 4946 102 4951 103
rect 5149 87 5154 92
rect 4669 77 4674 82
rect 5133 57 5138 62
rect 328 3 330 7
rect 330 3 333 7
rect 338 3 341 7
rect 341 3 343 7
rect 328 2 333 3
rect 338 2 343 3
rect 1352 3 1354 7
rect 1354 3 1357 7
rect 1362 3 1365 7
rect 1365 3 1367 7
rect 1352 2 1357 3
rect 1362 2 1367 3
rect 2384 3 2386 7
rect 2386 3 2389 7
rect 2394 3 2397 7
rect 2397 3 2399 7
rect 2384 2 2389 3
rect 2394 2 2399 3
rect 3400 3 3402 7
rect 3402 3 3405 7
rect 3410 3 3413 7
rect 3413 3 3415 7
rect 3400 2 3405 3
rect 3410 2 3415 3
rect 4424 3 4426 7
rect 4426 3 4429 7
rect 4434 3 4437 7
rect 4437 3 4439 7
rect 4424 2 4429 3
rect 4434 2 4439 3
<< metal6 >>
rect 328 5007 344 5130
rect 333 5002 338 5007
rect 343 5002 344 5007
rect 328 4807 344 5002
rect 333 4802 338 4807
rect 343 4802 344 4807
rect 328 4607 344 4802
rect 333 4602 338 4607
rect 343 4602 344 4607
rect 328 4407 344 4602
rect 333 4402 338 4407
rect 343 4402 344 4407
rect 328 4207 344 4402
rect 333 4202 338 4207
rect 343 4202 344 4207
rect 328 4007 344 4202
rect 333 4002 338 4007
rect 343 4002 344 4007
rect 328 3807 344 4002
rect 333 3802 338 3807
rect 343 3802 344 3807
rect 328 3607 344 3802
rect 333 3602 338 3607
rect 343 3602 344 3607
rect 328 3407 344 3602
rect 333 3402 338 3407
rect 343 3402 344 3407
rect 328 3207 344 3402
rect 333 3202 338 3207
rect 343 3202 344 3207
rect 328 3007 344 3202
rect 333 3002 338 3007
rect 343 3002 344 3007
rect 328 2807 344 3002
rect 848 5107 864 5130
rect 853 5102 858 5107
rect 863 5102 864 5107
rect 848 4907 864 5102
rect 853 4902 858 4907
rect 863 4902 864 4907
rect 848 4707 864 4902
rect 853 4702 858 4707
rect 863 4702 864 4707
rect 848 4507 864 4702
rect 853 4502 858 4507
rect 863 4502 864 4507
rect 848 4307 864 4502
rect 853 4302 858 4307
rect 863 4302 864 4307
rect 848 4107 864 4302
rect 853 4102 858 4107
rect 863 4102 864 4107
rect 848 3907 864 4102
rect 853 3902 858 3907
rect 863 3902 864 3907
rect 848 3707 864 3902
rect 1352 5007 1368 5130
rect 1357 5002 1362 5007
rect 1367 5002 1368 5007
rect 1352 4807 1368 5002
rect 1357 4802 1362 4807
rect 1367 4802 1368 4807
rect 1352 4607 1368 4802
rect 1357 4602 1362 4607
rect 1367 4602 1368 4607
rect 1352 4407 1368 4602
rect 1357 4402 1362 4407
rect 1367 4402 1368 4407
rect 1352 4207 1368 4402
rect 1872 5107 1888 5130
rect 1877 5102 1882 5107
rect 1887 5102 1888 5107
rect 1872 4907 1888 5102
rect 1877 4902 1882 4907
rect 1887 4902 1888 4907
rect 1872 4707 1888 4902
rect 1877 4702 1882 4707
rect 1887 4702 1888 4707
rect 1872 4507 1888 4702
rect 1877 4502 1882 4507
rect 1887 4502 1888 4507
rect 1357 4202 1362 4207
rect 1367 4202 1368 4207
rect 1352 4007 1368 4202
rect 1357 4002 1362 4007
rect 1367 4002 1368 4007
rect 1352 3807 1368 4002
rect 1357 3802 1362 3807
rect 1367 3802 1368 3807
rect 853 3702 858 3707
rect 863 3702 864 3707
rect 848 3507 864 3702
rect 853 3502 858 3507
rect 863 3502 864 3507
rect 848 3307 864 3502
rect 853 3302 858 3307
rect 863 3302 864 3307
rect 848 3107 864 3302
rect 853 3102 858 3107
rect 863 3102 864 3107
rect 848 2907 864 3102
rect 853 2902 858 2907
rect 863 2902 864 2907
rect 714 2867 722 2872
rect 333 2802 338 2807
rect 343 2802 344 2807
rect 328 2607 344 2802
rect 333 2602 338 2607
rect 343 2602 344 2607
rect 328 2407 344 2602
rect 333 2402 338 2407
rect 343 2402 344 2407
rect 328 2207 344 2402
rect 333 2202 338 2207
rect 343 2202 344 2207
rect 328 2007 344 2202
rect 333 2002 338 2007
rect 343 2002 344 2007
rect 328 1807 344 2002
rect 333 1802 338 1807
rect 343 1802 344 1807
rect 328 1607 344 1802
rect 333 1602 338 1607
rect 343 1602 344 1607
rect 328 1407 344 1602
rect 717 1532 722 2867
rect 848 2707 864 2902
rect 853 2702 858 2707
rect 863 2702 864 2707
rect 848 2507 864 2702
rect 853 2502 858 2507
rect 863 2502 864 2507
rect 333 1402 338 1407
rect 343 1402 344 1407
rect 328 1207 344 1402
rect 333 1202 338 1207
rect 343 1202 344 1207
rect 328 1007 344 1202
rect 333 1002 338 1007
rect 343 1002 344 1007
rect 328 807 344 1002
rect 813 972 818 2487
rect 848 2307 864 2502
rect 853 2302 858 2307
rect 863 2302 864 2307
rect 848 2107 864 2302
rect 853 2102 858 2107
rect 863 2102 864 2107
rect 848 1907 864 2102
rect 853 1902 858 1907
rect 863 1902 864 1907
rect 848 1707 864 1902
rect 853 1702 858 1707
rect 863 1702 864 1707
rect 848 1507 864 1702
rect 853 1502 858 1507
rect 863 1502 864 1507
rect 848 1307 864 1502
rect 853 1302 858 1307
rect 863 1302 864 1307
rect 848 1107 864 1302
rect 853 1102 858 1107
rect 863 1102 864 1107
rect 333 802 338 807
rect 343 802 344 807
rect 328 607 344 802
rect 333 602 338 607
rect 343 602 344 607
rect 328 407 344 602
rect 333 402 338 407
rect 343 402 344 407
rect 328 207 344 402
rect 333 202 338 207
rect 343 202 344 207
rect 328 7 344 202
rect 333 2 338 7
rect 343 2 344 7
rect 328 -30 344 2
rect 848 907 864 1102
rect 853 902 858 907
rect 863 902 864 907
rect 848 707 864 902
rect 853 702 858 707
rect 863 702 864 707
rect 848 507 864 702
rect 957 572 962 1997
rect 1069 1272 1074 3707
rect 1117 952 1122 3637
rect 1352 3607 1368 3802
rect 1357 3602 1362 3607
rect 1367 3602 1368 3607
rect 1325 2852 1330 3447
rect 1229 762 1234 1637
rect 1309 1202 1314 2837
rect 1325 1272 1330 2847
rect 1352 3407 1368 3602
rect 1357 3402 1362 3407
rect 1367 3402 1368 3407
rect 1352 3207 1368 3402
rect 1357 3202 1362 3207
rect 1367 3202 1368 3207
rect 1352 3007 1368 3202
rect 1357 3002 1362 3007
rect 1367 3002 1368 3007
rect 1352 2807 1368 3002
rect 1453 2952 1458 4357
rect 1872 4307 1888 4502
rect 2384 5007 2400 5130
rect 2389 5002 2394 5007
rect 2399 5002 2400 5007
rect 2384 4807 2400 5002
rect 2389 4802 2394 4807
rect 2399 4802 2400 4807
rect 2384 4607 2400 4802
rect 2389 4602 2394 4607
rect 2399 4602 2400 4607
rect 1877 4302 1882 4307
rect 1887 4302 1888 4307
rect 1677 4267 1685 4272
rect 1357 2802 1362 2807
rect 1367 2802 1368 2807
rect 1352 2607 1368 2802
rect 1373 2802 1378 2867
rect 1357 2602 1362 2607
rect 1367 2602 1368 2607
rect 1341 2542 1346 2597
rect 1352 2407 1368 2602
rect 1357 2402 1362 2407
rect 1367 2402 1368 2407
rect 1352 2207 1368 2402
rect 1421 2342 1426 2707
rect 1357 2202 1362 2207
rect 1367 2202 1368 2207
rect 1341 1192 1346 2057
rect 1352 2007 1368 2202
rect 1357 2002 1362 2007
rect 1367 2002 1368 2007
rect 1352 1807 1368 2002
rect 1357 1802 1362 1807
rect 1367 1802 1368 1807
rect 1352 1607 1368 1802
rect 1357 1602 1362 1607
rect 1367 1602 1368 1607
rect 1352 1407 1368 1602
rect 1357 1402 1362 1407
rect 1367 1402 1368 1407
rect 1352 1207 1368 1402
rect 1357 1202 1362 1207
rect 1367 1202 1368 1207
rect 1352 1007 1368 1202
rect 1357 1002 1362 1007
rect 1367 1002 1368 1007
rect 1352 807 1368 1002
rect 1357 802 1362 807
rect 1367 802 1368 807
rect 1352 607 1368 802
rect 1373 682 1378 1487
rect 1437 1282 1442 2497
rect 1453 2342 1458 2897
rect 1469 1852 1474 3997
rect 1485 2672 1490 3597
rect 1485 1752 1490 2667
rect 1517 1882 1522 3007
rect 1597 2972 1602 4057
rect 1517 1462 1522 1877
rect 1565 1632 1570 2457
rect 1581 1472 1586 2577
rect 1597 2182 1602 2967
rect 1437 952 1442 1277
rect 1613 862 1618 3737
rect 1645 3332 1650 3567
rect 1629 2422 1634 2457
rect 1645 1672 1650 2237
rect 1677 1692 1682 4267
rect 1872 4107 1888 4302
rect 1877 4102 1882 4107
rect 1887 4102 1888 4107
rect 1872 3907 1888 4102
rect 1877 3902 1882 3907
rect 1887 3902 1888 3907
rect 1872 3707 1888 3902
rect 1877 3702 1882 3707
rect 1887 3702 1888 3707
rect 1741 3562 1746 3647
rect 1741 2862 1746 3557
rect 1789 3647 1797 3652
rect 1773 2862 1778 2907
rect 1709 1122 1714 2117
rect 1725 1552 1730 2747
rect 1757 1352 1762 2317
rect 1789 2222 1794 3647
rect 1872 3507 1888 3702
rect 1877 3502 1882 3507
rect 1887 3502 1888 3507
rect 1872 3307 1888 3502
rect 1877 3302 1882 3307
rect 1887 3302 1888 3307
rect 1872 3107 1888 3302
rect 1877 3102 1882 3107
rect 1887 3102 1888 3107
rect 1872 2907 1888 3102
rect 1877 2902 1882 2907
rect 1887 2902 1888 2907
rect 1821 962 1826 2777
rect 1872 2707 1888 2902
rect 1877 2702 1882 2707
rect 1887 2702 1888 2707
rect 1837 1992 1842 2547
rect 1872 2507 1888 2702
rect 1877 2502 1882 2507
rect 1887 2502 1888 2507
rect 1853 1952 1858 2337
rect 1872 2307 1888 2502
rect 1877 2302 1882 2307
rect 1887 2302 1888 2307
rect 1872 2107 1888 2302
rect 1877 2102 1882 2107
rect 1887 2102 1888 2107
rect 1837 1502 1842 1947
rect 1872 1907 1888 2102
rect 1877 1902 1882 1907
rect 1887 1902 1888 1907
rect 1872 1707 1888 1902
rect 1877 1702 1882 1707
rect 1887 1702 1888 1707
rect 1872 1507 1888 1702
rect 1877 1502 1882 1507
rect 1887 1502 1888 1507
rect 1821 782 1826 957
rect 1872 1307 1888 1502
rect 1901 1462 1906 3497
rect 1917 2682 1922 3047
rect 1917 1802 1922 2677
rect 1949 2522 1954 3057
rect 1965 2852 1970 3857
rect 1965 2272 1970 2847
rect 1997 2162 2002 3867
rect 2061 2682 2066 4457
rect 2384 4407 2400 4602
rect 2888 5107 2904 5130
rect 2893 5102 2898 5107
rect 2903 5102 2904 5107
rect 2888 4907 2904 5102
rect 2893 4902 2898 4907
rect 2903 4902 2904 4907
rect 2888 4707 2904 4902
rect 2893 4702 2898 4707
rect 2903 4702 2904 4707
rect 2888 4507 2904 4702
rect 2893 4502 2898 4507
rect 2903 4502 2904 4507
rect 2389 4402 2394 4407
rect 2399 4402 2400 4407
rect 2045 2482 2050 2667
rect 2077 2652 2082 4287
rect 2384 4207 2400 4402
rect 2389 4202 2394 4207
rect 2399 4202 2400 4207
rect 2384 4007 2400 4202
rect 2389 4002 2394 4007
rect 2399 4002 2400 4007
rect 2384 3807 2400 4002
rect 2389 3802 2394 3807
rect 2399 3802 2400 3807
rect 2109 3152 2114 3627
rect 1877 1302 1882 1307
rect 1887 1302 1888 1307
rect 1872 1107 1888 1302
rect 1877 1102 1882 1107
rect 1887 1102 1888 1107
rect 1872 907 1888 1102
rect 1877 902 1882 907
rect 1887 902 1888 907
rect 1872 707 1888 902
rect 1877 702 1882 707
rect 1887 702 1888 707
rect 1357 602 1362 607
rect 1367 602 1368 607
rect 853 502 858 507
rect 863 502 864 507
rect 848 307 864 502
rect 853 302 858 307
rect 863 302 864 307
rect 848 107 864 302
rect 853 102 858 107
rect 863 102 864 107
rect 848 -30 864 102
rect 1352 407 1368 602
rect 1357 402 1362 407
rect 1367 402 1368 407
rect 1352 207 1368 402
rect 1357 202 1362 207
rect 1367 202 1368 207
rect 1352 7 1368 202
rect 1357 2 1362 7
rect 1367 2 1368 7
rect 1352 -30 1368 2
rect 1872 507 1888 702
rect 1877 502 1882 507
rect 1887 502 1888 507
rect 1872 307 1888 502
rect 1877 302 1882 307
rect 1887 302 1888 307
rect 1872 107 1888 302
rect 1965 922 1970 1797
rect 2013 1482 2018 2457
rect 2045 2312 2050 2477
rect 2061 1902 2066 2607
rect 1965 442 1970 917
rect 2029 562 2034 1777
rect 2061 1272 2066 1857
rect 2077 1622 2082 2647
rect 2109 2462 2114 2527
rect 2093 1382 2098 2437
rect 2125 2362 2130 3027
rect 2157 2872 2162 2917
rect 2173 2682 2178 3717
rect 2384 3607 2400 3802
rect 2389 3602 2394 3607
rect 2399 3602 2400 3607
rect 2253 3572 2258 3587
rect 2301 2792 2306 3487
rect 2384 3407 2400 3602
rect 2389 3402 2394 3407
rect 2399 3402 2400 3407
rect 2317 2792 2322 2857
rect 2141 2452 2146 2677
rect 2141 2437 2146 2447
rect 2157 2622 2162 2647
rect 2093 552 2098 1377
rect 2125 1112 2130 1937
rect 2141 1732 2146 2067
rect 2157 2012 2162 2617
rect 2157 1582 2162 2007
rect 2173 1562 2178 2307
rect 2189 2102 2194 2697
rect 2205 2412 2210 2427
rect 2253 1542 2258 2517
rect 2253 1192 2258 1537
rect 2269 1422 2274 2207
rect 2285 1712 2290 2737
rect 2301 2192 2306 2757
rect 2333 2202 2338 3307
rect 2384 3207 2400 3402
rect 2389 3202 2394 3207
rect 2399 3202 2400 3207
rect 2349 2842 2354 3077
rect 2384 3007 2400 3202
rect 2389 3002 2394 3007
rect 2399 3002 2400 3007
rect 2384 2807 2400 3002
rect 2389 2802 2394 2807
rect 2399 2802 2400 2807
rect 2384 2607 2400 2802
rect 2389 2602 2394 2607
rect 2399 2602 2400 2607
rect 2384 2407 2400 2602
rect 2389 2402 2394 2407
rect 2399 2402 2400 2407
rect 2384 2207 2400 2402
rect 2389 2202 2394 2207
rect 2399 2202 2400 2207
rect 2317 1452 2322 2147
rect 2317 962 2322 1447
rect 2384 2007 2400 2202
rect 2389 2002 2394 2007
rect 2399 2002 2400 2007
rect 2384 1807 2400 2002
rect 2389 1802 2394 1807
rect 2399 1802 2400 1807
rect 2384 1607 2400 1802
rect 2389 1602 2394 1607
rect 2399 1602 2400 1607
rect 2384 1407 2400 1602
rect 2389 1402 2394 1407
rect 2399 1402 2400 1407
rect 2384 1207 2400 1402
rect 2389 1202 2394 1207
rect 2399 1202 2400 1207
rect 2384 1007 2400 1202
rect 2413 1012 2418 3267
rect 2445 1252 2450 2277
rect 2461 1552 2466 2807
rect 2477 2462 2482 3507
rect 2493 3032 2498 3117
rect 2477 1572 2482 2267
rect 2509 1882 2514 2417
rect 2509 1352 2514 1367
rect 2525 1362 2530 2457
rect 2557 2422 2562 2997
rect 2573 2552 2578 4257
rect 2669 3022 2674 3057
rect 2685 2992 2690 3997
rect 2589 2092 2594 2727
rect 2541 1342 2546 1947
rect 2605 1702 2610 2687
rect 2621 2432 2626 2597
rect 2637 2582 2642 2927
rect 2637 1202 2642 2567
rect 2669 2382 2674 2807
rect 2669 2252 2674 2267
rect 2685 2252 2690 2927
rect 2701 2412 2706 3697
rect 2733 2932 2738 2947
rect 2749 2712 2754 4457
rect 2888 4307 2904 4502
rect 2893 4302 2898 4307
rect 2903 4302 2904 4307
rect 2888 4107 2904 4302
rect 3400 5007 3416 5130
rect 3405 5002 3410 5007
rect 3415 5002 3416 5007
rect 3400 4807 3416 5002
rect 3405 4802 3410 4807
rect 3415 4802 3416 4807
rect 3400 4607 3416 4802
rect 3405 4602 3410 4607
rect 3415 4602 3416 4607
rect 3400 4407 3416 4602
rect 3405 4402 3410 4407
rect 3415 4402 3416 4407
rect 3400 4207 3416 4402
rect 3920 5107 3936 5130
rect 3925 5102 3930 5107
rect 3935 5102 3936 5107
rect 3920 4907 3936 5102
rect 3925 4902 3930 4907
rect 3935 4902 3936 4907
rect 3920 4707 3936 4902
rect 3925 4702 3930 4707
rect 3935 4702 3936 4707
rect 3920 4507 3936 4702
rect 3925 4502 3930 4507
rect 3935 4502 3936 4507
rect 3920 4307 3936 4502
rect 4424 5007 4440 5130
rect 4936 5107 4952 5130
rect 4941 5102 4946 5107
rect 4951 5102 4952 5107
rect 4429 5002 4434 5007
rect 4439 5002 4440 5007
rect 4424 4807 4440 5002
rect 4429 4802 4434 4807
rect 4439 4802 4440 4807
rect 4424 4607 4440 4802
rect 4429 4602 4434 4607
rect 4439 4602 4440 4607
rect 4424 4407 4440 4602
rect 4429 4402 4434 4407
rect 4439 4402 4440 4407
rect 3925 4302 3930 4307
rect 3935 4302 3936 4307
rect 3405 4202 3410 4207
rect 3415 4202 3416 4207
rect 2893 4102 2898 4107
rect 2903 4102 2904 4107
rect 2888 3907 2904 4102
rect 2893 3902 2898 3907
rect 2903 3902 2904 3907
rect 2765 2302 2770 2767
rect 2781 2142 2786 3257
rect 2797 2762 2802 3647
rect 2877 3292 2882 3727
rect 2797 2342 2802 2377
rect 2389 1002 2394 1007
rect 2399 1002 2400 1007
rect 2384 807 2400 1002
rect 2389 802 2394 807
rect 2399 802 2400 807
rect 2384 607 2400 802
rect 2389 602 2394 607
rect 2399 602 2400 607
rect 1965 272 1970 437
rect 2384 407 2400 602
rect 2389 402 2394 407
rect 2399 402 2400 407
rect 1965 267 1973 272
rect 1877 102 1882 107
rect 1887 102 1888 107
rect 1872 -30 1888 102
rect 2384 207 2400 402
rect 2637 382 2642 1197
rect 2781 1142 2786 1927
rect 2813 1762 2818 2827
rect 2829 2392 2834 2667
rect 2845 1972 2850 2967
rect 2877 2952 2882 3287
rect 2888 3707 2904 3902
rect 3037 4112 3042 4157
rect 2893 3702 2898 3707
rect 2903 3702 2904 3707
rect 2888 3507 2904 3702
rect 2893 3502 2898 3507
rect 2903 3502 2904 3507
rect 2888 3307 2904 3502
rect 2893 3302 2898 3307
rect 2903 3302 2904 3307
rect 2888 3107 2904 3302
rect 2893 3102 2898 3107
rect 2903 3102 2904 3107
rect 2888 2907 2904 3102
rect 2893 2902 2898 2907
rect 2903 2902 2904 2907
rect 2888 2707 2904 2902
rect 2925 3352 2930 3777
rect 2925 2772 2930 3347
rect 2893 2702 2898 2707
rect 2903 2702 2904 2707
rect 2861 2482 2866 2537
rect 2888 2507 2904 2702
rect 2893 2502 2898 2507
rect 2903 2502 2904 2507
rect 2888 2307 2904 2502
rect 2893 2302 2898 2307
rect 2903 2302 2904 2307
rect 2888 2107 2904 2302
rect 2893 2102 2898 2107
rect 2903 2102 2904 2107
rect 2888 1907 2904 2102
rect 2893 1902 2898 1907
rect 2903 1902 2904 1907
rect 2781 932 2786 1137
rect 2888 1707 2904 1902
rect 2893 1702 2898 1707
rect 2903 1702 2904 1707
rect 2888 1507 2904 1702
rect 2893 1502 2898 1507
rect 2903 1502 2904 1507
rect 2888 1307 2904 1502
rect 2893 1302 2898 1307
rect 2903 1302 2904 1307
rect 2888 1107 2904 1302
rect 2909 1282 2914 1307
rect 2893 1102 2898 1107
rect 2903 1102 2904 1107
rect 2888 907 2904 1102
rect 2893 902 2898 907
rect 2903 902 2904 907
rect 2888 707 2904 902
rect 2925 892 2930 2527
rect 2973 2072 2978 3847
rect 3037 3152 3042 4107
rect 2973 912 2978 2067
rect 2989 1532 2994 2627
rect 3005 1972 3010 2477
rect 3021 1602 3026 2627
rect 3037 2492 3042 3127
rect 3037 2412 3042 2457
rect 3037 2332 3042 2367
rect 2989 862 2994 1527
rect 3053 1442 3058 2967
rect 3101 2542 3106 3527
rect 3165 2762 3170 3647
rect 3149 762 3154 2697
rect 3197 2482 3202 3827
rect 3213 2492 3218 3537
rect 3197 2382 3202 2397
rect 3229 1702 3234 2627
rect 3261 2232 3266 4007
rect 3400 4007 3416 4202
rect 3405 4002 3410 4007
rect 3415 4002 3416 4007
rect 3400 3807 3416 4002
rect 3405 3802 3410 3807
rect 3415 3802 3416 3807
rect 3309 3452 3314 3667
rect 3277 2192 3282 2277
rect 3261 1152 3266 1947
rect 3293 1942 3298 3277
rect 3309 2692 3314 3447
rect 3400 3607 3416 3802
rect 3405 3602 3410 3607
rect 3415 3602 3416 3607
rect 3400 3407 3416 3602
rect 3405 3402 3410 3407
rect 3415 3402 3416 3407
rect 3400 3207 3416 3402
rect 3405 3202 3410 3207
rect 3415 3202 3416 3207
rect 3293 1462 3298 1907
rect 3309 1232 3314 2527
rect 3325 2212 3330 2377
rect 3341 1362 3346 3007
rect 3400 3007 3416 3202
rect 3405 3002 3410 3007
rect 3415 3002 3416 3007
rect 3400 2807 3416 3002
rect 3405 2802 3410 2807
rect 3415 2802 3416 2807
rect 3400 2607 3416 2802
rect 3405 2602 3410 2607
rect 3415 2602 3416 2607
rect 3357 1572 3362 2517
rect 3357 1372 3362 1567
rect 3309 1152 3314 1227
rect 3373 1192 3378 2527
rect 3400 2407 3416 2602
rect 3405 2402 3410 2407
rect 3415 2402 3416 2407
rect 3400 2207 3416 2402
rect 3405 2202 3410 2207
rect 3415 2202 3416 2207
rect 3400 2007 3416 2202
rect 3405 2002 3410 2007
rect 3415 2002 3416 2007
rect 3400 1807 3416 2002
rect 3405 1802 3410 1807
rect 3415 1802 3416 1807
rect 3400 1607 3416 1802
rect 3405 1602 3410 1607
rect 3415 1602 3416 1607
rect 3400 1407 3416 1602
rect 3405 1402 3410 1407
rect 3415 1402 3416 1407
rect 3400 1207 3416 1402
rect 3405 1202 3410 1207
rect 3415 1202 3416 1207
rect 3400 1007 3416 1202
rect 3405 1002 3410 1007
rect 3415 1002 3416 1007
rect 3400 807 3416 1002
rect 3405 802 3410 807
rect 3415 802 3416 807
rect 2893 702 2898 707
rect 2903 702 2904 707
rect 2888 507 2904 702
rect 2893 502 2898 507
rect 2903 502 2904 507
rect 2389 202 2394 207
rect 2399 202 2400 207
rect 2384 7 2400 202
rect 2389 2 2394 7
rect 2399 2 2400 7
rect 2384 -30 2400 2
rect 2888 307 2904 502
rect 2893 302 2898 307
rect 2903 302 2904 307
rect 2888 107 2904 302
rect 2893 102 2898 107
rect 2903 102 2904 107
rect 2888 -30 2904 102
rect 3400 607 3416 802
rect 3453 682 3458 2767
rect 3485 2612 3490 3937
rect 3533 1582 3538 2637
rect 3549 2512 3554 4247
rect 3920 4107 3936 4302
rect 3925 4102 3930 4107
rect 3935 4102 3936 4107
rect 3920 3907 3936 4102
rect 3925 3902 3930 3907
rect 3935 3902 3936 3907
rect 3920 3707 3936 3902
rect 3925 3702 3930 3707
rect 3935 3702 3936 3707
rect 3901 3672 3906 3687
rect 3920 3507 3936 3702
rect 3925 3502 3930 3507
rect 3935 3502 3936 3507
rect 3920 3307 3936 3502
rect 3925 3302 3930 3307
rect 3935 3302 3936 3307
rect 3565 2832 3570 2877
rect 3565 2742 3570 2767
rect 3597 1372 3602 2057
rect 3629 1752 3634 2867
rect 3645 1472 3650 2687
rect 3805 1542 3810 2777
rect 3853 1812 3858 2237
rect 3885 2102 3890 3217
rect 3920 3107 3936 3302
rect 3925 3102 3930 3107
rect 3935 3102 3936 3107
rect 3920 2907 3936 3102
rect 3925 2902 3930 2907
rect 3935 2902 3936 2907
rect 3920 2707 3936 2902
rect 3925 2702 3930 2707
rect 3935 2702 3936 2707
rect 3920 2507 3936 2702
rect 3925 2502 3930 2507
rect 3935 2502 3936 2507
rect 3920 2307 3936 2502
rect 3925 2302 3930 2307
rect 3935 2302 3936 2307
rect 3920 2107 3936 2302
rect 3925 2102 3930 2107
rect 3935 2102 3936 2107
rect 3920 1907 3936 2102
rect 3925 1902 3930 1907
rect 3935 1902 3936 1907
rect 3920 1707 3936 1902
rect 3925 1702 3930 1707
rect 3935 1702 3936 1707
rect 3920 1507 3936 1702
rect 3925 1502 3930 1507
rect 3935 1502 3936 1507
rect 3920 1307 3936 1502
rect 3925 1302 3930 1307
rect 3935 1302 3936 1307
rect 3805 1262 3810 1297
rect 3920 1107 3936 1302
rect 3925 1102 3930 1107
rect 3935 1102 3936 1107
rect 3920 907 3936 1102
rect 3925 902 3930 907
rect 3935 902 3936 907
rect 3920 707 3936 902
rect 3925 702 3930 707
rect 3935 702 3936 707
rect 3405 602 3410 607
rect 3415 602 3416 607
rect 3400 407 3416 602
rect 3405 402 3410 407
rect 3415 402 3416 407
rect 3400 207 3416 402
rect 3405 202 3410 207
rect 3415 202 3416 207
rect 3400 7 3416 202
rect 3405 2 3410 7
rect 3415 2 3416 7
rect 3400 -30 3416 2
rect 3920 507 3936 702
rect 3925 502 3930 507
rect 3935 502 3936 507
rect 3920 307 3936 502
rect 3981 362 3986 1377
rect 3925 302 3930 307
rect 3935 302 3936 307
rect 3920 107 3936 302
rect 3997 282 4002 3377
rect 4045 1332 4050 2237
rect 4061 1762 4066 3047
rect 4093 652 4098 4357
rect 4424 4207 4440 4402
rect 4429 4202 4434 4207
rect 4439 4202 4440 4207
rect 4424 4007 4440 4202
rect 4429 4002 4434 4007
rect 4439 4002 4440 4007
rect 4424 3807 4440 4002
rect 4429 3802 4434 3807
rect 4439 3802 4440 3807
rect 4157 2162 4162 3617
rect 4424 3607 4440 3802
rect 4429 3602 4434 3607
rect 4439 3602 4440 3607
rect 4157 2072 4162 2157
rect 4173 1182 4178 3467
rect 4189 1052 4194 2947
rect 4205 1352 4210 3417
rect 4424 3407 4440 3602
rect 4429 3402 4434 3407
rect 4439 3402 4440 3407
rect 4424 3207 4440 3402
rect 4429 3202 4434 3207
rect 4439 3202 4440 3207
rect 4253 2447 4261 2452
rect 4253 1542 4258 2447
rect 4349 2027 4357 2032
rect 4205 572 4210 1347
rect 4349 1252 4354 2027
rect 4381 1572 4386 2627
rect 4365 1042 4370 1517
rect 4397 1512 4402 2677
rect 4413 1482 4418 3127
rect 4424 3007 4440 3202
rect 4429 3002 4434 3007
rect 4439 3002 4440 3007
rect 4424 2807 4440 3002
rect 4429 2802 4434 2807
rect 4439 2802 4440 2807
rect 4424 2607 4440 2802
rect 4429 2602 4434 2607
rect 4439 2602 4440 2607
rect 4424 2407 4440 2602
rect 4429 2402 4434 2407
rect 4439 2402 4440 2407
rect 4424 2207 4440 2402
rect 4429 2202 4434 2207
rect 4439 2202 4440 2207
rect 4424 2007 4440 2202
rect 4429 2002 4434 2007
rect 4439 2002 4440 2007
rect 4424 1807 4440 2002
rect 4477 1962 4482 3287
rect 4493 2872 4498 3977
rect 4509 2672 4514 5067
rect 4525 2842 4530 4127
rect 4541 3152 4546 5077
rect 4429 1802 4434 1807
rect 4439 1802 4440 1807
rect 4424 1607 4440 1802
rect 4493 1782 4498 2577
rect 4429 1602 4434 1607
rect 4439 1602 4440 1607
rect 4424 1407 4440 1602
rect 4525 1422 4530 2837
rect 4429 1402 4434 1407
rect 4439 1402 4440 1407
rect 4424 1207 4440 1402
rect 4429 1202 4434 1207
rect 4439 1202 4440 1207
rect 4424 1007 4440 1202
rect 4429 1002 4434 1007
rect 4439 1002 4440 1007
rect 4424 807 4440 1002
rect 4429 802 4434 807
rect 4439 802 4440 807
rect 4424 607 4440 802
rect 4429 602 4434 607
rect 4439 602 4440 607
rect 4424 407 4440 602
rect 4557 552 4562 1817
rect 4573 1572 4578 3327
rect 4589 1812 4594 4017
rect 4605 2032 4610 3227
rect 4621 892 4626 5057
rect 4653 4172 4658 4247
rect 4653 1942 4658 4167
rect 4429 402 4434 407
rect 4439 402 4440 407
rect 3925 102 3930 107
rect 3935 102 3936 107
rect 3920 -30 3936 102
rect 4424 207 4440 402
rect 4429 202 4434 207
rect 4439 202 4440 207
rect 4424 7 4440 202
rect 4669 82 4674 3637
rect 4685 762 4690 3957
rect 4701 2062 4706 3757
rect 4717 1372 4722 2257
rect 4733 1522 4738 2657
rect 4765 1922 4770 3467
rect 4813 2932 4818 4857
rect 4797 292 4802 2677
rect 4813 652 4818 2767
rect 4829 1132 4834 4717
rect 4845 2442 4850 5017
rect 4861 1472 4866 4337
rect 4877 262 4882 3497
rect 4893 2622 4898 3087
rect 4909 2642 4914 5047
rect 4925 2742 4930 5057
rect 4936 4907 4952 5102
rect 4941 4902 4946 4907
rect 4951 4902 4952 4907
rect 4936 4707 4952 4902
rect 4941 4702 4946 4707
rect 4951 4702 4952 4707
rect 4936 4507 4952 4702
rect 4941 4502 4946 4507
rect 4951 4502 4952 4507
rect 4936 4307 4952 4502
rect 4941 4302 4946 4307
rect 4951 4302 4952 4307
rect 4936 4107 4952 4302
rect 4941 4102 4946 4107
rect 4951 4102 4952 4107
rect 4936 3907 4952 4102
rect 4941 3902 4946 3907
rect 4951 3902 4952 3907
rect 4936 3707 4952 3902
rect 4941 3702 4946 3707
rect 4951 3702 4952 3707
rect 4936 3507 4952 3702
rect 4941 3502 4946 3507
rect 4951 3502 4952 3507
rect 4936 3307 4952 3502
rect 4941 3302 4946 3307
rect 4951 3302 4952 3307
rect 4936 3107 4952 3302
rect 4957 3192 4962 4467
rect 4973 3842 4978 4557
rect 4989 3852 4994 4537
rect 4941 3102 4946 3107
rect 4951 3102 4952 3107
rect 4936 2907 4952 3102
rect 4941 2902 4946 2907
rect 4951 2902 4952 2907
rect 4936 2707 4952 2902
rect 4941 2702 4946 2707
rect 4951 2702 4952 2707
rect 4936 2507 4952 2702
rect 4941 2502 4946 2507
rect 4951 2502 4952 2507
rect 4925 1072 4930 2377
rect 4936 2307 4952 2502
rect 4941 2302 4946 2307
rect 4951 2302 4952 2307
rect 4936 2107 4952 2302
rect 4941 2102 4946 2107
rect 4951 2102 4952 2107
rect 4936 1907 4952 2102
rect 4941 1902 4946 1907
rect 4951 1902 4952 1907
rect 4936 1707 4952 1902
rect 4941 1702 4946 1707
rect 4951 1702 4952 1707
rect 4936 1507 4952 1702
rect 4941 1502 4946 1507
rect 4951 1502 4952 1507
rect 4936 1307 4952 1502
rect 4941 1302 4946 1307
rect 4951 1302 4952 1307
rect 4936 1107 4952 1302
rect 4941 1102 4946 1107
rect 4951 1102 4952 1107
rect 4936 907 4952 1102
rect 4941 902 4946 907
rect 4951 902 4952 907
rect 4936 707 4952 902
rect 4957 772 4962 2957
rect 4941 702 4946 707
rect 4951 702 4952 707
rect 4936 507 4952 702
rect 4941 502 4946 507
rect 4951 502 4952 507
rect 4936 307 4952 502
rect 4941 302 4946 307
rect 4951 302 4952 307
rect 4936 107 4952 302
rect 4973 122 4978 3677
rect 4989 3392 4994 3837
rect 5005 3722 5010 4867
rect 5021 3972 5026 4587
rect 5037 3942 5042 4827
rect 4989 1432 4994 3367
rect 5005 2662 5010 3687
rect 5021 3002 5026 3507
rect 5037 3182 5042 3697
rect 5005 682 5010 2627
rect 5021 572 5026 2757
rect 5037 2702 5042 3167
rect 5037 1432 5042 2687
rect 5053 1902 5058 4267
rect 5037 272 5042 1227
rect 5069 972 5074 4927
rect 5085 2812 5090 4787
rect 5101 3562 5106 4287
rect 5085 1692 5090 2707
rect 5085 202 5090 1117
rect 5101 742 5106 3207
rect 5117 1862 5122 3997
rect 5133 3712 5138 4637
rect 5149 3932 5154 3997
rect 5133 1642 5138 3687
rect 5149 2982 5154 3717
rect 5165 3692 5170 4537
rect 4941 102 4946 107
rect 4951 102 4952 107
rect 4429 2 4434 7
rect 4439 2 4440 7
rect 4424 -30 4440 2
rect 4936 -30 4952 102
rect 5133 62 5138 1427
rect 5149 92 5154 2957
rect 5165 2502 5170 3557
rect 5165 1142 5170 2487
rect 5181 2132 5186 3867
rect 5197 2912 5202 4457
rect 5213 3192 5218 4117
rect 5197 2172 5202 2857
rect 5181 872 5186 1727
rect 5197 472 5202 2167
rect 5213 2142 5218 3167
rect 5229 2842 5234 3857
rect 5213 1182 5218 2127
rect 5229 2112 5234 2827
rect 5245 2572 5250 4697
rect 5245 2102 5250 2547
rect 5229 452 5234 2067
rect 5245 152 5250 1957
rect 5261 1862 5266 4077
rect 5277 3162 5282 4307
rect 5277 2232 5282 3127
rect 5293 1922 5298 3257
rect 5261 132 5266 1637
rect 5277 992 5282 1157
rect 5293 152 5298 977
use DFFPOSX1  DFFPOSX1_1027
timestamp 1607101874
transform -1 0 100 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_141
timestamp 1607101874
transform 1 0 100 0 -1 105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_57
timestamp 1607101874
transform 1 0 4 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_548
timestamp 1607101874
transform 1 0 76 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_128
timestamp 1607101874
transform -1 0 164 0 -1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_46
timestamp 1607101874
transform 1 0 164 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_87
timestamp 1607101874
transform -1 0 220 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1607101874
transform 1 0 172 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_735
timestamp 1607101874
transform 1 0 220 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_521
timestamp 1607101874
transform 1 0 268 0 1 105
box -2 -3 98 103
use FILL  FILL_0_0_0
timestamp 1607101874
transform 1 0 316 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1607101874
transform 1 0 324 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1031
timestamp 1607101874
transform 1 0 332 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_0_0
timestamp 1607101874
transform 1 0 364 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1607101874
transform 1 0 372 0 1 105
box -2 -3 10 103
use INVX1  INVX1_384
timestamp 1607101874
transform 1 0 380 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_148
timestamp 1607101874
transform 1 0 396 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_520
timestamp 1607101874
transform 1 0 428 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_235
timestamp 1607101874
transform -1 0 452 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_34
timestamp 1607101874
transform 1 0 452 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1030
timestamp 1607101874
transform 1 0 524 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_321
timestamp 1607101874
transform 1 0 524 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_151
timestamp 1607101874
transform 1 0 540 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_238
timestamp 1607101874
transform -1 0 596 0 1 105
box -2 -3 26 103
use INVX1  INVX1_142
timestamp 1607101874
transform 1 0 596 0 1 105
box -2 -3 18 103
use INVX1  INVX1_144
timestamp 1607101874
transform 1 0 620 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_131
timestamp 1607101874
transform 1 0 636 0 -1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_301
timestamp 1607101874
transform 1 0 684 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1028
timestamp 1607101874
transform -1 0 708 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_663
timestamp 1607101874
transform 1 0 708 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_737
timestamp 1607101874
transform -1 0 812 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_93
timestamp 1607101874
transform 1 0 740 0 1 105
box -2 -3 74 103
use AOI21X1  AOI21X1_440
timestamp 1607101874
transform 1 0 812 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_0
timestamp 1607101874
transform 1 0 844 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1607101874
transform 1 0 852 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_88
timestamp 1607101874
transform 1 0 860 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_47
timestamp 1607101874
transform -1 0 916 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1607101874
transform 1 0 812 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1607101874
transform 1 0 820 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1607101874
transform 1 0 828 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_874
timestamp 1607101874
transform 1 0 916 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_88
timestamp 1607101874
transform 1 0 1012 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_869
timestamp 1607101874
transform 1 0 924 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_148
timestamp 1607101874
transform -1 0 1068 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1607101874
transform 1 0 1068 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_106
timestamp 1607101874
transform 1 0 1020 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_93
timestamp 1607101874
transform -1 0 1084 0 1 105
box -2 -3 50 103
use NOR2X1  NOR2X1_599
timestamp 1607101874
transform 1 0 1084 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_861
timestamp 1607101874
transform 1 0 1108 0 1 105
box -2 -3 98 103
use INVX1  INVX1_314
timestamp 1607101874
transform 1 0 1164 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_335
timestamp 1607101874
transform 1 0 1180 0 -1 105
box -2 -3 50 103
use INVX1  INVX1_104
timestamp 1607101874
transform 1 0 1204 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_870
timestamp 1607101874
transform 1 0 1228 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_85
timestamp 1607101874
transform 1 0 1220 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_144
timestamp 1607101874
transform -1 0 1276 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_26
timestamp 1607101874
transform 1 0 1276 0 1 105
box -2 -3 74 103
use AOI21X1  AOI21X1_337
timestamp 1607101874
transform 1 0 1324 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1607101874
transform 1 0 1356 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1607101874
transform 1 0 1364 0 -1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_336
timestamp 1607101874
transform 1 0 1372 0 -1 105
box -2 -3 50 103
use FILL  FILL_1_2_0
timestamp 1607101874
transform 1 0 1348 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1607101874
transform 1 0 1356 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1607101874
transform 1 0 1364 0 1 105
box -2 -3 98 103
use INVX1  INVX1_355
timestamp 1607101874
transform -1 0 1436 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1607101874
transform -1 0 1532 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_567
timestamp 1607101874
transform 1 0 1460 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_679
timestamp 1607101874
transform -1 0 1516 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_767
timestamp 1607101874
transform -1 0 1548 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1607101874
transform 1 0 1532 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1607101874
transform 1 0 1548 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_561
timestamp 1607101874
transform 1 0 1628 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_673
timestamp 1607101874
transform 1 0 1660 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_278
timestamp 1607101874
transform -1 0 1780 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_354
timestamp 1607101874
transform 1 0 1644 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_333
timestamp 1607101874
transform -1 0 1708 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1607101874
transform -1 0 1804 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_280
timestamp 1607101874
transform 1 0 1780 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_247
timestamp 1607101874
transform 1 0 1804 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_334
timestamp 1607101874
transform 1 0 1820 0 1 105
box -2 -3 50 103
use FILL  FILL_0_3_0
timestamp 1607101874
transform -1 0 1884 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1607101874
transform -1 0 1892 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_678
timestamp 1607101874
transform -1 0 1916 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_855
timestamp 1607101874
transform 1 0 1916 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_3_0
timestamp 1607101874
transform 1 0 1868 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1607101874
transform 1 0 1876 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_566
timestamp 1607101874
transform 1 0 1884 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1607101874
transform 1 0 1916 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1607101874
transform 1 0 2012 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_352
timestamp 1607101874
transform 1 0 2012 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_34
timestamp 1607101874
transform -1 0 2156 0 -1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_330
timestamp 1607101874
transform 1 0 2028 0 1 105
box -2 -3 50 103
use INVX1  INVX1_244
timestamp 1607101874
transform 1 0 2076 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_329
timestamp 1607101874
transform -1 0 2140 0 1 105
box -2 -3 50 103
use INVX1  INVX1_42
timestamp 1607101874
transform -1 0 2172 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_689
timestamp 1607101874
transform -1 0 2268 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_281
timestamp 1607101874
transform 1 0 2140 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_398
timestamp 1607101874
transform 1 0 2268 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_422
timestamp 1607101874
transform 1 0 2236 0 1 105
box -2 -3 18 103
use INVX1  INVX1_246
timestamp 1607101874
transform 1 0 2252 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_332
timestamp 1607101874
transform 1 0 2268 0 1 105
box -2 -3 50 103
use NOR2X1  NOR2X1_136
timestamp 1607101874
transform 1 0 2316 0 1 105
box -2 -3 26 103
use FILL  FILL_0_4_0
timestamp 1607101874
transform 1 0 2364 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_4_1
timestamp 1607101874
transform 1 0 2372 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_688
timestamp 1607101874
transform 1 0 2380 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_79
timestamp 1607101874
transform -1 0 2372 0 1 105
box -2 -3 34 103
use FILL  FILL_1_4_0
timestamp 1607101874
transform -1 0 2380 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_1
timestamp 1607101874
transform -1 0 2388 0 1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_69
timestamp 1607101874
transform -1 0 2460 0 1 105
box -2 -3 74 103
use INVX1  INVX1_41
timestamp 1607101874
transform 1 0 2476 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_33
timestamp 1607101874
transform 1 0 2492 0 -1 105
box -2 -3 50 103
use CLKBUF1  CLKBUF1_70
timestamp 1607101874
transform 1 0 2460 0 1 105
box -2 -3 74 103
use AOI21X1  AOI21X1_29
timestamp 1607101874
transform 1 0 2540 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1607101874
transform -1 0 2596 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_696
timestamp 1607101874
transform -1 0 2692 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_441
timestamp 1607101874
transform 1 0 2532 0 1 105
box -2 -3 98 103
use INVX1  INVX1_361
timestamp 1607101874
transform 1 0 2628 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_687
timestamp 1607101874
transform 1 0 2692 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_271
timestamp 1607101874
transform 1 0 2644 0 1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_514
timestamp 1607101874
transform 1 0 2692 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_626
timestamp 1607101874
transform 1 0 2724 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_396
timestamp 1607101874
transform 1 0 2788 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_691
timestamp 1607101874
transform -1 0 2844 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_55
timestamp 1607101874
transform -1 0 2908 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_5_0
timestamp 1607101874
transform 1 0 2908 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1607101874
transform 1 0 2916 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_439
timestamp 1607101874
transform 1 0 2924 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_26
timestamp 1607101874
transform 1 0 2844 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1607101874
transform 1 0 2876 0 1 105
box -2 -3 26 103
use FILL  FILL_1_5_0
timestamp 1607101874
transform -1 0 2908 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_1
timestamp 1607101874
transform -1 0 2916 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_24
timestamp 1607101874
transform -1 0 2948 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1607101874
transform 1 0 3020 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_692
timestamp 1607101874
transform 1 0 2948 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_440
timestamp 1607101874
transform -1 0 3212 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_43
timestamp 1607101874
transform 1 0 3044 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_35
timestamp 1607101874
transform 1 0 3060 0 1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_515
timestamp 1607101874
transform 1 0 3108 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_630
timestamp 1607101874
transform -1 0 3236 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_627
timestamp 1607101874
transform 1 0 3140 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_43
timestamp 1607101874
transform 1 0 3164 0 1 105
box -2 -3 74 103
use AOI21X1  AOI21X1_518
timestamp 1607101874
transform -1 0 3268 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_695
timestamp 1607101874
transform 1 0 3268 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_94
timestamp 1607101874
transform 1 0 3236 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1607101874
transform 1 0 3308 0 1 105
box -2 -3 98 103
use FILL  FILL_0_6_0
timestamp 1607101874
transform 1 0 3364 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_6_1
timestamp 1607101874
transform 1 0 3372 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_397
timestamp 1607101874
transform 1 0 3380 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_6_0
timestamp 1607101874
transform 1 0 3404 0 1 105
box -2 -3 10 103
use FILL  FILL_1_6_1
timestamp 1607101874
transform 1 0 3412 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_517
timestamp 1607101874
transform 1 0 3420 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_711
timestamp 1607101874
transform -1 0 3572 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_629
timestamp 1607101874
transform 1 0 3452 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_513
timestamp 1607101874
transform 1 0 3476 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_625
timestamp 1607101874
transform -1 0 3532 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_401
timestamp 1607101874
transform 1 0 3532 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1607101874
transform 1 0 3572 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_72
timestamp 1607101874
transform -1 0 3628 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_714
timestamp 1607101874
transform 1 0 3628 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_699
timestamp 1607101874
transform 1 0 3556 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_61
timestamp 1607101874
transform 1 0 3588 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_28
timestamp 1607101874
transform -1 0 3644 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_33
timestamp 1607101874
transform 1 0 3724 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_554
timestamp 1607101874
transform 1 0 3644 0 1 105
box -2 -3 34 103
use INVX1  INVX1_304
timestamp 1607101874
transform 1 0 3676 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_267
timestamp 1607101874
transform 1 0 3692 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_702
timestamp 1607101874
transform -1 0 3836 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_67
timestamp 1607101874
transform -1 0 3780 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_704
timestamp 1607101874
transform 1 0 3780 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_823
timestamp 1607101874
transform -1 0 3868 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_179
timestamp 1607101874
transform 1 0 3876 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_276
timestamp 1607101874
transform -1 0 3932 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_7_0
timestamp 1607101874
transform -1 0 3940 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_7_1
timestamp 1607101874
transform -1 0 3948 0 -1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_36
timestamp 1607101874
transform 1 0 3868 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_71
timestamp 1607101874
transform 1 0 3900 0 1 105
box -2 -3 26 103
use FILL  FILL_1_7_0
timestamp 1607101874
transform 1 0 3924 0 1 105
box -2 -3 10 103
use FILL  FILL_1_7_1
timestamp 1607101874
transform 1 0 3932 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1607101874
transform 1 0 3940 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1607101874
transform -1 0 4044 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_176
timestamp 1607101874
transform 1 0 4036 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_163
timestamp 1607101874
transform -1 0 4092 0 -1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_187
timestamp 1607101874
transform 1 0 4092 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_284
timestamp 1607101874
transform -1 0 4148 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_303
timestamp 1607101874
transform 1 0 4052 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_273
timestamp 1607101874
transform -1 0 4116 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1607101874
transform 1 0 4116 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_646
timestamp 1607101874
transform 1 0 4148 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_11
timestamp 1607101874
transform -1 0 4276 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_24
timestamp 1607101874
transform -1 0 4284 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1607101874
transform 1 0 4276 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_31
timestamp 1607101874
transform 1 0 4284 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_80
timestamp 1607101874
transform 1 0 4308 0 1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_24
timestamp 1607101874
transform -1 0 4396 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1607101874
transform -1 0 4428 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_8_0
timestamp 1607101874
transform 1 0 4428 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_8_1
timestamp 1607101874
transform 1 0 4436 0 -1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_156
timestamp 1607101874
transform 1 0 4444 0 -1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_610
timestamp 1607101874
transform -1 0 4476 0 1 105
box -2 -3 98 103
use INVX1  INVX1_169
timestamp 1607101874
transform -1 0 4508 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1607101874
transform -1 0 4604 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_8_0
timestamp 1607101874
transform 1 0 4476 0 1 105
box -2 -3 10 103
use FILL  FILL_1_8_1
timestamp 1607101874
transform 1 0 4484 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1607101874
transform 1 0 4492 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_22
timestamp 1607101874
transform 1 0 4604 0 -1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_181
timestamp 1607101874
transform 1 0 4588 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_278
timestamp 1607101874
transform 1 0 4620 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_21
timestamp 1607101874
transform 1 0 4644 0 1 105
box -2 -3 74 103
use INVX1  INVX1_29
timestamp 1607101874
transform -1 0 4668 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_632
timestamp 1607101874
transform -1 0 4764 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_34
timestamp 1607101874
transform 1 0 4716 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1607101874
transform -1 0 4772 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1607101874
transform -1 0 4796 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1607101874
transform 1 0 4796 0 -1 105
box -2 -3 18 103
use INVX1  INVX1_171
timestamp 1607101874
transform -1 0 4828 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_338
timestamp 1607101874
transform -1 0 4924 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_651
timestamp 1607101874
transform -1 0 4868 0 1 105
box -2 -3 98 103
use FILL  FILL_0_9_0
timestamp 1607101874
transform -1 0 4932 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_9_1
timestamp 1607101874
transform -1 0 4940 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_653
timestamp 1607101874
transform -1 0 5036 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_636
timestamp 1607101874
transform 1 0 4868 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1607101874
transform 1 0 5036 0 -1 105
box -2 -3 74 103
use FILL  FILL_1_9_0
timestamp 1607101874
transform -1 0 4972 0 1 105
box -2 -3 10 103
use FILL  FILL_1_9_1
timestamp 1607101874
transform -1 0 4980 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_25
timestamp 1607101874
transform -1 0 5028 0 1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_24
timestamp 1607101874
transform 1 0 5028 0 1 105
box -2 -3 50 103
use CLKBUF1  CLKBUF1_84
timestamp 1607101874
transform 1 0 5108 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_634
timestamp 1607101874
transform -1 0 5172 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_5
timestamp 1607101874
transform 1 0 5180 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1607101874
transform 1 0 5204 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_30
timestamp 1607101874
transform 1 0 5172 0 1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_494
timestamp 1607101874
transform -1 0 5268 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1
timestamp 1607101874
transform -1 0 5308 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_109
timestamp 1607101874
transform -1 0 5292 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1607101874
transform 1 0 5292 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1607101874
transform 1 0 5300 0 1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_254
timestamp 1607101874
transform -1 0 28 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_163
timestamp 1607101874
transform -1 0 60 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_619
timestamp 1607101874
transform 1 0 60 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_731
timestamp 1607101874
transform -1 0 116 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1057
timestamp 1607101874
transform 1 0 116 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_531
timestamp 1607101874
transform 1 0 212 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_387
timestamp 1607101874
transform -1 0 292 0 -1 305
box -2 -3 50 103
use FILL  FILL_2_0_0
timestamp 1607101874
transform 1 0 292 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1607101874
transform 1 0 300 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_549
timestamp 1607101874
transform 1 0 308 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_386
timestamp 1607101874
transform -1 0 452 0 -1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_161
timestamp 1607101874
transform 1 0 452 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_252
timestamp 1607101874
transform -1 0 508 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1034
timestamp 1607101874
transform 1 0 508 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_129
timestamp 1607101874
transform 1 0 604 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_296
timestamp 1607101874
transform 1 0 652 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_457
timestamp 1607101874
transform 1 0 748 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_327
timestamp 1607101874
transform -1 0 812 0 -1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_532
timestamp 1607101874
transform 1 0 812 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1607101874
transform -1 0 852 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1607101874
transform -1 0 860 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_644
timestamp 1607101874
transform -1 0 884 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_299
timestamp 1607101874
transform -1 0 980 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_873
timestamp 1607101874
transform -1 0 1076 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_87
timestamp 1607101874
transform 1 0 1076 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_147
timestamp 1607101874
transform -1 0 1132 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_91
timestamp 1607101874
transform -1 0 1180 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_865
timestamp 1607101874
transform 1 0 1180 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_141
timestamp 1607101874
transform -1 0 1300 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1607101874
transform -1 0 1332 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_2_0
timestamp 1607101874
transform 1 0 1332 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1607101874
transform 1 0 1340 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_862
timestamp 1607101874
transform 1 0 1348 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1607101874
transform 1 0 1444 0 -1 305
box -2 -3 98 103
use BUFX4  BUFX4_329
timestamp 1607101874
transform -1 0 1572 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_568
timestamp 1607101874
transform 1 0 1572 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_680
timestamp 1607101874
transform -1 0 1628 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1607101874
transform 1 0 1628 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_569
timestamp 1607101874
transform -1 0 1756 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_681
timestamp 1607101874
transform -1 0 1780 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_399
timestamp 1607101874
transform 1 0 1780 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_924
timestamp 1607101874
transform -1 0 1844 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_3_0
timestamp 1607101874
transform -1 0 1852 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1607101874
transform -1 0 1860 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1607101874
transform -1 0 1956 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_176
timestamp 1607101874
transform 1 0 1956 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_671
timestamp 1607101874
transform -1 0 2004 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_559
timestamp 1607101874
transform -1 0 2036 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1607101874
transform 1 0 2036 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_372
timestamp 1607101874
transform -1 0 2156 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_547
timestamp 1607101874
transform 1 0 2156 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_331
timestamp 1607101874
transform -1 0 2228 0 -1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_268
timestamp 1607101874
transform 1 0 2228 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_397
timestamp 1607101874
transform -1 0 2284 0 -1 305
box -2 -3 26 103
use BUFX4  BUFX4_351
timestamp 1607101874
transform 1 0 2284 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_847
timestamp 1607101874
transform -1 0 2412 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_4_0
timestamp 1607101874
transform 1 0 2412 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1607101874
transform 1 0 2420 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1019
timestamp 1607101874
transform 1 0 2428 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_437
timestamp 1607101874
transform -1 0 2492 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_693
timestamp 1607101874
transform 1 0 2492 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_36
timestamp 1607101874
transform -1 0 2636 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_398
timestamp 1607101874
transform -1 0 2652 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_71
timestamp 1607101874
transform -1 0 2684 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_72
timestamp 1607101874
transform -1 0 2716 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1607101874
transform -1 0 2812 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_821
timestamp 1607101874
transform -1 0 2844 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_358
timestamp 1607101874
transform -1 0 2876 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_332
timestamp 1607101874
transform -1 0 2892 0 -1 305
box -2 -3 18 103
use FILL  FILL_2_5_0
timestamp 1607101874
transform 1 0 2892 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1607101874
transform 1 0 2900 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_519
timestamp 1607101874
transform 1 0 2908 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_631
timestamp 1607101874
transform -1 0 2964 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_442
timestamp 1607101874
transform 1 0 2964 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_69
timestamp 1607101874
transform 1 0 3060 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1607101874
transform -1 0 3124 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1607101874
transform -1 0 3220 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_68
timestamp 1607101874
transform 1 0 3220 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_67
timestamp 1607101874
transform 1 0 3252 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1265
timestamp 1607101874
transform 1 0 3284 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1266
timestamp 1607101874
transform -1 0 3348 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1607101874
transform 1 0 3348 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_6_0
timestamp 1607101874
transform 1 0 3444 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1607101874
transform 1 0 3452 0 -1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_269
timestamp 1607101874
transform 1 0 3460 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1607101874
transform 1 0 3508 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_222
timestamp 1607101874
transform 1 0 3604 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_743
timestamp 1607101874
transform 1 0 3620 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_170
timestamp 1607101874
transform -1 0 3676 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_742
timestamp 1607101874
transform 1 0 3676 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_575
timestamp 1607101874
transform 1 0 3708 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_327
timestamp 1607101874
transform -1 0 3764 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1607101874
transform -1 0 3796 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1607101874
transform -1 0 3828 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_77
timestamp 1607101874
transform 1 0 3828 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_78
timestamp 1607101874
transform -1 0 3892 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_7_0
timestamp 1607101874
transform -1 0 3900 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_7_1
timestamp 1607101874
transform -1 0 3908 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_700
timestamp 1607101874
transform -1 0 4004 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_69
timestamp 1607101874
transform -1 0 4028 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_35
timestamp 1607101874
transform -1 0 4060 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_706
timestamp 1607101874
transform -1 0 4156 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1274
timestamp 1607101874
transform -1 0 4188 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1273
timestamp 1607101874
transform 1 0 4188 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1607101874
transform 1 0 4220 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_223
timestamp 1607101874
transform 1 0 4316 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_250
timestamp 1607101874
transform 1 0 4332 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_556
timestamp 1607101874
transform 1 0 4364 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_864
timestamp 1607101874
transform 1 0 4396 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_8_0
timestamp 1607101874
transform 1 0 4428 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_8_1
timestamp 1607101874
transform 1 0 4436 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_17
timestamp 1607101874
transform 1 0 4444 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_12
timestamp 1607101874
transform -1 0 4508 0 -1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_381
timestamp 1607101874
transform 1 0 4508 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_98
timestamp 1607101874
transform 1 0 4540 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_179
timestamp 1607101874
transform 1 0 4564 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_388
timestamp 1607101874
transform 1 0 4580 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1607101874
transform -1 0 4708 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_285
timestamp 1607101874
transform 1 0 4708 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_452
timestamp 1607101874
transform 1 0 4732 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1053
timestamp 1607101874
transform 1 0 4764 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_152
timestamp 1607101874
transform 1 0 4796 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_165
timestamp 1607101874
transform -1 0 4860 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1607101874
transform -1 0 4956 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_9_0
timestamp 1607101874
transform -1 0 4964 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_9_1
timestamp 1607101874
transform -1 0 4972 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_480
timestamp 1607101874
transform -1 0 5004 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_709
timestamp 1607101874
transform 1 0 5004 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_33
timestamp 1607101874
transform -1 0 5044 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_652
timestamp 1607101874
transform 1 0 5044 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_355
timestamp 1607101874
transform 1 0 5140 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_342
timestamp 1607101874
transform 1 0 5172 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_191
timestamp 1607101874
transform 1 0 5188 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_2
timestamp 1607101874
transform 1 0 5220 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1607101874
transform -1 0 5276 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_177
timestamp 1607101874
transform -1 0 5292 0 -1 305
box -2 -3 18 103
use FILL  FILL_3_1
timestamp 1607101874
transform -1 0 5300 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1607101874
transform -1 0 5308 0 -1 305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_52
timestamp 1607101874
transform 1 0 4 0 1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1607101874
transform 1 0 76 0 1 305
box -2 -3 98 103
use INVX1  INVX1_145
timestamp 1607101874
transform 1 0 172 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_350
timestamp 1607101874
transform 1 0 188 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1607101874
transform -1 0 308 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_643
timestamp 1607101874
transform 1 0 308 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1607101874
transform 1 0 332 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1607101874
transform 1 0 340 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_162
timestamp 1607101874
transform 1 0 348 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_253
timestamp 1607101874
transform 1 0 380 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_620
timestamp 1607101874
transform 1 0 404 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_732
timestamp 1607101874
transform 1 0 436 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_553
timestamp 1607101874
transform 1 0 460 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1056
timestamp 1607101874
transform 1 0 556 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_294
timestamp 1607101874
transform 1 0 652 0 1 305
box -2 -3 98 103
use INVX1  INVX1_455
timestamp 1607101874
transform -1 0 764 0 1 305
box -2 -3 18 103
use INVX1  INVX1_251
timestamp 1607101874
transform -1 0 780 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_298
timestamp 1607101874
transform -1 0 876 0 1 305
box -2 -3 98 103
use FILL  FILL_3_1_0
timestamp 1607101874
transform 1 0 876 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1607101874
transform 1 0 884 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_349
timestamp 1607101874
transform 1 0 892 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_1256
timestamp 1607101874
transform -1 0 948 0 1 305
box -2 -3 34 103
use INVX1  INVX1_313
timestamp 1607101874
transform 1 0 948 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_322
timestamp 1607101874
transform -1 0 1012 0 1 305
box -2 -3 50 103
use CLKBUF1  CLKBUF1_32
timestamp 1607101874
transform 1 0 1012 0 1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_860
timestamp 1607101874
transform 1 0 1084 0 1 305
box -2 -3 98 103
use INVX1  INVX1_103
timestamp 1607101874
transform 1 0 1180 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_90
timestamp 1607101874
transform -1 0 1244 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_188
timestamp 1607101874
transform 1 0 1244 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_189
timestamp 1607101874
transform -1 0 1308 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_191
timestamp 1607101874
transform 1 0 1308 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_190
timestamp 1607101874
transform 1 0 1340 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1607101874
transform 1 0 1372 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1607101874
transform 1 0 1380 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_866
timestamp 1607101874
transform 1 0 1388 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1218
timestamp 1607101874
transform 1 0 1484 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_598
timestamp 1607101874
transform 1 0 1516 0 1 305
box -2 -3 26 103
use OAI22X1  OAI22X1_79
timestamp 1607101874
transform -1 0 1580 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_1219
timestamp 1607101874
transform 1 0 1580 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1384
timestamp 1607101874
transform 1 0 1612 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1385
timestamp 1607101874
transform -1 0 1676 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1607101874
transform 1 0 1676 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_278
timestamp 1607101874
transform -1 0 1796 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_925
timestamp 1607101874
transform 1 0 1796 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1386
timestamp 1607101874
transform 1 0 1828 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1607101874
transform -1 0 1868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1607101874
transform -1 0 1876 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_400
timestamp 1607101874
transform -1 0 1908 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1387
timestamp 1607101874
transform 1 0 1908 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1607101874
transform 1 0 1940 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_472
timestamp 1607101874
transform -1 0 2060 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_588
timestamp 1607101874
transform 1 0 2060 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_674
timestamp 1607101874
transform 1 0 2092 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_562
timestamp 1607101874
transform -1 0 2148 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_354
timestamp 1607101874
transform -1 0 2180 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_269
timestamp 1607101874
transform 1 0 2180 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_356
timestamp 1607101874
transform 1 0 2212 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_587
timestamp 1607101874
transform -1 0 2276 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1607101874
transform -1 0 2372 0 1 305
box -2 -3 98 103
use FILL  FILL_3_4_0
timestamp 1607101874
transform -1 0 2380 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1607101874
transform -1 0 2388 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1383
timestamp 1607101874
transform -1 0 2420 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_89
timestamp 1607101874
transform 1 0 2420 0 1 305
box -2 -3 50 103
use INVX1  INVX1_102
timestamp 1607101874
transform -1 0 2484 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_859
timestamp 1607101874
transform -1 0 2580 0 1 305
box -2 -3 98 103
use INVX1  INVX1_44
timestamp 1607101874
transform 1 0 2580 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_132
timestamp 1607101874
transform 1 0 2596 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_76
timestamp 1607101874
transform -1 0 2652 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_670
timestamp 1607101874
transform 1 0 2652 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_558
timestamp 1607101874
transform -1 0 2708 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_279
timestamp 1607101874
transform -1 0 2804 0 1 305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_31
timestamp 1607101874
transform -1 0 2876 0 1 305
box -2 -3 74 103
use FILL  FILL_3_5_0
timestamp 1607101874
transform 1 0 2876 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1607101874
transform 1 0 2884 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_575
timestamp 1607101874
transform 1 0 2892 0 1 305
box -2 -3 98 103
use INVX1  INVX1_270
timestamp 1607101874
transform -1 0 3004 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_521
timestamp 1607101874
transform -1 0 3028 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_700
timestamp 1607101874
transform 1 0 3028 0 1 305
box -2 -3 34 103
use INVX1  INVX1_328
timestamp 1607101874
transform -1 0 3076 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_576
timestamp 1607101874
transform -1 0 3172 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_268
timestamp 1607101874
transform -1 0 3220 0 1 305
box -2 -3 50 103
use INVX1  INVX1_412
timestamp 1607101874
transform -1 0 3236 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_399
timestamp 1607101874
transform -1 0 3332 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_709
timestamp 1607101874
transform -1 0 3428 0 1 305
box -2 -3 98 103
use FILL  FILL_3_6_0
timestamp 1607101874
transform 1 0 3428 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1607101874
transform 1 0 3436 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1607101874
transform 1 0 3444 0 1 305
box -2 -3 98 103
use OAI22X1  OAI22X1_16
timestamp 1607101874
transform 1 0 3540 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_400
timestamp 1607101874
transform 1 0 3580 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_363
timestamp 1607101874
transform 1 0 3604 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_364
timestamp 1607101874
transform 1 0 3628 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_555
timestamp 1607101874
transform -1 0 3684 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_744
timestamp 1607101874
transform 1 0 3684 0 1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_68
timestamp 1607101874
transform 1 0 3716 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_574
timestamp 1607101874
transform -1 0 3780 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_745
timestamp 1607101874
transform 1 0 3780 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_445
timestamp 1607101874
transform 1 0 3812 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_444
timestamp 1607101874
transform -1 0 3860 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_1183
timestamp 1607101874
transform -1 0 3892 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_352
timestamp 1607101874
transform -1 0 3924 0 1 305
box -2 -3 34 103
use FILL  FILL_3_7_0
timestamp 1607101874
transform -1 0 3932 0 1 305
box -2 -3 10 103
use FILL  FILL_3_7_1
timestamp 1607101874
transform -1 0 3940 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1607101874
transform -1 0 4036 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_699
timestamp 1607101874
transform -1 0 4132 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_76
timestamp 1607101874
transform 1 0 4132 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_75
timestamp 1607101874
transform -1 0 4196 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_272
timestamp 1607101874
transform 1 0 4196 0 1 305
box -2 -3 50 103
use INVX1  INVX1_224
timestamp 1607101874
transform -1 0 4260 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1607101874
transform 1 0 4260 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_632
timestamp 1607101874
transform -1 0 4380 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_520
timestamp 1607101874
transform -1 0 4412 0 1 305
box -2 -3 34 103
use FILL  FILL_3_8_0
timestamp 1607101874
transform 1 0 4412 0 1 305
box -2 -3 10 103
use FILL  FILL_3_8_1
timestamp 1607101874
transform 1 0 4420 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_382
timestamp 1607101874
transform 1 0 4428 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_865
timestamp 1607101874
transform -1 0 4556 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1607101874
transform -1 0 4652 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1040
timestamp 1607101874
transform 1 0 4652 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_188
timestamp 1607101874
transform 1 0 4684 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_349
timestamp 1607101874
transform 1 0 4716 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_326
timestamp 1607101874
transform 1 0 4748 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_630
timestamp 1607101874
transform 1 0 4780 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_4
timestamp 1607101874
transform 1 0 4876 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_20
timestamp 1607101874
transform -1 0 4932 0 1 305
box -2 -3 26 103
use FILL  FILL_3_9_0
timestamp 1607101874
transform 1 0 4932 0 1 305
box -2 -3 10 103
use FILL  FILL_3_9_1
timestamp 1607101874
transform 1 0 4940 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1141
timestamp 1607101874
transform 1 0 4948 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_184
timestamp 1607101874
transform 1 0 4980 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_281
timestamp 1607101874
transform -1 0 5036 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1607101874
transform -1 0 5132 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_813
timestamp 1607101874
transform 1 0 5132 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1607101874
transform -1 0 5196 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_288
timestamp 1607101874
transform -1 0 5220 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_812
timestamp 1607101874
transform -1 0 5252 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_178
timestamp 1607101874
transform 1 0 5252 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_506
timestamp 1607101874
transform -1 0 5308 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1607101874
transform 1 0 4 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_147
timestamp 1607101874
transform 1 0 100 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_132
timestamp 1607101874
transform -1 0 164 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_134
timestamp 1607101874
transform 1 0 164 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1055
timestamp 1607101874
transform 1 0 212 0 -1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_160
timestamp 1607101874
transform 1 0 308 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1607101874
transform 1 0 340 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1607101874
transform 1 0 348 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_251
timestamp 1607101874
transform 1 0 356 0 -1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_56
timestamp 1607101874
transform 1 0 380 0 -1 505
box -2 -3 74 103
use MUX2X1  MUX2X1_396
timestamp 1607101874
transform -1 0 500 0 -1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_723
timestamp 1607101874
transform 1 0 500 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_611
timestamp 1607101874
transform -1 0 556 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_523
timestamp 1607101874
transform 1 0 556 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_291
timestamp 1607101874
transform -1 0 676 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_612
timestamp 1607101874
transform 1 0 676 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_325
timestamp 1607101874
transform -1 0 756 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_180
timestamp 1607101874
transform -1 0 780 0 -1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_321
timestamp 1607101874
transform -1 0 828 0 -1 505
box -2 -3 50 103
use FILL  FILL_4_1_0
timestamp 1607101874
transform -1 0 836 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1607101874
transform -1 0 844 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1032
timestamp 1607101874
transform -1 0 940 0 -1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_326
timestamp 1607101874
transform 1 0 940 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_456
timestamp 1607101874
transform -1 0 1004 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_295
timestamp 1607101874
transform -1 0 1100 0 -1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_614
timestamp 1607101874
transform 1 0 1100 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_726
timestamp 1607101874
transform -1 0 1156 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_526
timestamp 1607101874
transform 1 0 1156 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_339
timestamp 1607101874
transform -1 0 1276 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_301
timestamp 1607101874
transform 1 0 1276 0 -1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_328
timestamp 1607101874
transform 1 0 1300 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_458
timestamp 1607101874
transform -1 0 1364 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_2_0
timestamp 1607101874
transform 1 0 1364 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1607101874
transform 1 0 1372 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_297
timestamp 1607101874
transform 1 0 1380 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_286
timestamp 1607101874
transform 1 0 1476 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_845
timestamp 1607101874
transform 1 0 1572 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_768
timestamp 1607101874
transform -1 0 1700 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_766
timestamp 1607101874
transform -1 0 1732 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_427
timestamp 1607101874
transform 1 0 1732 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1607101874
transform -1 0 1852 0 -1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_563
timestamp 1607101874
transform 1 0 1852 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_675
timestamp 1607101874
transform 1 0 1900 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_922
timestamp 1607101874
transform 1 0 1924 0 -1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_37
timestamp 1607101874
transform -1 0 1996 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_923
timestamp 1607101874
transform 1 0 1996 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_245
timestamp 1607101874
transform 1 0 2028 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_585
timestamp 1607101874
transform 1 0 2044 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_267
timestamp 1607101874
transform -1 0 2108 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_586
timestamp 1607101874
transform 1 0 2108 0 -1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_5
timestamp 1607101874
transform 1 0 2140 0 -1 505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1607101874
transform -1 0 2276 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1389
timestamp 1607101874
transform 1 0 2276 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1388
timestamp 1607101874
transform -1 0 2340 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1382
timestamp 1607101874
transform -1 0 2372 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_4_0
timestamp 1607101874
transform 1 0 2372 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1607101874
transform 1 0 2380 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_185
timestamp 1607101874
transform 1 0 2388 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_184
timestamp 1607101874
transform 1 0 2420 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_214
timestamp 1607101874
transform -1 0 2476 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_863
timestamp 1607101874
transform -1 0 2572 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_694
timestamp 1607101874
transform -1 0 2668 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_59
timestamp 1607101874
transform 1 0 2668 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_27
timestamp 1607101874
transform -1 0 2724 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1607101874
transform -1 0 2820 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_73
timestamp 1607101874
transform -1 0 2852 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_74
timestamp 1607101874
transform -1 0 2884 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_5_0
timestamp 1607101874
transform 1 0 2884 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1607101874
transform 1 0 2892 0 -1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_404
timestamp 1607101874
transform 1 0 2900 0 -1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_286
timestamp 1607101874
transform 1 0 2948 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_616
timestamp 1607101874
transform 1 0 2980 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_405
timestamp 1607101874
transform 1 0 3012 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1607101874
transform 1 0 3060 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1272
timestamp 1607101874
transform 1 0 3156 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1271
timestamp 1607101874
transform -1 0 3220 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1607101874
transform -1 0 3252 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1607101874
transform -1 0 3284 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1607101874
transform -1 0 3316 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1268
timestamp 1607101874
transform 1 0 3316 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1267
timestamp 1607101874
transform 1 0 3348 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1607101874
transform -1 0 3412 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_710
timestamp 1607101874
transform 1 0 3428 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_420
timestamp 1607101874
transform -1 0 3548 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_90
timestamp 1607101874
transform 1 0 3548 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1607101874
transform -1 0 3612 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1607101874
transform 1 0 3612 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1275
timestamp 1607101874
transform 1 0 3708 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1276
timestamp 1607101874
transform -1 0 3772 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_417
timestamp 1607101874
transform -1 0 3796 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_328
timestamp 1607101874
transform -1 0 3828 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_419
timestamp 1607101874
transform 1 0 3828 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_418
timestamp 1607101874
transform 1 0 3852 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_741
timestamp 1607101874
transform -1 0 3908 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_7_0
timestamp 1607101874
transform 1 0 3908 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_7_1
timestamp 1607101874
transform 1 0 3916 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_1283
timestamp 1607101874
transform 1 0 3924 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1284
timestamp 1607101874
transform -1 0 3988 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1607101874
transform -1 0 4012 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_32
timestamp 1607101874
transform -1 0 4044 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_703
timestamp 1607101874
transform -1 0 4140 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_334
timestamp 1607101874
transform -1 0 4172 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_326
timestamp 1607101874
transform -1 0 4204 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_740
timestamp 1607101874
transform -1 0 4236 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_383
timestamp 1607101874
transform -1 0 4332 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_633
timestamp 1607101874
transform 1 0 4332 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_521
timestamp 1607101874
transform -1 0 4388 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_449
timestamp 1607101874
transform -1 0 4412 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_866
timestamp 1607101874
transform 1 0 4412 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_8_0
timestamp 1607101874
transform 1 0 4444 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_8_1
timestamp 1607101874
transform 1 0 4452 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_382
timestamp 1607101874
transform 1 0 4460 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_383
timestamp 1607101874
transform -1 0 4524 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1607101874
transform -1 0 4620 0 -1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_5
timestamp 1607101874
transform -1 0 4652 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1235
timestamp 1607101874
transform -1 0 4684 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_193
timestamp 1607101874
transform -1 0 4708 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_343
timestamp 1607101874
transform -1 0 4740 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1233
timestamp 1607101874
transform 1 0 4740 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1607101874
transform -1 0 4868 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_387
timestamp 1607101874
transform 1 0 4868 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_386
timestamp 1607101874
transform -1 0 4932 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_9_0
timestamp 1607101874
transform 1 0 4932 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_9_1
timestamp 1607101874
transform 1 0 4940 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1607101874
transform 1 0 4948 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_12
timestamp 1607101874
transform 1 0 5044 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1607101874
transform 1 0 5076 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_442
timestamp 1607101874
transform -1 0 5132 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_814
timestamp 1607101874
transform 1 0 5132 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_624
timestamp 1607101874
transform -1 0 5260 0 -1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_15
timestamp 1607101874
transform -1 0 5292 0 -1 505
box -2 -3 34 103
use FILL  FILL_5_1
timestamp 1607101874
transform -1 0 5300 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1607101874
transform -1 0 5308 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1029
timestamp 1607101874
transform 1 0 4 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1054
timestamp 1607101874
transform 1 0 100 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_522
timestamp 1607101874
transform 1 0 196 0 1 505
box -2 -3 98 103
use INVX1  INVX1_437
timestamp 1607101874
transform 1 0 292 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_388
timestamp 1607101874
transform -1 0 356 0 1 505
box -2 -3 50 103
use FILL  FILL_5_0_0
timestamp 1607101874
transform 1 0 356 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1607101874
transform 1 0 364 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1051
timestamp 1607101874
transform 1 0 372 0 1 505
box -2 -3 98 103
use INVX1  INVX1_282
timestamp 1607101874
transform 1 0 468 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_655
timestamp 1607101874
transform 1 0 484 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_207
timestamp 1607101874
transform 1 0 516 0 1 505
box -2 -3 26 103
use INVX1  INVX1_388
timestamp 1607101874
transform -1 0 556 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1052
timestamp 1607101874
transform 1 0 556 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_266
timestamp 1607101874
transform 1 0 652 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_524
timestamp 1607101874
transform 1 0 676 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_724
timestamp 1607101874
transform 1 0 772 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_969
timestamp 1607101874
transform 1 0 796 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_592
timestamp 1607101874
transform 1 0 828 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1607101874
transform -1 0 868 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1607101874
transform -1 0 876 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_243
timestamp 1607101874
transform -1 0 900 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_784
timestamp 1607101874
transform 1 0 900 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_236
timestamp 1607101874
transform 1 0 932 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_149
timestamp 1607101874
transform -1 0 988 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_424
timestamp 1607101874
transform -1 0 1020 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_613
timestamp 1607101874
transform 1 0 1020 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_511
timestamp 1607101874
transform -1 0 1148 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_725
timestamp 1607101874
transform -1 0 1172 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_525
timestamp 1607101874
transform -1 0 1268 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1167
timestamp 1607101874
transform 1 0 1268 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1004
timestamp 1607101874
transform 1 0 1300 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_302
timestamp 1607101874
transform 1 0 1332 0 1 505
box -2 -3 26 103
use FILL  FILL_5_2_0
timestamp 1607101874
transform 1 0 1356 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1607101874
transform 1 0 1364 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_1005
timestamp 1607101874
transform 1 0 1372 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_837
timestamp 1607101874
transform 1 0 1404 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1367
timestamp 1607101874
transform 1 0 1500 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1366
timestamp 1607101874
transform -1 0 1564 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_173
timestamp 1607101874
transform 1 0 1564 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1607101874
transform 1 0 1596 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1370
timestamp 1607101874
transform 1 0 1628 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1371
timestamp 1607101874
transform -1 0 1692 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_288
timestamp 1607101874
transform 1 0 1692 0 1 505
box -2 -3 98 103
use INVX1  INVX1_394
timestamp 1607101874
transform 1 0 1788 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_545
timestamp 1607101874
transform 1 0 1804 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1002
timestamp 1607101874
transform 1 0 1828 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1607101874
transform -1 0 1868 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1607101874
transform -1 0 1876 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_398
timestamp 1607101874
transform -1 0 1908 0 1 505
box -2 -3 34 103
use INVX1  INVX1_353
timestamp 1607101874
transform 1 0 1908 0 1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_477
timestamp 1607101874
transform 1 0 1924 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_150
timestamp 1607101874
transform -1 0 1988 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1123
timestamp 1607101874
transform -1 0 2020 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1125
timestamp 1607101874
transform -1 0 2052 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_584
timestamp 1607101874
transform -1 0 2084 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_476
timestamp 1607101874
transform 1 0 2084 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1372
timestamp 1607101874
transform 1 0 2116 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1373
timestamp 1607101874
transform -1 0 2180 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_289
timestamp 1607101874
transform -1 0 2276 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_169
timestamp 1607101874
transform 1 0 2276 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_843
timestamp 1607101874
transform 1 0 2308 0 1 505
box -2 -3 98 103
use FILL  FILL_5_4_0
timestamp 1607101874
transform -1 0 2412 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1607101874
transform -1 0 2420 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_168
timestamp 1607101874
transform -1 0 2452 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_571
timestamp 1607101874
transform -1 0 2476 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1182
timestamp 1607101874
transform -1 0 2508 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_690
timestamp 1607101874
transform -1 0 2604 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_56
timestamp 1607101874
transform 1 0 2604 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1607101874
transform -1 0 2660 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_697
timestamp 1607101874
transform -1 0 2756 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_30
timestamp 1607101874
transform 1 0 2756 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_63
timestamp 1607101874
transform 1 0 2788 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_270
timestamp 1607101874
transform -1 0 2860 0 1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_359
timestamp 1607101874
transform -1 0 2892 0 1 505
box -2 -3 34 103
use FILL  FILL_5_5_0
timestamp 1607101874
transform -1 0 2900 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1607101874
transform -1 0 2908 0 1 505
box -2 -3 10 103
use INVX1  INVX1_362
timestamp 1607101874
transform -1 0 2924 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1607101874
transform -1 0 3020 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_247
timestamp 1607101874
transform 1 0 3020 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_822
timestamp 1607101874
transform -1 0 3076 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_583
timestamp 1607101874
transform -1 0 3172 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1087
timestamp 1607101874
transform 1 0 3172 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_465
timestamp 1607101874
transform -1 0 3236 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_35
timestamp 1607101874
transform 1 0 3236 0 1 505
box -2 -3 74 103
use BUFX4  BUFX4_301
timestamp 1607101874
transform 1 0 3308 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1607101874
transform 1 0 3340 0 1 505
box -2 -3 98 103
use FILL  FILL_5_6_0
timestamp 1607101874
transform 1 0 3436 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1607101874
transform 1 0 3444 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_524
timestamp 1607101874
transform 1 0 3452 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_636
timestamp 1607101874
transform 1 0 3484 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_523
timestamp 1607101874
transform 1 0 3508 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1184
timestamp 1607101874
transform 1 0 3532 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1090
timestamp 1607101874
transform -1 0 3596 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_299
timestamp 1607101874
transform 1 0 3596 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_249
timestamp 1607101874
transform -1 0 3660 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_43
timestamp 1607101874
transform 1 0 3660 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1138
timestamp 1607101874
transform -1 0 3724 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_614
timestamp 1607101874
transform -1 0 3820 0 1 505
box -2 -3 98 103
use INVX1  INVX1_21
timestamp 1607101874
transform 1 0 3820 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_16
timestamp 1607101874
transform -1 0 3884 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_703
timestamp 1607101874
transform -1 0 3916 0 1 505
box -2 -3 34 103
use FILL  FILL_5_7_0
timestamp 1607101874
transform 1 0 3916 0 1 505
box -2 -3 10 103
use FILL  FILL_5_7_1
timestamp 1607101874
transform 1 0 3924 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_404
timestamp 1607101874
transform 1 0 3932 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_701
timestamp 1607101874
transform -1 0 3988 0 1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_17
timestamp 1607101874
transform -1 0 4028 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_403
timestamp 1607101874
transform -1 0 4052 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1607101874
transform -1 0 4148 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_635
timestamp 1607101874
transform 1 0 4148 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_523
timestamp 1607101874
transform -1 0 4204 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_385
timestamp 1607101874
transform -1 0 4300 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1607101874
transform -1 0 4396 0 1 505
box -2 -3 98 103
use FILL  FILL_5_8_0
timestamp 1607101874
transform -1 0 4404 0 1 505
box -2 -3 10 103
use FILL  FILL_5_8_1
timestamp 1607101874
transform -1 0 4412 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1607101874
transform -1 0 4508 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_180
timestamp 1607101874
transform 1 0 4508 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_277
timestamp 1607101874
transform 1 0 4540 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_421
timestamp 1607101874
transform -1 0 4596 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1607101874
transform -1 0 4620 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_635
timestamp 1607101874
transform -1 0 4716 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_159
timestamp 1607101874
transform 1 0 4716 0 1 505
box -2 -3 34 103
use INVX1  INVX1_170
timestamp 1607101874
transform -1 0 4764 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1607101874
transform -1 0 4860 0 1 505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_91
timestamp 1607101874
transform -1 0 4932 0 1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_605
timestamp 1607101874
transform -1 0 4956 0 1 505
box -2 -3 26 103
use FILL  FILL_5_9_0
timestamp 1607101874
transform 1 0 4956 0 1 505
box -2 -3 10 103
use FILL  FILL_5_9_1
timestamp 1607101874
transform 1 0 4964 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_375
timestamp 1607101874
transform 1 0 4972 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_290
timestamp 1607101874
transform -1 0 5036 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_505
timestamp 1607101874
transform -1 0 5068 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_93
timestamp 1607101874
transform 1 0 5068 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_816
timestamp 1607101874
transform 1 0 5092 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_356
timestamp 1607101874
transform -1 0 5156 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1607101874
transform 1 0 5156 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_5
timestamp 1607101874
transform -1 0 5212 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_599
timestamp 1607101874
transform -1 0 5308 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_130
timestamp 1607101874
transform -1 0 52 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_143
timestamp 1607101874
transform -1 0 68 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_335
timestamp 1607101874
transform 1 0 68 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_334
timestamp 1607101874
transform -1 0 132 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_444
timestamp 1607101874
transform 1 0 132 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_1258
timestamp 1607101874
transform 1 0 148 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_387
timestamp 1607101874
transform 1 0 180 0 -1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_458
timestamp 1607101874
transform 1 0 196 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_329
timestamp 1607101874
transform 1 0 228 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_328
timestamp 1607101874
transform 1 0 260 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_330
timestamp 1607101874
transform 1 0 292 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1607101874
transform -1 0 332 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1607101874
transform -1 0 340 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_331
timestamp 1607101874
transform -1 0 372 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_292
timestamp 1607101874
transform -1 0 396 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_547
timestamp 1607101874
transform 1 0 396 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_970
timestamp 1607101874
transform -1 0 524 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1033
timestamp 1607101874
transform 1 0 524 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_150
timestamp 1607101874
transform 1 0 620 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_237
timestamp 1607101874
transform -1 0 676 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_340
timestamp 1607101874
transform 1 0 676 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_886
timestamp 1607101874
transform 1 0 692 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_330
timestamp 1607101874
transform 1 0 724 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_303
timestamp 1607101874
transform 1 0 748 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_1_0
timestamp 1607101874
transform -1 0 852 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1607101874
transform -1 0 860 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_234
timestamp 1607101874
transform -1 0 884 0 -1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_62
timestamp 1607101874
transform 1 0 884 0 -1 705
box -2 -3 74 103
use NAND2X1  NAND2X1_188
timestamp 1607101874
transform -1 0 980 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_378
timestamp 1607101874
transform -1 0 1012 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_381
timestamp 1607101874
transform -1 0 1060 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_266
timestamp 1607101874
transform -1 0 1076 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1022
timestamp 1607101874
transform -1 0 1172 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_287
timestamp 1607101874
transform -1 0 1196 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_92
timestamp 1607101874
transform -1 0 1244 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_867
timestamp 1607101874
transform 1 0 1244 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_105
timestamp 1607101874
transform 1 0 1340 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_2_0
timestamp 1607101874
transform 1 0 1356 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1607101874
transform 1 0 1364 0 -1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_82
timestamp 1607101874
transform 1 0 1372 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_95
timestamp 1607101874
transform -1 0 1436 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_1009
timestamp 1607101874
transform 1 0 1436 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_306
timestamp 1607101874
transform -1 0 1492 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_145
timestamp 1607101874
transform -1 0 1516 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_272
timestamp 1607101874
transform 1 0 1516 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1379
timestamp 1607101874
transform -1 0 1644 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1378
timestamp 1607101874
transform -1 0 1676 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_351
timestamp 1607101874
transform 1 0 1676 0 -1 705
box -2 -3 18 103
use BUFX4  BUFX4_130
timestamp 1607101874
transform -1 0 1724 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_127
timestamp 1607101874
transform 1 0 1724 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_423
timestamp 1607101874
transform 1 0 1756 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_921
timestamp 1607101874
transform 1 0 1772 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1001
timestamp 1607101874
transform -1 0 1836 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_393
timestamp 1607101874
transform -1 0 1852 0 -1 705
box -2 -3 18 103
use BUFX4  BUFX4_129
timestamp 1607101874
transform 1 0 1852 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_180
timestamp 1607101874
transform 1 0 1900 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_181
timestamp 1607101874
transform -1 0 1964 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_853
timestamp 1607101874
transform -1 0 2060 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1126
timestamp 1607101874
transform -1 0 2092 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_243
timestamp 1607101874
transform -1 0 2108 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_270
timestamp 1607101874
transform -1 0 2204 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1374
timestamp 1607101874
transform -1 0 2236 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1375
timestamp 1607101874
transform -1 0 2268 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_685
timestamp 1607101874
transform -1 0 2300 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1607101874
transform -1 0 2396 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_4_0
timestamp 1607101874
transform -1 0 2404 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1607101874
transform -1 0 2412 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1181
timestamp 1607101874
transform -1 0 2444 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_67
timestamp 1607101874
transform -1 0 2484 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_572
timestamp 1607101874
transform -1 0 2508 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_698
timestamp 1607101874
transform -1 0 2604 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_64
timestamp 1607101874
transform 1 0 2604 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1607101874
transform -1 0 2660 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_57
timestamp 1607101874
transform -1 0 2684 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1556
timestamp 1607101874
transform 1 0 2684 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_584
timestamp 1607101874
transform 1 0 2716 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_796
timestamp 1607101874
transform 1 0 2812 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1555
timestamp 1607101874
transform -1 0 2876 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_349
timestamp 1607101874
transform -1 0 2908 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_5_0
timestamp 1607101874
transform 1 0 2908 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1607101874
transform 1 0 2916 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1554
timestamp 1607101874
transform 1 0 2924 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1553
timestamp 1607101874
transform 1 0 2956 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1607101874
transform 1 0 2988 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1287
timestamp 1607101874
transform -1 0 3116 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1288
timestamp 1607101874
transform -1 0 3148 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_628
timestamp 1607101874
transform 1 0 3148 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_516
timestamp 1607101874
transform -1 0 3204 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1607101874
transform -1 0 3300 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_60
timestamp 1607101874
transform -1 0 3324 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_42
timestamp 1607101874
transform -1 0 3356 0 -1 705
box -2 -3 34 103
use INVX8  INVX8_12
timestamp 1607101874
transform -1 0 3396 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_6_0
timestamp 1607101874
transform 1 0 3396 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1607101874
transform 1 0 3404 0 -1 705
box -2 -3 10 103
use OAI22X1  OAI22X1_49
timestamp 1607101874
transform 1 0 3412 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_522
timestamp 1607101874
transform 1 0 3452 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_157
timestamp 1607101874
transform -1 0 3508 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1607101874
transform 1 0 3508 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1607101874
transform -1 0 3564 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1607101874
transform -1 0 3660 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1279
timestamp 1607101874
transform -1 0 3692 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1280
timestamp 1607101874
transform -1 0 3724 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_602
timestamp 1607101874
transform 1 0 3724 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_8
timestamp 1607101874
transform 1 0 3820 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1607101874
transform -1 0 3876 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_7_0
timestamp 1607101874
transform -1 0 3884 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_7_1
timestamp 1607101874
transform -1 0 3892 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1607101874
transform -1 0 3988 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1282
timestamp 1607101874
transform 1 0 3988 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1281
timestamp 1607101874
transform 1 0 4020 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_557
timestamp 1607101874
transform 1 0 4052 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1607101874
transform -1 0 4108 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_251
timestamp 1607101874
transform -1 0 4140 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_393
timestamp 1607101874
transform 1 0 4140 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_394
timestamp 1607101874
transform -1 0 4204 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1607101874
transform -1 0 4228 0 -1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_76
timestamp 1607101874
transform -1 0 4300 0 -1 705
box -2 -3 74 103
use NOR2X1  NOR2X1_505
timestamp 1607101874
transform -1 0 4324 0 -1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_28
timestamp 1607101874
transform -1 0 4396 0 -1 705
box -2 -3 74 103
use OAI21X1  OAI21X1_404
timestamp 1607101874
transform 1 0 4396 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_8_0
timestamp 1607101874
transform -1 0 4436 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_8_1
timestamp 1607101874
transform -1 0 4444 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1607101874
transform -1 0 4540 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_287
timestamp 1607101874
transform 1 0 4540 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_190
timestamp 1607101874
transform -1 0 4596 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1041
timestamp 1607101874
transform -1 0 4628 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_45
timestamp 1607101874
transform 1 0 4628 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_628
timestamp 1607101874
transform 1 0 4668 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_157
timestamp 1607101874
transform 1 0 4700 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_603
timestamp 1607101874
transform 1 0 4748 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_8
timestamp 1607101874
transform 1 0 4844 0 -1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_5
timestamp 1607101874
transform -1 0 4908 0 -1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_622
timestamp 1607101874
transform 1 0 4908 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_9_0
timestamp 1607101874
transform 1 0 4940 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_9_1
timestamp 1607101874
transform 1 0 4948 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1142
timestamp 1607101874
transform 1 0 4956 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_274
timestamp 1607101874
transform -1 0 5004 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_401
timestamp 1607101874
transform 1 0 5004 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_402
timestamp 1607101874
transform -1 0 5068 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1607101874
transform -1 0 5164 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_29
timestamp 1607101874
transform 1 0 5164 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_648
timestamp 1607101874
transform -1 0 5292 0 -1 705
box -2 -3 98 103
use FILL  FILL_7_1
timestamp 1607101874
transform -1 0 5300 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1607101874
transform -1 0 5308 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_6
timestamp 1607101874
transform -1 0 36 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_97
timestamp 1607101874
transform 1 0 36 0 1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_545
timestamp 1607101874
transform 1 0 108 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1534
timestamp 1607101874
transform -1 0 236 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_519
timestamp 1607101874
transform 1 0 236 0 1 705
box -2 -3 98 103
use FILL  FILL_7_0_0
timestamp 1607101874
transform 1 0 332 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1607101874
transform 1 0 340 0 1 705
box -2 -3 10 103
use INVX1  INVX1_267
timestamp 1607101874
transform 1 0 348 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_385
timestamp 1607101874
transform 1 0 364 0 1 705
box -2 -3 50 103
use AOI21X1  AOI21X1_618
timestamp 1607101874
transform 1 0 412 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_730
timestamp 1607101874
transform -1 0 468 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_250
timestamp 1607101874
transform 1 0 468 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_222
timestamp 1607101874
transform 1 0 492 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_731
timestamp 1607101874
transform 1 0 516 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_306
timestamp 1607101874
transform -1 0 708 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_233
timestamp 1607101874
transform -1 0 732 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1072
timestamp 1607101874
transform -1 0 764 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_555
timestamp 1607101874
transform 1 0 764 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_667
timestamp 1607101874
transform -1 0 820 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_238
timestamp 1607101874
transform 1 0 820 0 1 705
box -2 -3 50 103
use FILL  FILL_7_1_0
timestamp 1607101874
transform 1 0 868 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1607101874
transform 1 0 876 0 1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_2
timestamp 1607101874
transform 1 0 884 0 1 705
box -2 -3 74 103
use OAI21X1  OAI21X1_612
timestamp 1607101874
transform -1 0 988 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_762
timestamp 1607101874
transform 1 0 988 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_236
timestamp 1607101874
transform -1 0 1044 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_515
timestamp 1607101874
transform 1 0 1044 0 1 705
box -2 -3 98 103
use INVX1  INVX1_140
timestamp 1607101874
transform 1 0 1140 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_127
timestamp 1607101874
transform -1 0 1204 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_964
timestamp 1607101874
transform -1 0 1236 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_142
timestamp 1607101874
transform -1 0 1260 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1255
timestamp 1607101874
transform 1 0 1260 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_140
timestamp 1607101874
transform -1 0 1316 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_379
timestamp 1607101874
transform -1 0 1348 0 1 705
box -2 -3 34 103
use FILL  FILL_7_2_0
timestamp 1607101874
transform -1 0 1356 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1607101874
transform -1 0 1364 0 1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_265
timestamp 1607101874
transform -1 0 1412 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_86
timestamp 1607101874
transform 1 0 1412 0 1 705
box -2 -3 50 103
use INVX1  INVX1_99
timestamp 1607101874
transform -1 0 1476 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_841
timestamp 1607101874
transform -1 0 1572 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_241
timestamp 1607101874
transform -1 0 1620 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_273
timestamp 1607101874
transform 1 0 1620 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1380
timestamp 1607101874
transform 1 0 1716 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1381
timestamp 1607101874
transform -1 0 1780 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_433
timestamp 1607101874
transform 1 0 1780 0 1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_58
timestamp 1607101874
transform 1 0 1812 0 1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_544
timestamp 1607101874
transform 1 0 1852 0 1 705
box -2 -3 26 103
use FILL  FILL_7_3_0
timestamp 1607101874
transform -1 0 1884 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1607101874
transform -1 0 1892 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1607101874
transform -1 0 1988 0 1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_564
timestamp 1607101874
transform 1 0 1988 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_676
timestamp 1607101874
transform 1 0 2020 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_131
timestamp 1607101874
transform 1 0 2044 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_78
timestamp 1607101874
transform 1 0 2076 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_134
timestamp 1607101874
transform -1 0 2132 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_850
timestamp 1607101874
transform 1 0 2132 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_396
timestamp 1607101874
transform -1 0 2252 0 1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_14
timestamp 1607101874
transform -1 0 2292 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_686
timestamp 1607101874
transform 1 0 2292 0 1 705
box -2 -3 34 103
use INVX1  INVX1_150
timestamp 1607101874
transform 1 0 2324 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_764
timestamp 1607101874
transform -1 0 2372 0 1 705
box -2 -3 34 103
use FILL  FILL_7_4_0
timestamp 1607101874
transform -1 0 2380 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1607101874
transform -1 0 2388 0 1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_137
timestamp 1607101874
transform -1 0 2436 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_1020
timestamp 1607101874
transform 1 0 2436 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_309
timestamp 1607101874
transform -1 0 2492 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_559
timestamp 1607101874
transform 1 0 2492 0 1 705
box -2 -3 98 103
use INVX1  INVX1_268
timestamp 1607101874
transform 1 0 2588 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_405
timestamp 1607101874
transform -1 0 2636 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_934
timestamp 1607101874
transform -1 0 2668 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1607101874
transform -1 0 2764 0 1 705
box -2 -3 98 103
use INVX1  INVX1_153
timestamp 1607101874
transform 1 0 2764 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_140
timestamp 1607101874
transform -1 0 2828 0 1 705
box -2 -3 50 103
use AOI21X1  AOI21X1_406
timestamp 1607101874
transform -1 0 2860 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_935
timestamp 1607101874
transform -1 0 2892 0 1 705
box -2 -3 34 103
use FILL  FILL_7_5_0
timestamp 1607101874
transform -1 0 2900 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1607101874
transform -1 0 2908 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_76
timestamp 1607101874
transform -1 0 2940 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_256
timestamp 1607101874
transform -1 0 2988 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_1089
timestamp 1607101874
transform -1 0 3020 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1088
timestamp 1607101874
transform -1 0 3052 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1091
timestamp 1607101874
transform 1 0 3052 0 1 705
box -2 -3 34 103
use INVX1  INVX1_46
timestamp 1607101874
transform -1 0 3100 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_713
timestamp 1607101874
transform -1 0 3196 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_38
timestamp 1607101874
transform -1 0 3244 0 1 705
box -2 -3 50 103
use CLKBUF1  CLKBUF1_19
timestamp 1607101874
transform 1 0 3244 0 1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1607101874
transform -1 0 3412 0 1 705
box -2 -3 98 103
use FILL  FILL_7_6_0
timestamp 1607101874
transform 1 0 3412 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1607101874
transform 1 0 3420 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1270
timestamp 1607101874
transform 1 0 3428 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1269
timestamp 1607101874
transform -1 0 3492 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_54
timestamp 1607101874
transform -1 0 3516 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_68
timestamp 1607101874
transform 1 0 3516 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1607101874
transform -1 0 3572 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_705
timestamp 1607101874
transform -1 0 3668 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_79
timestamp 1607101874
transform 1 0 3668 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_701
timestamp 1607101874
transform -1 0 3796 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_80
timestamp 1607101874
transform -1 0 3828 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_707
timestamp 1607101874
transform 1 0 3828 0 1 705
box -2 -3 98 103
use FILL  FILL_7_7_0
timestamp 1607101874
transform 1 0 3924 0 1 705
box -2 -3 10 103
use FILL  FILL_7_7_1
timestamp 1607101874
transform 1 0 3932 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_83
timestamp 1607101874
transform 1 0 3940 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_84
timestamp 1607101874
transform -1 0 4004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_702
timestamp 1607101874
transform 1 0 4004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1277
timestamp 1607101874
transform -1 0 4068 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1278
timestamp 1607101874
transform -1 0 4100 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_8
timestamp 1607101874
transform 1 0 4100 0 1 705
box -2 -3 50 103
use INVX1  INVX1_11
timestamp 1607101874
transform -1 0 4164 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_558
timestamp 1607101874
transform -1 0 4196 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1607101874
transform -1 0 4292 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_606
timestamp 1607101874
transform -1 0 4388 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_555
timestamp 1607101874
transform -1 0 4412 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_403
timestamp 1607101874
transform -1 0 4444 0 1 705
box -2 -3 34 103
use FILL  FILL_7_8_0
timestamp 1607101874
transform 1 0 4444 0 1 705
box -2 -3 10 103
use FILL  FILL_7_8_1
timestamp 1607101874
transform 1 0 4452 0 1 705
box -2 -3 10 103
use BUFX4  BUFX4_7
timestamp 1607101874
transform 1 0 4460 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1607101874
transform -1 0 4588 0 1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_40
timestamp 1607101874
transform -1 0 4660 0 1 705
box -2 -3 74 103
use INVX1  INVX1_166
timestamp 1607101874
transform -1 0 4676 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1607101874
transform -1 0 4772 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_604
timestamp 1607101874
transform -1 0 4796 0 1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_83
timestamp 1607101874
transform -1 0 4836 0 1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_626
timestamp 1607101874
transform 1 0 4836 0 1 705
box -2 -3 98 103
use FILL  FILL_7_9_0
timestamp 1607101874
transform -1 0 4940 0 1 705
box -2 -3 10 103
use FILL  FILL_7_9_1
timestamp 1607101874
transform -1 0 4948 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1143
timestamp 1607101874
transform -1 0 4980 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_558
timestamp 1607101874
transform -1 0 5004 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_17
timestamp 1607101874
transform 1 0 5004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_16
timestamp 1607101874
transform -1 0 5068 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_295
timestamp 1607101874
transform 1 0 5068 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1607101874
transform 1 0 5100 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1607101874
transform -1 0 5164 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_647
timestamp 1607101874
transform -1 0 5260 0 1 705
box -2 -3 98 103
use INVX1  INVX1_180
timestamp 1607101874
transform -1 0 5276 0 1 705
box -2 -3 18 103
use INVX1  INVX1_167
timestamp 1607101874
transform -1 0 5292 0 1 705
box -2 -3 18 103
use FILL  FILL_8_1
timestamp 1607101874
transform 1 0 5292 0 1 705
box -2 -3 10 103
use FILL  FILL_8_2
timestamp 1607101874
transform 1 0 5300 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_550
timestamp 1607101874
transform 1 0 4 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_621
timestamp 1607101874
transform 1 0 100 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_733
timestamp 1607101874
transform -1 0 156 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1533
timestamp 1607101874
transform 1 0 156 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1077
timestamp 1607101874
transform 1 0 188 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1076
timestamp 1607101874
transform -1 0 252 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_557
timestamp 1607101874
transform 1 0 252 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_0_0
timestamp 1607101874
transform -1 0 356 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1607101874
transform -1 0 364 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1607101874
transform -1 0 460 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_135
timestamp 1607101874
transform 1 0 460 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_46
timestamp 1607101874
transform -1 0 556 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_704
timestamp 1607101874
transform -1 0 588 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1607101874
transform -1 0 604 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1358
timestamp 1607101874
transform 1 0 604 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1359
timestamp 1607101874
transform -1 0 668 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_556
timestamp 1607101874
transform 1 0 668 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_668
timestamp 1607101874
transform -1 0 724 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_307
timestamp 1607101874
transform 1 0 724 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1361
timestamp 1607101874
transform 1 0 820 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_1_0
timestamp 1607101874
transform -1 0 860 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1607101874
transform -1 0 868 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_1360
timestamp 1607101874
transform -1 0 900 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_125
timestamp 1607101874
transform -1 0 924 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_235
timestamp 1607101874
transform -1 0 948 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1024
timestamp 1607101874
transform 1 0 948 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1506
timestamp 1607101874
transform 1 0 1044 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1505
timestamp 1607101874
transform -1 0 1108 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1026
timestamp 1607101874
transform 1 0 1108 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_310
timestamp 1607101874
transform 1 0 1204 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_311
timestamp 1607101874
transform -1 0 1268 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_348
timestamp 1607101874
transform 1 0 1268 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_842
timestamp 1607101874
transform 1 0 1292 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_2_0
timestamp 1607101874
transform 1 0 1388 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1607101874
transform 1 0 1396 0 -1 905
box -2 -3 10 103
use INVX1  INVX1_100
timestamp 1607101874
transform 1 0 1404 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_87
timestamp 1607101874
transform -1 0 1468 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_684
timestamp 1607101874
transform 1 0 1468 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_136
timestamp 1607101874
transform 1 0 1500 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1607101874
transform 1 0 1532 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_677
timestamp 1607101874
transform -1 0 1652 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_565
timestamp 1607101874
transform -1 0 1684 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1124
timestamp 1607101874
transform 1 0 1684 0 -1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_44
timestamp 1607101874
transform -1 0 1756 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_1003
timestamp 1607101874
transform -1 0 1788 0 -1 905
box -2 -3 34 103
use AND2X2  AND2X2_44
timestamp 1607101874
transform -1 0 1820 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_849
timestamp 1607101874
transform -1 0 1916 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_3_0
timestamp 1607101874
transform 1 0 1916 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1607101874
transform 1 0 1924 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_133
timestamp 1607101874
transform 1 0 1932 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_77
timestamp 1607101874
transform -1 0 1988 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_846
timestamp 1607101874
transform -1 0 2084 0 -1 905
box -2 -3 98 103
use BUFX4  BUFX4_133
timestamp 1607101874
transform 1 0 2084 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_361
timestamp 1607101874
transform 1 0 2116 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1216
timestamp 1607101874
transform 1 0 2148 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_177
timestamp 1607101874
transform 1 0 2180 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1607101874
transform 1 0 2212 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_851
timestamp 1607101874
transform 1 0 2244 0 -1 905
box -2 -3 98 103
use BUFX4  BUFX4_154
timestamp 1607101874
transform -1 0 2372 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_4_0
timestamp 1607101874
transform -1 0 2380 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1607101874
transform -1 0 2388 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_683
timestamp 1607101874
transform -1 0 2420 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_571
timestamp 1607101874
transform 1 0 2420 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_438
timestamp 1607101874
transform -1 0 2548 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_398
timestamp 1607101874
transform -1 0 2596 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_613
timestamp 1607101874
transform 1 0 2596 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_284
timestamp 1607101874
transform -1 0 2660 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1607101874
transform -1 0 2756 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_322
timestamp 1607101874
transform -1 0 2780 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_263
timestamp 1607101874
transform 1 0 2780 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_168
timestamp 1607101874
transform -1 0 2836 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_1
timestamp 1607101874
transform -1 0 2868 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_5_0
timestamp 1607101874
transform 1 0 2868 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1607101874
transform 1 0 2876 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_708
timestamp 1607101874
transform 1 0 2884 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_824
timestamp 1607101874
transform -1 0 3012 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_85
timestamp 1607101874
transform -1 0 3044 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1607101874
transform -1 0 3076 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_270
timestamp 1607101874
transform -1 0 3100 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_141
timestamp 1607101874
transform 1 0 3100 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1607101874
transform 1 0 3148 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_154
timestamp 1607101874
transform 1 0 3244 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1607101874
transform 1 0 3260 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_177
timestamp 1607101874
transform 1 0 3356 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_274
timestamp 1607101874
transform -1 0 3412 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_501
timestamp 1607101874
transform 1 0 3428 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1224
timestamp 1607101874
transform 1 0 3460 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_500
timestamp 1607101874
transform 1 0 3492 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1021
timestamp 1607101874
transform -1 0 3548 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_562
timestamp 1607101874
transform -1 0 3644 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_559
timestamp 1607101874
transform 1 0 3644 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_124
timestamp 1607101874
transform 1 0 3676 0 -1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_62
timestamp 1607101874
transform -1 0 3748 0 -1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_556
timestamp 1607101874
transform 1 0 3748 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_933
timestamp 1607101874
transform -1 0 3804 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_475
timestamp 1607101874
transform -1 0 3828 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_474
timestamp 1607101874
transform 1 0 3828 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1285
timestamp 1607101874
transform -1 0 3884 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1286
timestamp 1607101874
transform -1 0 3916 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_7_0
timestamp 1607101874
transform -1 0 3924 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_7_1
timestamp 1607101874
transform -1 0 3932 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_1139
timestamp 1607101874
transform -1 0 3964 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_448
timestamp 1607101874
transform 1 0 3964 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_618
timestamp 1607101874
transform -1 0 4092 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_26
timestamp 1607101874
transform 1 0 4092 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_20
timestamp 1607101874
transform -1 0 4156 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_384
timestamp 1607101874
transform 1 0 4156 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_385
timestamp 1607101874
transform -1 0 4220 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_188
timestamp 1607101874
transform 1 0 4220 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_1236
timestamp 1607101874
transform -1 0 4300 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_280
timestamp 1607101874
transform 1 0 4300 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_183
timestamp 1607101874
transform -1 0 4356 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_263
timestamp 1607101874
transform -1 0 4404 0 -1 905
box -2 -3 50 103
use BUFX4  BUFX4_294
timestamp 1607101874
transform -1 0 4436 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_8_0
timestamp 1607101874
transform 1 0 4436 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_8_1
timestamp 1607101874
transform 1 0 4444 0 -1 905
box -2 -3 10 103
use OAI22X1  OAI22X1_84
timestamp 1607101874
transform 1 0 4452 0 -1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_192
timestamp 1607101874
transform 1 0 4492 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_289
timestamp 1607101874
transform -1 0 4548 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_607
timestamp 1607101874
transform 1 0 4548 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_332
timestamp 1607101874
transform -1 0 4604 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_153
timestamp 1607101874
transform 1 0 4604 0 -1 905
box -2 -3 50 103
use BUFX4  BUFX4_293
timestamp 1607101874
transform 1 0 4652 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1607101874
transform 1 0 4684 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_19
timestamp 1607101874
transform -1 0 4740 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_638
timestamp 1607101874
transform 1 0 4740 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1607101874
transform -1 0 4932 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_178
timestamp 1607101874
transform 1 0 4932 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_9_0
timestamp 1607101874
transform -1 0 4956 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_9_1
timestamp 1607101874
transform -1 0 4964 0 -1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_165
timestamp 1607101874
transform -1 0 5012 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_1230
timestamp 1607101874
transform 1 0 5012 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1607101874
transform 1 0 5044 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1607101874
transform 1 0 5076 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1607101874
transform 1 0 5100 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_35
timestamp 1607101874
transform -1 0 5156 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_149
timestamp 1607101874
transform 1 0 5156 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1607101874
transform -1 0 5300 0 -1 905
box -2 -3 98 103
use FILL  FILL_9_1
timestamp 1607101874
transform -1 0 5308 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1053
timestamp 1607101874
transform 1 0 4 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_333
timestamp 1607101874
transform 1 0 100 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1607101874
transform -1 0 164 0 1 905
box -2 -3 34 103
use INVX1  INVX1_406
timestamp 1607101874
transform 1 0 164 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_656
timestamp 1607101874
transform -1 0 212 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1078
timestamp 1607101874
transform 1 0 212 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_49
timestamp 1607101874
transform -1 0 276 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1542
timestamp 1607101874
transform 1 0 276 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_351
timestamp 1607101874
transform 1 0 308 0 1 905
box -2 -3 26 103
use FILL  FILL_9_0_0
timestamp 1607101874
transform 1 0 332 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1607101874
transform 1 0 340 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_322
timestamp 1607101874
transform 1 0 348 0 1 905
box -2 -3 34 103
use INVX1  INVX1_148
timestamp 1607101874
transform 1 0 380 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1259
timestamp 1607101874
transform -1 0 428 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_198
timestamp 1607101874
transform -1 0 476 0 1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_314
timestamp 1607101874
transform 1 0 476 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_530
timestamp 1607101874
transform 1 0 572 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_642
timestamp 1607101874
transform -1 0 628 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_453
timestamp 1607101874
transform -1 0 660 0 1 905
box -2 -3 34 103
use INVX1  INVX1_250
timestamp 1607101874
transform 1 0 660 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_591
timestamp 1607101874
transform 1 0 676 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_304
timestamp 1607101874
transform 1 0 708 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_893
timestamp 1607101874
transform 1 0 804 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_269
timestamp 1607101874
transform -1 0 860 0 1 905
box -2 -3 26 103
use FILL  FILL_9_1_0
timestamp 1607101874
transform -1 0 868 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1607101874
transform -1 0 876 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_266
timestamp 1607101874
transform -1 0 924 0 1 905
box -2 -3 50 103
use INVX1  INVX1_312
timestamp 1607101874
transform 1 0 924 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_761
timestamp 1607101874
transform -1 0 972 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_210
timestamp 1607101874
transform 1 0 972 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_268
timestamp 1607101874
transform -1 0 1044 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_307
timestamp 1607101874
transform 1 0 1044 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_306
timestamp 1607101874
transform -1 0 1108 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_611
timestamp 1607101874
transform 1 0 1108 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1607101874
transform -1 0 1164 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_185
timestamp 1607101874
transform 1 0 1164 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_1511
timestamp 1607101874
transform 1 0 1212 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1512
timestamp 1607101874
transform -1 0 1276 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_518
timestamp 1607101874
transform -1 0 1372 0 1 905
box -2 -3 98 103
use FILL  FILL_9_2_0
timestamp 1607101874
transform -1 0 1380 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1607101874
transform -1 0 1388 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_467
timestamp 1607101874
transform -1 0 1420 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_86
timestamp 1607101874
transform 1 0 1420 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_146
timestamp 1607101874
transform -1 0 1476 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_215
timestamp 1607101874
transform 1 0 1476 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_871
timestamp 1607101874
transform -1 0 1596 0 1 905
box -2 -3 98 103
use BUFX4  BUFX4_297
timestamp 1607101874
transform 1 0 1596 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_179
timestamp 1607101874
transform -1 0 1676 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_623
timestamp 1607101874
transform -1 0 1700 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_138
timestamp 1607101874
transform -1 0 1724 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_81
timestamp 1607101874
transform -1 0 1756 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_857
timestamp 1607101874
transform -1 0 1852 0 1 905
box -2 -3 98 103
use FILL  FILL_9_3_0
timestamp 1607101874
transform 1 0 1852 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1607101874
transform 1 0 1860 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_858
timestamp 1607101874
transform 1 0 1868 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_82
timestamp 1607101874
transform 1 0 1964 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_139
timestamp 1607101874
transform 1 0 1996 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_174
timestamp 1607101874
transform -1 0 2052 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_175
timestamp 1607101874
transform -1 0 2084 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_88
timestamp 1607101874
transform 1 0 2084 0 1 905
box -2 -3 50 103
use INVX1  INVX1_101
timestamp 1607101874
transform -1 0 2148 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_848
timestamp 1607101874
transform -1 0 2244 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_135
timestamp 1607101874
transform 1 0 2244 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_131
timestamp 1607101874
transform 1 0 2268 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_200
timestamp 1607101874
transform -1 0 2340 0 1 905
box -2 -3 50 103
use CLKBUF1  CLKBUF1_53
timestamp 1607101874
transform -1 0 2412 0 1 905
box -2 -3 74 103
use FILL  FILL_9_4_0
timestamp 1607101874
transform 1 0 2412 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1607101874
transform 1 0 2420 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_624
timestamp 1607101874
transform 1 0 2428 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_736
timestamp 1607101874
transform -1 0 2484 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_563
timestamp 1607101874
transform 1 0 2484 0 1 905
box -2 -3 98 103
use INVX1  INVX1_269
timestamp 1607101874
transform 1 0 2580 0 1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_401
timestamp 1607101874
transform -1 0 2644 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_614
timestamp 1607101874
transform 1 0 2644 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_285
timestamp 1607101874
transform -1 0 2708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_615
timestamp 1607101874
transform 1 0 2708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1056
timestamp 1607101874
transform 1 0 2740 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1607101874
transform 1 0 2772 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1058
timestamp 1607101874
transform 1 0 2796 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_324
timestamp 1607101874
transform -1 0 2852 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_273
timestamp 1607101874
transform 1 0 2852 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_176
timestamp 1607101874
transform -1 0 2908 0 1 905
box -2 -3 34 103
use FILL  FILL_9_5_0
timestamp 1607101874
transform -1 0 2916 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1607101874
transform -1 0 2924 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1607101874
transform -1 0 3020 0 1 905
box -2 -3 98 103
use INVX1  INVX1_329
timestamp 1607101874
transform -1 0 3036 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_580
timestamp 1607101874
transform -1 0 3132 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_360
timestamp 1607101874
transform -1 0 3164 0 1 905
box -2 -3 34 103
use INVX1  INVX1_45
timestamp 1607101874
transform -1 0 3180 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_712
timestamp 1607101874
transform -1 0 3276 0 1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_37
timestamp 1607101874
transform -1 0 3324 0 1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_574
timestamp 1607101874
transform 1 0 3324 0 1 905
box -2 -3 98 103
use FILL  FILL_9_6_0
timestamp 1607101874
transform 1 0 3420 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1607101874
transform 1 0 3428 0 1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_549
timestamp 1607101874
transform 1 0 3436 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_627
timestamp 1607101874
transform 1 0 3460 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_739
timestamp 1607101874
transform -1 0 3516 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_499
timestamp 1607101874
transform -1 0 3540 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_468
timestamp 1607101874
transform 1 0 3540 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_734
timestamp 1607101874
transform 1 0 3572 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_622
timestamp 1607101874
transform -1 0 3628 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_622
timestamp 1607101874
transform 1 0 3628 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_9
timestamp 1607101874
transform 1 0 3724 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1607101874
transform -1 0 3780 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1137
timestamp 1607101874
transform -1 0 3812 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1607101874
transform 1 0 3812 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1607101874
transform -1 0 3932 0 1 905
box -2 -3 98 103
use FILL  FILL_9_7_0
timestamp 1607101874
transform 1 0 3932 0 1 905
box -2 -3 10 103
use FILL  FILL_9_7_1
timestamp 1607101874
transform 1 0 3940 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_125
timestamp 1607101874
transform 1 0 3948 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_643
timestamp 1607101874
transform 1 0 3980 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_8
timestamp 1607101874
transform 1 0 4076 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1607101874
transform -1 0 4132 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_503
timestamp 1607101874
transform -1 0 4156 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_504
timestamp 1607101874
transform 1 0 4156 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_192
timestamp 1607101874
transform 1 0 4180 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_318
timestamp 1607101874
transform -1 0 4228 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_627
timestamp 1607101874
transform -1 0 4260 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1038
timestamp 1607101874
transform -1 0 4292 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1607101874
transform -1 0 4388 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1229
timestamp 1607101874
transform -1 0 4420 0 1 905
box -2 -3 34 103
use FILL  FILL_9_8_0
timestamp 1607101874
transform -1 0 4428 0 1 905
box -2 -3 10 103
use FILL  FILL_9_8_1
timestamp 1607101874
transform -1 0 4436 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_1228
timestamp 1607101874
transform -1 0 4468 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_606
timestamp 1607101874
transform -1 0 4492 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_603
timestamp 1607101874
transform 1 0 4492 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1607101874
transform 1 0 4516 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1144
timestamp 1607101874
transform 1 0 4612 0 1 905
box -2 -3 34 103
use INVX1  INVX1_273
timestamp 1607101874
transform -1 0 4660 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_629
timestamp 1607101874
transform 1 0 4660 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_18
timestamp 1607101874
transform -1 0 4788 0 1 905
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1607101874
transform -1 0 4804 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1234
timestamp 1607101874
transform -1 0 4836 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_561
timestamp 1607101874
transform -1 0 4860 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_493
timestamp 1607101874
transform -1 0 4884 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_279
timestamp 1607101874
transform -1 0 4908 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_182
timestamp 1607101874
transform -1 0 4940 0 1 905
box -2 -3 34 103
use FILL  FILL_9_9_0
timestamp 1607101874
transform -1 0 4948 0 1 905
box -2 -3 10 103
use FILL  FILL_9_9_1
timestamp 1607101874
transform -1 0 4956 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1607101874
transform -1 0 5052 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_654
timestamp 1607101874
transform -1 0 5148 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1607101874
transform -1 0 5244 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_275
timestamp 1607101874
transform -1 0 5268 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_227
timestamp 1607101874
transform -1 0 5292 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1607101874
transform 1 0 5292 0 1 905
box -2 -3 10 103
use FILL  FILL_10_2
timestamp 1607101874
transform 1 0 5300 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_315
timestamp 1607101874
transform 1 0 4 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_299
timestamp 1607101874
transform 1 0 100 0 -1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_285
timestamp 1607101874
transform -1 0 164 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1607101874
transform 1 0 164 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_340
timestamp 1607101874
transform 1 0 260 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1541
timestamp 1607101874
transform 1 0 292 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1607101874
transform 1 0 324 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1607101874
transform 1 0 332 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_734
timestamp 1607101874
transform 1 0 340 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_341
timestamp 1607101874
transform -1 0 404 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1607101874
transform 1 0 404 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_302
timestamp 1607101874
transform 1 0 500 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_554
timestamp 1607101874
transform 1 0 596 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_666
timestamp 1607101874
transform -1 0 652 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_252
timestamp 1607101874
transform 1 0 652 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_179
timestamp 1607101874
transform -1 0 708 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_834
timestamp 1607101874
transform 1 0 708 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_67
timestamp 1607101874
transform -1 0 836 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1607101874
transform 1 0 836 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1607101874
transform 1 0 844 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_308
timestamp 1607101874
transform 1 0 852 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_183
timestamp 1607101874
transform -1 0 972 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_283
timestamp 1607101874
transform -1 0 996 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_892
timestamp 1607101874
transform 1 0 996 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_125
timestamp 1607101874
transform 1 0 1028 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_138
timestamp 1607101874
transform -1 0 1092 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1020
timestamp 1607101874
transform 1 0 1092 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_514
timestamp 1607101874
transform 1 0 1188 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_436
timestamp 1607101874
transform 1 0 1284 0 -1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_384
timestamp 1607101874
transform 1 0 1300 0 -1 1105
box -2 -3 50 103
use FILL  FILL_10_2_0
timestamp 1607101874
transform 1 0 1348 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1607101874
transform 1 0 1356 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_167
timestamp 1607101874
transform 1 0 1364 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_830
timestamp 1607101874
transform 1 0 1396 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_868
timestamp 1607101874
transform 1 0 1492 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_143
timestamp 1607101874
transform 1 0 1588 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_84
timestamp 1607101874
transform -1 0 1644 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_248
timestamp 1607101874
transform -1 0 1676 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_260
timestamp 1607101874
transform 1 0 1676 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_94
timestamp 1607101874
transform 1 0 1708 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_872
timestamp 1607101874
transform -1 0 1852 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1220
timestamp 1607101874
transform 1 0 1852 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_560
timestamp 1607101874
transform 1 0 1900 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_672
timestamp 1607101874
transform -1 0 1956 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_80
timestamp 1607101874
transform 1 0 1956 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_137
timestamp 1607101874
transform -1 0 2012 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_856
timestamp 1607101874
transform 1 0 2012 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_258
timestamp 1607101874
transform 1 0 2108 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_862
timestamp 1607101874
transform 1 0 2132 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_251
timestamp 1607101874
transform 1 0 2164 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_246
timestamp 1607101874
transform 1 0 2196 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_567
timestamp 1607101874
transform 1 0 2228 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1546
timestamp 1607101874
transform 1 0 2324 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1545
timestamp 1607101874
transform -1 0 2388 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_4_0
timestamp 1607101874
transform 1 0 2388 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1607101874
transform 1 0 2396 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_626
timestamp 1607101874
transform 1 0 2404 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_573
timestamp 1607101874
transform 1 0 2436 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_65
timestamp 1607101874
transform -1 0 2564 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_587
timestamp 1607101874
transform 1 0 2564 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1561
timestamp 1607101874
transform 1 0 2660 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1562
timestamp 1607101874
transform -1 0 2724 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1563
timestamp 1607101874
transform 1 0 2724 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1564
timestamp 1607101874
transform -1 0 2788 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_588
timestamp 1607101874
transform 1 0 2788 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_5_0
timestamp 1607101874
transform -1 0 2892 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1607101874
transform -1 0 2900 0 -1 1105
box -2 -3 10 103
use BUFX4  BUFX4_426
timestamp 1607101874
transform -1 0 2932 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_409
timestamp 1607101874
transform -1 0 2980 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_407
timestamp 1607101874
transform 1 0 2980 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_461
timestamp 1607101874
transform -1 0 3044 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_578
timestamp 1607101874
transform 1 0 3044 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_590
timestamp 1607101874
transform -1 0 3236 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1568
timestamp 1607101874
transform 1 0 3236 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1567
timestamp 1607101874
transform -1 0 3300 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1132
timestamp 1607101874
transform 1 0 3300 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1134
timestamp 1607101874
transform -1 0 3364 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_551
timestamp 1607101874
transform 1 0 3364 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_6_0
timestamp 1607101874
transform 1 0 3388 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1607101874
transform 1 0 3396 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_582
timestamp 1607101874
transform 1 0 3404 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_64
timestamp 1607101874
transform -1 0 3532 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1135
timestamp 1607101874
transform 1 0 3532 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_63
timestamp 1607101874
transform -1 0 3604 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_554
timestamp 1607101874
transform 1 0 3604 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1140
timestamp 1607101874
transform -1 0 3660 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_61
timestamp 1607101874
transform -1 0 3700 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_552
timestamp 1607101874
transform -1 0 3724 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_553
timestamp 1607101874
transform -1 0 3748 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_476
timestamp 1607101874
transform 1 0 3748 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_363
timestamp 1607101874
transform -1 0 3804 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_594
timestamp 1607101874
transform -1 0 3900 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_3
timestamp 1607101874
transform 1 0 3900 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_7_0
timestamp 1607101874
transform -1 0 3932 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_7_1
timestamp 1607101874
transform -1 0 3940 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_1
timestamp 1607101874
transform -1 0 3972 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_372
timestamp 1607101874
transform -1 0 4004 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_634
timestamp 1607101874
transform -1 0 4028 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_522
timestamp 1607101874
transform -1 0 4060 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_274
timestamp 1607101874
transform -1 0 4108 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_360
timestamp 1607101874
transform -1 0 4124 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_319
timestamp 1607101874
transform 1 0 4124 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_447
timestamp 1607101874
transform -1 0 4180 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1607101874
transform 1 0 4180 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1039
timestamp 1607101874
transform -1 0 4236 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_291
timestamp 1607101874
transform -1 0 4268 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_591
timestamp 1607101874
transform -1 0 4364 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_361
timestamp 1607101874
transform 1 0 4364 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1569
timestamp 1607101874
transform -1 0 4420 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_8_0
timestamp 1607101874
transform 1 0 4420 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_8_1
timestamp 1607101874
transform 1 0 4428 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1607101874
transform 1 0 4436 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_33
timestamp 1607101874
transform -1 0 4556 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_371
timestamp 1607101874
transform 1 0 4556 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1607101874
transform -1 0 4612 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1145
timestamp 1607101874
transform -1 0 4644 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_64
timestamp 1607101874
transform -1 0 4684 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_33
timestamp 1607101874
transform 1 0 4684 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1607101874
transform -1 0 4748 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_650
timestamp 1607101874
transform -1 0 4844 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_25
timestamp 1607101874
transform 1 0 4844 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_7
timestamp 1607101874
transform -1 0 4900 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_9_0
timestamp 1607101874
transform -1 0 4908 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_9_1
timestamp 1607101874
transform -1 0 4916 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_637
timestamp 1607101874
transform -1 0 5012 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_639
timestamp 1607101874
transform -1 0 5108 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_36
timestamp 1607101874
transform 1 0 5108 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_395
timestamp 1607101874
transform 1 0 5124 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_164
timestamp 1607101874
transform 1 0 5156 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1607101874
transform -1 0 5300 0 -1 1105
box -2 -3 98 103
use FILL  FILL_11_1
timestamp 1607101874
transform -1 0 5308 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1607101874
transform 1 0 4 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_337
timestamp 1607101874
transform -1 0 132 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_336
timestamp 1607101874
transform -1 0 164 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_208
timestamp 1607101874
transform 1 0 164 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_343
timestamp 1607101874
transform -1 0 220 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_342
timestamp 1607101874
transform 1 0 220 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_308
timestamp 1607101874
transform 1 0 252 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1607101874
transform -1 0 380 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_0_0
timestamp 1607101874
transform 1 0 380 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1607101874
transform 1 0 388 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_339
timestamp 1607101874
transform 1 0 396 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_338
timestamp 1607101874
transform 1 0 428 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1607101874
transform 1 0 460 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_146
timestamp 1607101874
transform 1 0 556 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_133
timestamp 1607101874
transform -1 0 620 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_394
timestamp 1607101874
transform 1 0 620 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_887
timestamp 1607101874
transform 1 0 668 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_267
timestamp 1607101874
transform 1 0 700 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_75
timestamp 1607101874
transform 1 0 724 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_129
timestamp 1607101874
transform -1 0 780 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_226
timestamp 1607101874
transform -1 0 828 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_1026
timestamp 1607101874
transform 1 0 828 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1607101874
transform 1 0 860 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1607101874
transform 1 0 868 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_1363
timestamp 1607101874
transform 1 0 876 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1362
timestamp 1607101874
transform 1 0 908 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_372
timestamp 1607101874
transform 1 0 940 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_948
timestamp 1607101874
transform 1 0 956 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_227
timestamp 1607101874
transform -1 0 1036 0 1 1105
box -2 -3 50 103
use BUFX4  BUFX4_454
timestamp 1607101874
transform -1 0 1068 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_557
timestamp 1607101874
transform 1 0 1068 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_669
timestamp 1607101874
transform -1 0 1124 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_305
timestamp 1607101874
transform 1 0 1124 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_439
timestamp 1607101874
transform 1 0 1220 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_338
timestamp 1607101874
transform -1 0 1276 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1166
timestamp 1607101874
transform -1 0 1308 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_259
timestamp 1607101874
transform 1 0 1308 0 1 1105
box -2 -3 50 103
use FILL  FILL_11_2_0
timestamp 1607101874
transform 1 0 1356 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1607101874
transform 1 0 1364 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_1120
timestamp 1607101874
transform 1 0 1372 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_166
timestamp 1607101874
transform 1 0 1404 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1214
timestamp 1607101874
transform -1 0 1468 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_593
timestamp 1607101874
transform 1 0 1468 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_77
timestamp 1607101874
transform -1 0 1532 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_594
timestamp 1607101874
transform 1 0 1532 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_330
timestamp 1607101874
transform -1 0 1588 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_325
timestamp 1607101874
transform -1 0 1620 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_732
timestamp 1607101874
transform 1 0 1620 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_57
timestamp 1607101874
transform 1 0 1716 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_107
timestamp 1607101874
transform -1 0 1748 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_262
timestamp 1607101874
transform -1 0 1780 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_273
timestamp 1607101874
transform 1 0 1780 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_221
timestamp 1607101874
transform -1 0 1844 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_257
timestamp 1607101874
transform -1 0 1876 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_3_0
timestamp 1607101874
transform 1 0 1876 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1607101874
transform 1 0 1884 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1607101874
transform 1 0 1892 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_441
timestamp 1607101874
transform -1 0 2020 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_269
timestamp 1607101874
transform -1 0 2052 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_596
timestamp 1607101874
transform 1 0 2052 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_595
timestamp 1607101874
transform 1 0 2076 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_80
timestamp 1607101874
transform -1 0 2140 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_597
timestamp 1607101874
transform 1 0 2140 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_78
timestamp 1607101874
transform -1 0 2204 0 1 1105
box -2 -3 42 103
use BUFX4  BUFX4_21
timestamp 1607101874
transform -1 0 2236 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1607101874
transform -1 0 2268 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_687
timestamp 1607101874
transform 1 0 2268 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_308
timestamp 1607101874
transform -1 0 2332 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_570
timestamp 1607101874
transform 1 0 2332 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_4_0
timestamp 1607101874
transform 1 0 2428 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1607101874
transform 1 0 2436 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_1552
timestamp 1607101874
transform 1 0 2444 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1551
timestamp 1607101874
transform -1 0 2508 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_738
timestamp 1607101874
transform -1 0 2532 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_294
timestamp 1607101874
transform -1 0 2556 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1024
timestamp 1607101874
transform 1 0 2556 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_321
timestamp 1607101874
transform 1 0 2588 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_579
timestamp 1607101874
transform 1 0 2620 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_271
timestamp 1607101874
transform 1 0 2716 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_408
timestamp 1607101874
transform -1 0 2780 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_617
timestamp 1607101874
transform -1 0 2812 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_287
timestamp 1607101874
transform -1 0 2844 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_826
timestamp 1607101874
transform -1 0 2876 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_618
timestamp 1607101874
transform -1 0 2908 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_5_0
timestamp 1607101874
transform 1 0 2908 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1607101874
transform 1 0 2916 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_288
timestamp 1607101874
transform 1 0 2924 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_797
timestamp 1607101874
transform 1 0 2956 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_350
timestamp 1607101874
transform -1 0 3020 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_798
timestamp 1607101874
transform 1 0 3020 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1607101874
transform 1 0 3052 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1023
timestamp 1607101874
transform -1 0 3108 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_825
timestamp 1607101874
transform -1 0 3140 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_439
timestamp 1607101874
transform 1 0 3140 0 1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_72
timestamp 1607101874
transform 1 0 3172 0 1 1105
box -2 -3 74 103
use OAI21X1  OAI21X1_1022
timestamp 1607101874
transform -1 0 3276 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1130
timestamp 1607101874
transform 1 0 3276 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1607101874
transform -1 0 3332 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_479
timestamp 1607101874
transform -1 0 3364 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_411
timestamp 1607101874
transform 1 0 3364 0 1 1105
box -2 -3 50 103
use FILL  FILL_11_6_0
timestamp 1607101874
transform -1 0 3420 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1607101874
transform -1 0 3428 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_425
timestamp 1607101874
transform -1 0 3444 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_1131
timestamp 1607101874
transform 1 0 3444 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_550
timestamp 1607101874
transform -1 0 3500 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1129
timestamp 1607101874
transform 1 0 3500 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1185
timestamp 1607101874
transform -1 0 3564 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_4
timestamp 1607101874
transform 1 0 3564 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_7
timestamp 1607101874
transform -1 0 3628 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_1136
timestamp 1607101874
transform -1 0 3660 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_598
timestamp 1607101874
transform -1 0 3756 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_280
timestamp 1607101874
transform -1 0 3780 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_314
timestamp 1607101874
transform 1 0 3780 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_28
timestamp 1607101874
transform -1 0 3844 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1607101874
transform -1 0 3860 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_615
timestamp 1607101874
transform -1 0 3956 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_7_0
timestamp 1607101874
transform 1 0 3956 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_7_1
timestamp 1607101874
transform 1 0 3964 0 1 1105
box -2 -3 10 103
use BUFX4  BUFX4_323
timestamp 1607101874
transform 1 0 3972 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_932
timestamp 1607101874
transform 1 0 4004 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_384
timestamp 1607101874
transform -1 0 4132 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1042
timestamp 1607101874
transform -1 0 4164 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_404
timestamp 1607101874
transform 1 0 4164 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1607101874
transform -1 0 4292 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_346
timestamp 1607101874
transform 1 0 4292 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_452
timestamp 1607101874
transform -1 0 4348 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_72
timestamp 1607101874
transform 1 0 4348 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1607101874
transform -1 0 4412 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_8_0
timestamp 1607101874
transform 1 0 4412 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_8_1
timestamp 1607101874
transform 1 0 4420 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_625
timestamp 1607101874
transform 1 0 4428 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_14
timestamp 1607101874
transform -1 0 4556 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1607101874
transform -1 0 4588 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_506
timestamp 1607101874
transform -1 0 4620 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1231
timestamp 1607101874
transform -1 0 4652 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_81
timestamp 1607101874
transform -1 0 4684 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1607101874
transform 1 0 4684 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_1
timestamp 1607101874
transform -1 0 4748 0 1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_560
timestamp 1607101874
transform -1 0 4772 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_642
timestamp 1607101874
transform -1 0 4868 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_25
timestamp 1607101874
transform -1 0 4900 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1607101874
transform -1 0 4932 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_286
timestamp 1607101874
transform -1 0 4956 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_9_0
timestamp 1607101874
transform -1 0 4964 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_9_1
timestamp 1607101874
transform -1 0 4972 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_189
timestamp 1607101874
transform -1 0 5004 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1607101874
transform -1 0 5100 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_19
timestamp 1607101874
transform -1 0 5132 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1607101874
transform -1 0 5164 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_145
timestamp 1607101874
transform 1 0 5164 0 1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1607101874
transform -1 0 5308 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_543
timestamp 1607101874
transform 1 0 4 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1530
timestamp 1607101874
transform -1 0 132 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1529
timestamp 1607101874
transform -1 0 164 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_84
timestamp 1607101874
transform -1 0 188 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_262
timestamp 1607101874
transform 1 0 188 0 -1 1305
box -2 -3 18 103
use BUFX4  BUFX4_309
timestamp 1607101874
transform -1 0 236 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_48
timestamp 1607101874
transform -1 0 284 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_58
timestamp 1607101874
transform -1 0 300 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_0_0
timestamp 1607101874
transform -1 0 308 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1607101874
transform -1 0 316 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_733
timestamp 1607101874
transform -1 0 412 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_343
timestamp 1607101874
transform 1 0 412 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_544
timestamp 1607101874
transform -1 0 540 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_551
timestamp 1607101874
transform 1 0 540 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_263
timestamp 1607101874
transform 1 0 636 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_833
timestamp 1607101874
transform 1 0 652 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_74
timestamp 1607101874
transform 1 0 748 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1607101874
transform -1 0 804 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_399
timestamp 1607101874
transform 1 0 804 0 -1 1305
box -2 -3 18 103
use BUFX4  BUFX4_381
timestamp 1607101874
transform -1 0 852 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1607101874
transform 1 0 852 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1607101874
transform 1 0 860 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_305
timestamp 1607101874
transform 1 0 868 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1025
timestamp 1607101874
transform 1 0 892 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1027
timestamp 1607101874
transform -1 0 956 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_607
timestamp 1607101874
transform 1 0 956 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_185
timestamp 1607101874
transform -1 0 1020 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_284
timestamp 1607101874
transform -1 0 1044 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_164
timestamp 1607101874
transform 1 0 1044 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_165
timestamp 1607101874
transform -1 0 1108 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_829
timestamp 1607101874
transform 1 0 1108 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_309
timestamp 1607101874
transform 1 0 1204 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1365
timestamp 1607101874
transform 1 0 1300 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1364
timestamp 1607101874
transform -1 0 1364 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_2_0
timestamp 1607101874
transform -1 0 1372 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1607101874
transform -1 0 1380 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_542
timestamp 1607101874
transform -1 0 1404 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_57
timestamp 1607101874
transform -1 0 1444 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_543
timestamp 1607101874
transform 1 0 1444 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_262
timestamp 1607101874
transform 1 0 1468 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_86
timestamp 1607101874
transform -1 0 1540 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_137
timestamp 1607101874
transform 1 0 1540 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_120
timestamp 1607101874
transform -1 0 1604 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1607101874
transform 1 0 1604 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_186
timestamp 1607101874
transform 1 0 1652 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_187
timestamp 1607101874
transform -1 0 1716 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_864
timestamp 1607101874
transform -1 0 1812 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_509
timestamp 1607101874
transform 1 0 1812 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_546
timestamp 1607101874
transform -1 0 1868 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_3_0
timestamp 1607101874
transform -1 0 1876 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1607101874
transform -1 0 1884 0 -1 1305
box -2 -3 10 103
use INVX8  INVX8_20
timestamp 1607101874
transform -1 0 1924 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_56
timestamp 1607101874
transform 1 0 1924 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_128
timestamp 1607101874
transform 1 0 1948 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_171
timestamp 1607101874
transform 1 0 1980 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_170
timestamp 1607101874
transform 1 0 2012 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_844
timestamp 1607101874
transform 1 0 2044 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_854
timestamp 1607101874
transform 1 0 2140 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_183
timestamp 1607101874
transform 1 0 2236 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_182
timestamp 1607101874
transform -1 0 2300 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_337
timestamp 1607101874
transform 1 0 2300 0 -1 1305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_5
timestamp 1607101874
transform -1 0 2388 0 -1 1305
box -2 -3 74 103
use FILL  FILL_12_4_0
timestamp 1607101874
transform 1 0 2388 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1607101874
transform 1 0 2396 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_268
timestamp 1607101874
transform 1 0 2404 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_172
timestamp 1607101874
transform -1 0 2460 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_349
timestamp 1607101874
transform 1 0 2460 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_390
timestamp 1607101874
transform 1 0 2492 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_972
timestamp 1607101874
transform 1 0 2508 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_348
timestamp 1607101874
transform 1 0 2540 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1607101874
transform 1 0 2572 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_403
timestamp 1607101874
transform 1 0 2668 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1057
timestamp 1607101874
transform 1 0 2684 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1607101874
transform -1 0 2740 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_250
timestamp 1607101874
transform -1 0 2788 0 -1 1305
box -2 -3 50 103
use CLKBUF1  CLKBUF1_25
timestamp 1607101874
transform 1 0 2788 0 -1 1305
box -2 -3 74 103
use BUFX4  BUFX4_195
timestamp 1607101874
transform -1 0 2892 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_5_0
timestamp 1607101874
transform 1 0 2892 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1607101874
transform 1 0 2900 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_356
timestamp 1607101874
transform 1 0 2908 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_357
timestamp 1607101874
transform -1 0 2972 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1607101874
transform 1 0 2972 0 -1 1305
box -2 -3 98 103
use BUFX4  BUFX4_196
timestamp 1607101874
transform 1 0 3068 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_389
timestamp 1607101874
transform -1 0 3116 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_561
timestamp 1607101874
transform -1 0 3212 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_400
timestamp 1607101874
transform 1 0 3212 0 -1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_292
timestamp 1607101874
transform -1 0 3292 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_405
timestamp 1607101874
transform -1 0 3316 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_402
timestamp 1607101874
transform 1 0 3316 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1607101874
transform 1 0 3340 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_6_0
timestamp 1607101874
transform 1 0 3436 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1607101874
transform 1 0 3444 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_174
timestamp 1607101874
transform 1 0 3452 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_161
timestamp 1607101874
transform -1 0 3516 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_566
timestamp 1607101874
transform 1 0 3516 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1607101874
transform 1 0 3612 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_6
timestamp 1607101874
transform 1 0 3708 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1607101874
transform -1 0 3764 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_619
timestamp 1607101874
transform -1 0 3796 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_289
timestamp 1607101874
transform -1 0 3828 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_376
timestamp 1607101874
transform 1 0 3828 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1607101874
transform -1 0 3884 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_17
timestamp 1607101874
transform -1 0 3932 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_7_0
timestamp 1607101874
transform 1 0 3932 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_7_1
timestamp 1607101874
transform 1 0 3940 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1607101874
transform 1 0 3948 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_294
timestamp 1607101874
transform 1 0 4044 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_450
timestamp 1607101874
transform 1 0 4076 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_442
timestamp 1607101874
transform -1 0 4140 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_611
timestamp 1607101874
transform 1 0 4140 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_18
timestamp 1607101874
transform 1 0 4236 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_13
timestamp 1607101874
transform -1 0 4300 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_620
timestamp 1607101874
transform 1 0 4300 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_624
timestamp 1607101874
transform 1 0 4332 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_621
timestamp 1607101874
transform 1 0 4364 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1232
timestamp 1607101874
transform 1 0 4396 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_8_0
timestamp 1607101874
transform 1 0 4428 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_8_1
timestamp 1607101874
transform 1 0 4436 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_296
timestamp 1607101874
transform 1 0 4444 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1607101874
transform -1 0 4572 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_369
timestamp 1607101874
transform 1 0 4572 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_189
timestamp 1607101874
transform -1 0 4628 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_438
timestamp 1607101874
transform 1 0 4628 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_595
timestamp 1607101874
transform -1 0 4756 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_627
timestamp 1607101874
transform -1 0 4852 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_17
timestamp 1607101874
transform 1 0 4852 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_1
timestamp 1607101874
transform -1 0 4908 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_204
timestamp 1607101874
transform 1 0 4908 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_9_0
timestamp 1607101874
transform -1 0 4940 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_9_1
timestamp 1607101874
transform -1 0 4948 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_644
timestamp 1607101874
transform -1 0 5044 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_389
timestamp 1607101874
transform 1 0 5044 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_390
timestamp 1607101874
transform -1 0 5108 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1607101874
transform -1 0 5204 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1607101874
transform -1 0 5300 0 -1 1305
box -2 -3 98 103
use FILL  FILL_13_1
timestamp 1607101874
transform -1 0 5308 0 -1 1305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_92
timestamp 1607101874
transform -1 0 76 0 1 1305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_741
timestamp 1607101874
transform 1 0 76 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_98
timestamp 1607101874
transform 1 0 172 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1607101874
transform -1 0 236 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_322
timestamp 1607101874
transform -1 0 268 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1300
timestamp 1607101874
transform 1 0 268 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1607101874
transform -1 0 308 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1607101874
transform -1 0 316 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1607101874
transform -1 0 412 0 1 1305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_90
timestamp 1607101874
transform -1 0 484 0 1 1305
box -2 -3 74 103
use INVX1  INVX1_322
timestamp 1607101874
transform 1 0 484 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1532
timestamp 1607101874
transform -1 0 532 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1301
timestamp 1607101874
transform -1 0 564 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_555
timestamp 1607101874
transform 1 0 564 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_745
timestamp 1607101874
transform 1 0 660 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_106
timestamp 1607101874
transform 1 0 756 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1607101874
transform -1 0 820 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1607101874
transform 1 0 820 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1607101874
transform 1 0 828 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_832
timestamp 1607101874
transform 1 0 836 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_127
timestamp 1607101874
transform 1 0 932 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_73
timestamp 1607101874
transform -1 0 988 0 1 1305
box -2 -3 34 103
use AND2X2  AND2X2_45
timestamp 1607101874
transform -1 0 1020 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_949
timestamp 1607101874
transform -1 0 1052 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_233
timestamp 1607101874
transform 1 0 1052 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_184
timestamp 1607101874
transform -1 0 1124 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_608
timestamp 1607101874
transform 1 0 1124 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1008
timestamp 1607101874
transform -1 0 1188 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_396
timestamp 1607101874
transform -1 0 1204 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_183
timestamp 1607101874
transform -1 0 1252 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_180
timestamp 1607101874
transform 1 0 1252 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_163
timestamp 1607101874
transform 1 0 1284 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1607101874
transform -1 0 1348 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_2_0
timestamp 1607101874
transform -1 0 1356 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1607101874
transform -1 0 1364 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_828
timestamp 1607101874
transform -1 0 1460 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_317
timestamp 1607101874
transform 1 0 1460 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_413
timestamp 1607101874
transform 1 0 1556 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_161
timestamp 1607101874
transform 1 0 1572 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_160
timestamp 1607101874
transform 1 0 1604 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_117
timestamp 1607101874
transform -1 0 1660 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_186
timestamp 1607101874
transform -1 0 1692 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_827
timestamp 1607101874
transform 1 0 1692 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_244
timestamp 1607101874
transform 1 0 1788 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_93
timestamp 1607101874
transform -1 0 1852 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_3_0
timestamp 1607101874
transform 1 0 1852 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1607101874
transform 1 0 1860 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_835
timestamp 1607101874
transform 1 0 1868 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_860
timestamp 1607101874
transform 1 0 1964 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_257
timestamp 1607101874
transform 1 0 1996 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_831
timestamp 1607101874
transform 1 0 2020 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_287
timestamp 1607101874
transform 1 0 2052 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1369
timestamp 1607101874
transform 1 0 2148 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1368
timestamp 1607101874
transform 1 0 2180 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1217
timestamp 1607101874
transform -1 0 2244 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_424
timestamp 1607101874
transform -1 0 2268 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_425
timestamp 1607101874
transform 1 0 2268 0 1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_21
timestamp 1607101874
transform 1 0 2292 0 1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_220
timestamp 1607101874
transform 1 0 2332 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_4_0
timestamp 1607101874
transform 1 0 2380 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1607101874
transform 1 0 2388 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_863
timestamp 1607101874
transform 1 0 2396 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_472
timestamp 1607101874
transform 1 0 2428 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1377
timestamp 1607101874
transform 1 0 2460 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1376
timestamp 1607101874
transform 1 0 2492 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_765
timestamp 1607101874
transform -1 0 2556 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1549
timestamp 1607101874
transform 1 0 2556 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1550
timestamp 1607101874
transform 1 0 2588 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_569
timestamp 1607101874
transform -1 0 2716 0 1 1305
box -2 -3 98 103
use BUFX4  BUFX4_385
timestamp 1607101874
transform -1 0 2748 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_271
timestamp 1607101874
transform -1 0 2844 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1607101874
transform 1 0 2844 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_5_0
timestamp 1607101874
transform 1 0 2940 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1607101874
transform 1 0 2948 0 1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_251
timestamp 1607101874
transform 1 0 2956 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_239
timestamp 1607101874
transform -1 0 3052 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_971
timestamp 1607101874
transform -1 0 3084 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_198
timestamp 1607101874
transform 1 0 3084 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1560
timestamp 1607101874
transform 1 0 3116 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1559
timestamp 1607101874
transform 1 0 3148 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_586
timestamp 1607101874
transform 1 0 3180 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_404
timestamp 1607101874
transform 1 0 3276 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1059
timestamp 1607101874
transform 1 0 3292 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1133
timestamp 1607101874
transform 1 0 3324 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_365
timestamp 1607101874
transform 1 0 3356 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_364
timestamp 1607101874
transform 1 0 3388 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_6_0
timestamp 1607101874
transform -1 0 3428 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1607101874
transform -1 0 3436 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_325
timestamp 1607101874
transform -1 0 3460 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1607101874
transform -1 0 3556 0 1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_478
timestamp 1607101874
transform -1 0 3588 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_424
timestamp 1607101874
transform 1 0 3588 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_403
timestamp 1607101874
transform -1 0 3652 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_173
timestamp 1607101874
transform 1 0 3652 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_602
timestamp 1607101874
transform -1 0 3708 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_269
timestamp 1607101874
transform 1 0 3708 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_31
timestamp 1607101874
transform 1 0 3732 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1227
timestamp 1607101874
transform 1 0 3756 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_504
timestamp 1607101874
transform 1 0 3788 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_173
timestamp 1607101874
transform 1 0 3820 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_619
timestamp 1607101874
transform -1 0 3948 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_7_0
timestamp 1607101874
transform -1 0 3956 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_7_1
timestamp 1607101874
transform -1 0 3964 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1607101874
transform -1 0 4060 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_23
timestamp 1607101874
transform 1 0 4060 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_633
timestamp 1607101874
transform 1 0 4108 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_30
timestamp 1607101874
transform 1 0 4204 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_430
timestamp 1607101874
transform 1 0 4220 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_16
timestamp 1607101874
transform -1 0 4276 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_146
timestamp 1607101874
transform 1 0 4276 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_159
timestamp 1607101874
transform -1 0 4340 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1607101874
transform -1 0 4436 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_8_0
timestamp 1607101874
transform -1 0 4444 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_8_1
timestamp 1607101874
transform -1 0 4452 0 1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_455
timestamp 1607101874
transform -1 0 4476 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_22
timestamp 1607101874
transform -1 0 4500 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_982
timestamp 1607101874
transform -1 0 4532 0 1 1305
box -2 -3 34 103
use INVX8  INVX8_5
timestamp 1607101874
transform 1 0 4532 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_87
timestamp 1607101874
transform 1 0 4572 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_190
timestamp 1607101874
transform -1 0 4620 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1146
timestamp 1607101874
transform -1 0 4652 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_213
timestamp 1607101874
transform 1 0 4652 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_984
timestamp 1607101874
transform -1 0 4716 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_490
timestamp 1607101874
transform -1 0 4740 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_983
timestamp 1607101874
transform -1 0 4772 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_217
timestamp 1607101874
transform 1 0 4772 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_649
timestamp 1607101874
transform -1 0 4916 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_32
timestamp 1607101874
transform 1 0 4916 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_9_0
timestamp 1607101874
transform -1 0 4956 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_9_1
timestamp 1607101874
transform -1 0 4964 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_31
timestamp 1607101874
transform -1 0 4996 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_815
timestamp 1607101874
transform 1 0 4996 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_29
timestamp 1607101874
transform 1 0 5028 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_817
timestamp 1607101874
transform 1 0 5052 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_9
timestamp 1607101874
transform -1 0 5116 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_292
timestamp 1607101874
transform 1 0 5116 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_397
timestamp 1607101874
transform 1 0 5148 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_398
timestamp 1607101874
transform -1 0 5212 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1607101874
transform 1 0 5212 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1607101874
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1291
timestamp 1607101874
transform -1 0 132 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1290
timestamp 1607101874
transform -1 0 164 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_225
timestamp 1607101874
transform 1 0 164 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_255
timestamp 1607101874
transform -1 0 204 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1607101874
transform 1 0 204 0 -1 1505
box -2 -3 98 103
use AND2X2  AND2X2_28
timestamp 1607101874
transform 1 0 300 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_0_0
timestamp 1607101874
transform -1 0 340 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1607101874
transform -1 0 348 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_736
timestamp 1607101874
transform -1 0 380 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1537
timestamp 1607101874
transform 1 0 380 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1538
timestamp 1607101874
transform -1 0 444 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1531
timestamp 1607101874
transform 1 0 444 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_787
timestamp 1607101874
transform -1 0 508 0 -1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_48
timestamp 1607101874
transform 1 0 508 0 -1 1505
box -2 -3 74 103
use AND2X2  AND2X2_21
timestamp 1607101874
transform 1 0 580 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_560
timestamp 1607101874
transform 1 0 612 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_301
timestamp 1607101874
transform 1 0 644 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_323
timestamp 1607101874
transform -1 0 788 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_454
timestamp 1607101874
transform 1 0 788 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_324
timestamp 1607101874
transform -1 0 852 0 -1 1505
box -2 -3 50 103
use FILL  FILL_14_1_0
timestamp 1607101874
transform 1 0 852 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1607101874
transform 1 0 860 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_440
timestamp 1607101874
transform 1 0 868 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_377
timestamp 1607101874
transform 1 0 900 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_812
timestamp 1607101874
transform 1 0 932 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_91
timestamp 1607101874
transform 1 0 1028 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_142
timestamp 1607101874
transform 1 0 1044 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_49
timestamp 1607101874
transform -1 0 1100 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_858
timestamp 1607101874
transform 1 0 1100 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_513
timestamp 1607101874
transform 1 0 1132 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_383
timestamp 1607101874
transform 1 0 1228 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_383
timestamp 1607101874
transform 1 0 1244 0 -1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_378
timestamp 1607101874
transform -1 0 1324 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1121
timestamp 1607101874
transform 1 0 1324 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_2_0
timestamp 1607101874
transform 1 0 1356 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1607101874
transform 1 0 1364 0 -1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_395
timestamp 1607101874
transform 1 0 1372 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_287
timestamp 1607101874
transform -1 0 1452 0 -1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_307
timestamp 1607101874
transform 1 0 1452 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_679
timestamp 1607101874
transform -1 0 1516 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_80
timestamp 1607101874
transform -1 0 1564 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_861
timestamp 1607101874
transform 1 0 1564 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_740
timestamp 1607101874
transform 1 0 1596 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_379
timestamp 1607101874
transform -1 0 1724 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1607101874
transform 1 0 1724 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1607101874
transform -1 0 1788 0 -1 1505
box -2 -3 34 103
use INVX8  INVX8_13
timestamp 1607101874
transform 1 0 1788 0 -1 1505
box -2 -3 42 103
use BUFX4  BUFX4_214
timestamp 1607101874
transform -1 0 1860 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1607101874
transform 1 0 1860 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1607101874
transform 1 0 1868 0 -1 1505
box -2 -3 10 103
use AND2X2  AND2X2_31
timestamp 1607101874
transform 1 0 1876 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_179
timestamp 1607101874
transform -1 0 1940 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_380
timestamp 1607101874
transform -1 0 1972 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_221
timestamp 1607101874
transform -1 0 2020 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_832
timestamp 1607101874
transform 1 0 2020 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_179
timestamp 1607101874
transform 1 0 2052 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1607101874
transform -1 0 2116 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_568
timestamp 1607101874
transform -1 0 2212 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1548
timestamp 1607101874
transform -1 0 2244 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1547
timestamp 1607101874
transform -1 0 2276 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1607101874
transform 1 0 2276 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_350
timestamp 1607101874
transform 1 0 2308 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_4_0
timestamp 1607101874
transform 1 0 2340 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1607101874
transform 1 0 2348 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1607101874
transform 1 0 2356 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_573
timestamp 1607101874
transform 1 0 2452 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_199
timestamp 1607101874
transform -1 0 2508 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_623
timestamp 1607101874
transform 1 0 2508 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_735
timestamp 1607101874
transform -1 0 2564 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_565
timestamp 1607101874
transform 1 0 2564 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_473
timestamp 1607101874
transform -1 0 2692 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_171
timestamp 1607101874
transform 1 0 2692 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_267
timestamp 1607101874
transform -1 0 2748 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_355
timestamp 1607101874
transform 1 0 2748 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1607101874
transform 1 0 2780 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_354
timestamp 1607101874
transform -1 0 2908 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_5_0
timestamp 1607101874
transform -1 0 2916 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1607101874
transform -1 0 2924 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_260
timestamp 1607101874
transform -1 0 2948 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_252
timestamp 1607101874
transform 1 0 2948 0 -1 1505
box -2 -3 50 103
use NOR2X1  NOR2X1_265
timestamp 1607101874
transform -1 0 3020 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1607101874
transform 1 0 3020 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_367
timestamp 1607101874
transform 1 0 3116 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_366
timestamp 1607101874
transform -1 0 3180 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1607101874
transform 1 0 3180 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_178
timestamp 1607101874
transform 1 0 3276 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_259
timestamp 1607101874
transform -1 0 3332 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_165
timestamp 1607101874
transform -1 0 3364 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_6_0
timestamp 1607101874
transform 1 0 3364 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1607101874
transform 1 0 3372 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1607101874
transform 1 0 3380 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_169
timestamp 1607101874
transform 1 0 3476 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_264
timestamp 1607101874
transform -1 0 3532 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1607101874
transform 1 0 3532 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_379
timestamp 1607101874
transform 1 0 3628 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_97
timestamp 1607101874
transform -1 0 3684 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_572
timestamp 1607101874
transform -1 0 3780 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_377
timestamp 1607101874
transform 1 0 3780 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_95
timestamp 1607101874
transform -1 0 3836 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_265
timestamp 1607101874
transform 1 0 3836 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_378
timestamp 1607101874
transform 1 0 3860 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_96
timestamp 1607101874
transform -1 0 3916 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_7_0
timestamp 1607101874
transform 1 0 3916 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_7_1
timestamp 1607101874
transform 1 0 3924 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1607101874
transform 1 0 3932 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_634
timestamp 1607101874
transform 1 0 4028 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1607101874
transform -1 0 4156 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_392
timestamp 1607101874
transform -1 0 4188 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_391
timestamp 1607101874
transform -1 0 4220 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1607101874
transform -1 0 4316 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_160
timestamp 1607101874
transform 1 0 4316 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_147
timestamp 1607101874
transform -1 0 4380 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_626
timestamp 1607101874
transform -1 0 4412 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_8_0
timestamp 1607101874
transform 1 0 4412 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_8_1
timestamp 1607101874
transform 1 0 4420 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_21
timestamp 1607101874
transform 1 0 4428 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_28
timestamp 1607101874
transform -1 0 4492 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_631
timestamp 1607101874
transform -1 0 4588 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_143
timestamp 1607101874
transform 1 0 4588 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_156
timestamp 1607101874
transform -1 0 4652 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1607101874
transform -1 0 4748 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_986
timestamp 1607101874
transform -1 0 4780 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_40
timestamp 1607101874
transform 1 0 4780 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_492
timestamp 1607101874
transform -1 0 4844 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_10
timestamp 1607101874
transform 1 0 4844 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_23
timestamp 1607101874
transform 1 0 4876 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1607101874
transform -1 0 4940 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_9_0
timestamp 1607101874
transform -1 0 4948 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_9_1
timestamp 1607101874
transform -1 0 4956 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_641
timestamp 1607101874
transform -1 0 5052 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_649
timestamp 1607101874
transform 1 0 5052 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1607101874
transform -1 0 5100 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_443
timestamp 1607101874
transform -1 0 5124 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1607101874
transform 1 0 5124 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_162
timestamp 1607101874
transform 1 0 5156 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1607101874
transform -1 0 5300 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1607101874
transform -1 0 5308 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1607101874
transform 1 0 4 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1293
timestamp 1607101874
transform -1 0 132 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_558
timestamp 1607101874
transform 1 0 4 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1544
timestamp 1607101874
transform -1 0 132 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1292
timestamp 1607101874
transform -1 0 164 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_300
timestamp 1607101874
transform 1 0 164 0 1 1505
box -2 -3 18 103
use BUFX4  BUFX4_312
timestamp 1607101874
transform -1 0 212 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1543
timestamp 1607101874
transform -1 0 164 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1536
timestamp 1607101874
transform 1 0 164 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1535
timestamp 1607101874
transform -1 0 228 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1607101874
transform 1 0 212 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1607101874
transform 1 0 244 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_476
timestamp 1607101874
transform -1 0 308 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_739
timestamp 1607101874
transform 1 0 228 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_45
timestamp 1607101874
transform 1 0 340 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_0_1
timestamp 1607101874
transform 1 0 332 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_0
timestamp 1607101874
transform 1 0 324 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1607101874
transform -1 0 340 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_0
timestamp 1607101874
transform -1 0 332 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_226
timestamp 1607101874
transform 1 0 308 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1539
timestamp 1607101874
transform 1 0 396 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_85
timestamp 1607101874
transform -1 0 396 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_735
timestamp 1607101874
transform 1 0 388 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_288
timestamp 1607101874
transform -1 0 388 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_1540
timestamp 1607101874
transform -1 0 452 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_194
timestamp 1607101874
transform -1 0 484 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1607101874
transform 1 0 484 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_556
timestamp 1607101874
transform 1 0 428 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1299
timestamp 1607101874
transform 1 0 580 0 1 1505
box -2 -3 34 103
use AND2X2  AND2X2_30
timestamp 1607101874
transform -1 0 556 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_189
timestamp 1607101874
transform -1 0 588 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1607101874
transform -1 0 620 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_562
timestamp 1607101874
transform 1 0 612 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_561
timestamp 1607101874
transform 1 0 644 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_478
timestamp 1607101874
transform -1 0 708 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_300
timestamp 1607101874
transform 1 0 708 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1298
timestamp 1607101874
transform -1 0 652 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_746
timestamp 1607101874
transform 1 0 652 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_373
timestamp 1607101874
transform 1 0 804 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_108
timestamp 1607101874
transform 1 0 748 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1607101874
transform -1 0 812 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_193
timestamp 1607101874
transform 1 0 820 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_1_0
timestamp 1607101874
transform 1 0 852 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1607101874
transform 1 0 860 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_329
timestamp 1607101874
transform 1 0 868 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1302
timestamp 1607101874
transform 1 0 812 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_1_0
timestamp 1607101874
transform -1 0 852 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1607101874
transform -1 0 860 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_1303
timestamp 1607101874
transform -1 0 892 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_569
timestamp 1607101874
transform 1 0 892 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_663
timestamp 1607101874
transform 1 0 964 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_551
timestamp 1607101874
transform -1 0 1020 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1607101874
transform 1 0 916 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_742
timestamp 1607101874
transform -1 0 1108 0 -1 1705
box -2 -3 98 103
use BUFX4  BUFX4_455
timestamp 1607101874
transform -1 0 1052 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_479
timestamp 1607101874
transform 1 0 1052 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1607101874
transform -1 0 1116 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_100
timestamp 1607101874
transform -1 0 1140 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_74
timestamp 1607101874
transform 1 0 1116 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_857
timestamp 1607101874
transform -1 0 1180 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_217
timestamp 1607101874
transform 1 0 1180 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_316
timestamp 1607101874
transform 1 0 1212 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_336
timestamp 1607101874
transform 1 0 1140 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_826
timestamp 1607101874
transform 1 0 1156 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_349
timestamp 1607101874
transform 1 0 1308 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_592
timestamp 1607101874
transform 1 0 1252 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_539
timestamp 1607101874
transform -1 0 1300 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_38
timestamp 1607101874
transform 1 0 1300 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_286
timestamp 1607101874
transform -1 0 1372 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_2_0
timestamp 1607101874
transform -1 0 1380 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1607101874
transform -1 0 1388 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_918
timestamp 1607101874
transform -1 0 1420 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_76
timestamp 1607101874
transform 1 0 1332 0 -1 1705
box -2 -3 42 103
use FILL  FILL_16_2_0
timestamp 1607101874
transform 1 0 1372 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1607101874
transform 1 0 1380 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_1212
timestamp 1607101874
transform 1 0 1388 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_236
timestamp 1607101874
transform -1 0 1468 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_963
timestamp 1607101874
transform 1 0 1468 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_53
timestamp 1607101874
transform -1 0 1524 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_591
timestamp 1607101874
transform -1 0 1444 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_119
timestamp 1607101874
transform 1 0 1444 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_67
timestamp 1607101874
transform -1 0 1500 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_94
timestamp 1607101874
transform -1 0 1516 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_836
timestamp 1607101874
transform -1 0 1612 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1294
timestamp 1607101874
transform 1 0 1524 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1295
timestamp 1607101874
transform -1 0 1588 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1607101874
transform 1 0 1588 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_81
timestamp 1607101874
transform -1 0 1660 0 -1 1705
box -2 -3 50 103
use BUFX4  BUFX4_153
timestamp 1607101874
transform -1 0 1716 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1607101874
transform 1 0 1716 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_1092
timestamp 1607101874
transform 1 0 1660 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_920
timestamp 1607101874
transform -1 0 1724 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1305
timestamp 1607101874
transform 1 0 1740 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1304
timestamp 1607101874
transform 1 0 1772 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1607101874
transform 1 0 1804 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_350
timestamp 1607101874
transform 1 0 1724 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_919
timestamp 1607101874
transform 1 0 1740 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1607101874
transform 1 0 1772 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_3_0
timestamp 1607101874
transform -1 0 1908 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1607101874
transform -1 0 1916 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_57
timestamp 1607101874
transform -1 0 1940 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_3_0
timestamp 1607101874
transform 1 0 1868 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1607101874
transform 1 0 1876 0 -1 1705
box -2 -3 10 103
use INVX1  INVX1_414
timestamp 1607101874
transform 1 0 1884 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_289
timestamp 1607101874
transform -1 0 1948 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_58
timestamp 1607101874
transform 1 0 1940 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_769
timestamp 1607101874
transform 1 0 1964 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_770
timestamp 1607101874
transform 1 0 1996 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_497
timestamp 1607101874
transform -1 0 1972 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1093
timestamp 1607101874
transform 1 0 1972 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_467
timestamp 1607101874
transform -1 0 2036 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_426
timestamp 1607101874
transform 1 0 2028 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_852
timestamp 1607101874
transform 1 0 2052 0 1 1505
box -2 -3 98 103
use INVX4  INVX4_5
timestamp 1607101874
transform 1 0 2036 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_336
timestamp 1607101874
transform 1 0 2060 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1215
timestamp 1607101874
transform -1 0 2124 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_96
timestamp 1607101874
transform 1 0 2124 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_83
timestamp 1607101874
transform 1 0 2148 0 1 1505
box -2 -3 50 103
use BUFX4  BUFX4_382
timestamp 1607101874
transform 1 0 2196 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_838
timestamp 1607101874
transform 1 0 2140 0 -1 1705
box -2 -3 98 103
use BUFX4  BUFX4_249
timestamp 1607101874
transform -1 0 2260 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_274
timestamp 1607101874
transform 1 0 2260 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1607101874
transform 1 0 2292 0 1 1505
box -2 -3 98 103
use BUFX4  BUFX4_250
timestamp 1607101874
transform -1 0 2268 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_263
timestamp 1607101874
transform 1 0 2268 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_233
timestamp 1607101874
transform 1 0 2300 0 -1 1705
box -2 -3 34 103
use FILL  FILL_15_4_0
timestamp 1607101874
transform 1 0 2388 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_1
timestamp 1607101874
transform 1 0 2396 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_259
timestamp 1607101874
transform 1 0 2404 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_276
timestamp 1607101874
transform 1 0 2332 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_4_0
timestamp 1607101874
transform -1 0 2372 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_1
timestamp 1607101874
transform -1 0 2380 0 -1 1705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_14
timestamp 1607101874
transform -1 0 2452 0 -1 1705
box -2 -3 74 103
use OAI21X1  OAI21X1_347
timestamp 1607101874
transform 1 0 2428 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_346
timestamp 1607101874
transform -1 0 2492 0 1 1505
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1607101874
transform 1 0 2492 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_82
timestamp 1607101874
transform -1 0 2540 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_399
timestamp 1607101874
transform -1 0 2500 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_560
timestamp 1607101874
transform 1 0 2500 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_344
timestamp 1607101874
transform 1 0 2540 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_345
timestamp 1607101874
transform -1 0 2604 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1607101874
transform 1 0 2604 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_326
timestamp 1607101874
transform 1 0 2596 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_876
timestamp 1607101874
transform 1 0 2612 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1607101874
transform 1 0 2700 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_164
timestamp 1607101874
transform 1 0 2644 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_258
timestamp 1607101874
transform -1 0 2700 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1607101874
transform 1 0 2700 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_793
timestamp 1607101874
transform 1 0 2796 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_454
timestamp 1607101874
transform 1 0 2828 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_453
timestamp 1607101874
transform 1 0 2796 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_347
timestamp 1607101874
transform -1 0 2852 0 -1 1705
box -2 -3 34 103
use INVX8  INVX8_27
timestamp 1607101874
transform 1 0 2852 0 1 1505
box -2 -3 42 103
use FILL  FILL_15_5_0
timestamp 1607101874
transform 1 0 2892 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_1
timestamp 1607101874
transform 1 0 2900 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_878
timestamp 1607101874
transform 1 0 2908 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_29
timestamp 1607101874
transform 1 0 2852 0 -1 1705
box -2 -3 42 103
use FILL  FILL_16_5_0
timestamp 1607101874
transform -1 0 2900 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_5_1
timestamp 1607101874
transform -1 0 2908 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_875
timestamp 1607101874
transform -1 0 2940 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_197
timestamp 1607101874
transform 1 0 2940 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_293
timestamp 1607101874
transform -1 0 2996 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_385
timestamp 1607101874
transform -1 0 3028 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_339
timestamp 1607101874
transform -1 0 3044 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1607101874
transform -1 0 3036 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_362
timestamp 1607101874
transform 1 0 3044 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_363
timestamp 1607101874
transform -1 0 3108 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1607101874
transform -1 0 3204 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_167
timestamp 1607101874
transform 1 0 3036 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_262
timestamp 1607101874
transform 1 0 3068 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_263
timestamp 1607101874
transform 1 0 3092 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_877
timestamp 1607101874
transform -1 0 3148 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_443
timestamp 1607101874
transform 1 0 3204 0 1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_77
timestamp 1607101874
transform 1 0 3220 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_795
timestamp 1607101874
transform 1 0 3148 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_245
timestamp 1607101874
transform 1 0 3180 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_502
timestamp 1607101874
transform -1 0 3236 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_170
timestamp 1607101874
transform 1 0 3252 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_266
timestamp 1607101874
transform -1 0 3308 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_277
timestamp 1607101874
transform 1 0 3308 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_643
timestamp 1607101874
transform 1 0 3324 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1607101874
transform -1 0 3332 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_272
timestamp 1607101874
transform 1 0 3332 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_200
timestamp 1607101874
transform 1 0 3356 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_6_0
timestamp 1607101874
transform 1 0 3380 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_6_1
timestamp 1607101874
transform 1 0 3388 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1607101874
transform 1 0 3396 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_175
timestamp 1607101874
transform -1 0 3388 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1226
timestamp 1607101874
transform -1 0 3420 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_6_0
timestamp 1607101874
transform 1 0 3420 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_1
timestamp 1607101874
transform 1 0 3428 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_15
timestamp 1607101874
transform 1 0 3436 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_1223
timestamp 1607101874
transform 1 0 3492 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_191
timestamp 1607101874
transform -1 0 3556 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1607101874
transform -1 0 3500 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_613
timestamp 1607101874
transform -1 0 3596 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_601
timestamp 1607101874
transform 1 0 3556 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_82
timestamp 1607101874
transform 1 0 3580 0 1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_1222
timestamp 1607101874
transform -1 0 3652 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_347
timestamp 1607101874
transform -1 0 3620 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_348
timestamp 1607101874
transform 1 0 3620 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_794
timestamp 1607101874
transform -1 0 3684 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_737
timestamp 1607101874
transform 1 0 3684 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_625
timestamp 1607101874
transform -1 0 3740 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_564
timestamp 1607101874
transform -1 0 3836 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_402
timestamp 1607101874
transform 1 0 3652 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_327
timestamp 1607101874
transform -1 0 3716 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_597
timestamp 1607101874
transform 1 0 3716 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_253
timestamp 1607101874
transform 1 0 3836 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_6
timestamp 1607101874
transform 1 0 3812 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_3
timestamp 1607101874
transform -1 0 3876 0 -1 1705
box -2 -3 50 103
use BUFX4  BUFX4_333
timestamp 1607101874
transform -1 0 3916 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_7_0
timestamp 1607101874
transform 1 0 3916 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_7_1
timestamp 1607101874
transform 1 0 3924 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1607101874
transform 1 0 3932 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_7_0
timestamp 1607101874
transform 1 0 3876 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_7_1
timestamp 1607101874
transform 1 0 3884 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1607101874
transform 1 0 3892 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_161
timestamp 1607101874
transform 1 0 4028 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_91
timestamp 1607101874
transform 1 0 3988 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_373
timestamp 1607101874
transform -1 0 4044 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_148
timestamp 1607101874
transform -1 0 4092 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_19
timestamp 1607101874
transform -1 0 4116 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_491
timestamp 1607101874
transform 1 0 4116 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_883
timestamp 1607101874
transform 1 0 4140 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1607101874
transform 1 0 4044 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_92
timestamp 1607101874
transform 1 0 4140 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_987
timestamp 1607101874
transform -1 0 4204 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1607101874
transform 1 0 4204 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_24
timestamp 1607101874
transform -1 0 4252 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_374
timestamp 1607101874
transform -1 0 4196 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_375
timestamp 1607101874
transform 1 0 4196 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_451
timestamp 1607101874
transform 1 0 4228 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_456
timestamp 1607101874
transform -1 0 4276 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_30
timestamp 1607101874
transform 1 0 4276 0 1 1505
box -2 -3 42 103
use MUX2X1  MUX2X1_187
timestamp 1607101874
transform 1 0 4316 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_191
timestamp 1607101874
transform 1 0 4260 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_283
timestamp 1607101874
transform -1 0 4308 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_186
timestamp 1607101874
transform -1 0 4340 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1607101874
transform -1 0 4436 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_321
timestamp 1607101874
transform 1 0 4364 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_399
timestamp 1607101874
transform -1 0 4420 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_8_0
timestamp 1607101874
transform -1 0 4428 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_8_1
timestamp 1607101874
transform -1 0 4436 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_400
timestamp 1607101874
transform -1 0 4468 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_8_0
timestamp 1607101874
transform -1 0 4444 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_8_1
timestamp 1607101874
transform -1 0 4452 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_1055
timestamp 1607101874
transform -1 0 4500 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_374
timestamp 1607101874
transform 1 0 4500 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_625
timestamp 1607101874
transform 1 0 4524 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1052
timestamp 1607101874
transform -1 0 4484 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_9
timestamp 1607101874
transform 1 0 4484 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_12
timestamp 1607101874
transform -1 0 4548 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_607
timestamp 1607101874
transform -1 0 4644 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_272
timestamp 1607101874
transform -1 0 4572 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1054
timestamp 1607101874
transform -1 0 4604 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_453
timestamp 1607101874
transform 1 0 4604 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_882
timestamp 1607101874
transform -1 0 4668 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_509
timestamp 1607101874
transform -1 0 4668 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_149
timestamp 1607101874
transform 1 0 4668 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_623
timestamp 1607101874
transform -1 0 4796 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_510
timestamp 1607101874
transform 1 0 4668 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_360
timestamp 1607101874
transform -1 0 4724 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_88
timestamp 1607101874
transform 1 0 4724 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_370
timestamp 1607101874
transform -1 0 4780 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1607101874
transform 1 0 4796 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_10
timestamp 1607101874
transform -1 0 4860 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1607101874
transform -1 0 4876 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_30
timestamp 1607101874
transform -1 0 4884 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_985
timestamp 1607101874
transform -1 0 4916 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_9_0
timestamp 1607101874
transform -1 0 4924 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_9_1
timestamp 1607101874
transform -1 0 4932 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_645
timestamp 1607101874
transform -1 0 5028 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1050
timestamp 1607101874
transform -1 0 4908 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_9_0
timestamp 1607101874
transform 1 0 4908 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_9_1
timestamp 1607101874
transform 1 0 4916 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1607101874
transform 1 0 4924 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_278
timestamp 1607101874
transform -1 0 5044 0 1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_160
timestamp 1607101874
transform 1 0 5044 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_380
timestamp 1607101874
transform 1 0 5020 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_381
timestamp 1607101874
transform -1 0 5084 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1607101874
transform -1 0 5188 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1607101874
transform -1 0 5180 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_158
timestamp 1607101874
transform -1 0 5204 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_640
timestamp 1607101874
transform -1 0 5300 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_142
timestamp 1607101874
transform 1 0 5180 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_175
timestamp 1607101874
transform -1 0 5244 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_155
timestamp 1607101874
transform -1 0 5260 0 -1 1705
box -2 -3 18 103
use FILL  FILL_16_1
timestamp 1607101874
transform 1 0 5300 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_111
timestamp 1607101874
transform -1 0 5284 0 -1 1705
box -2 -3 26 103
use FILL  FILL_17_1
timestamp 1607101874
transform -1 0 5292 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_2
timestamp 1607101874
transform -1 0 5300 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_3
timestamp 1607101874
transform -1 0 5308 0 -1 1705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_75
timestamp 1607101874
transform 1 0 4 0 1 1705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_23
timestamp 1607101874
transform 1 0 76 0 1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_546
timestamp 1607101874
transform 1 0 148 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_734
timestamp 1607101874
transform 1 0 244 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_0_0
timestamp 1607101874
transform 1 0 340 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1607101874
transform 1 0 348 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_289
timestamp 1607101874
transform 1 0 356 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_81
timestamp 1607101874
transform -1 0 396 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_80
timestamp 1607101874
transform 1 0 396 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_705
timestamp 1607101874
transform 1 0 420 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_223
timestamp 1607101874
transform -1 0 476 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_743
timestamp 1607101874
transform -1 0 572 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_102
timestamp 1607101874
transform 1 0 572 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_738
timestamp 1607101874
transform 1 0 604 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_60
timestamp 1607101874
transform 1 0 700 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_1178
timestamp 1607101874
transform 1 0 716 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_126
timestamp 1607101874
transform -1 0 772 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_72
timestamp 1607101874
transform -1 0 804 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_1_0
timestamp 1607101874
transform 1 0 804 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1607101874
transform 1 0 812 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_831
timestamp 1607101874
transform 1 0 820 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1180
timestamp 1607101874
transform -1 0 948 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1179
timestamp 1607101874
transform -1 0 980 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_816
timestamp 1607101874
transform 1 0 980 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_147
timestamp 1607101874
transform 1 0 1076 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_146
timestamp 1607101874
transform -1 0 1140 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_183
timestamp 1607101874
transform 1 0 1140 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_71
timestamp 1607101874
transform 1 0 1172 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_124
timestamp 1607101874
transform -1 0 1228 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_818
timestamp 1607101874
transform 1 0 1228 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_151
timestamp 1607101874
transform 1 0 1324 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_2_0
timestamp 1607101874
transform -1 0 1364 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1607101874
transform -1 0 1372 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_150
timestamp 1607101874
transform -1 0 1404 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_394
timestamp 1607101874
transform 1 0 1404 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_814
timestamp 1607101874
transform -1 0 1524 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_681
timestamp 1607101874
transform -1 0 1556 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_286
timestamp 1607101874
transform -1 0 1580 0 1 1705
box -2 -3 26 103
use INVX8  INVX8_19
timestamp 1607101874
transform -1 0 1620 0 1 1705
box -2 -3 42 103
use INVX8  INVX8_16
timestamp 1607101874
transform -1 0 1660 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_477
timestamp 1607101874
transform 1 0 1660 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1607101874
transform -1 0 1716 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_680
timestamp 1607101874
transform -1 0 1748 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_36
timestamp 1607101874
transform -1 0 1772 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1297
timestamp 1607101874
transform 1 0 1772 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1607101874
transform 1 0 1804 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_3_0
timestamp 1607101874
transform -1 0 1908 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1607101874
transform -1 0 1916 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_1296
timestamp 1607101874
transform -1 0 1948 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_466
timestamp 1607101874
transform -1 0 1980 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1607101874
transform 1 0 1980 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1094
timestamp 1607101874
transform 1 0 2012 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1607101874
transform 1 0 2044 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_763
timestamp 1607101874
transform -1 0 2108 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_49
timestamp 1607101874
transform 1 0 2108 0 1 1705
box -2 -3 50 103
use NOR2X1  NOR2X1_570
timestamp 1607101874
transform -1 0 2180 0 1 1705
box -2 -3 26 103
use BUFX4  BUFX4_39
timestamp 1607101874
transform -1 0 2212 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_8
timestamp 1607101874
transform 1 0 2212 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_252
timestamp 1607101874
transform 1 0 2252 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1607101874
transform -1 0 2316 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_232
timestamp 1607101874
transform -1 0 2348 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_255
timestamp 1607101874
transform 1 0 2348 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_4_0
timestamp 1607101874
transform 1 0 2380 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1607101874
transform 1 0 2388 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_434
timestamp 1607101874
transform 1 0 2396 0 1 1705
box -2 -3 98 103
use OAI22X1  OAI22X1_69
timestamp 1607101874
transform -1 0 2532 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_34
timestamp 1607101874
transform 1 0 2532 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1607101874
transform -1 0 2596 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1607101874
transform 1 0 2596 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_359
timestamp 1607101874
transform 1 0 2620 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1607101874
transform 1 0 2652 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_358
timestamp 1607101874
transform -1 0 2780 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1607101874
transform 1 0 2780 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1225
timestamp 1607101874
transform 1 0 2804 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_83
timestamp 1607101874
transform 1 0 2836 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_5_0
timestamp 1607101874
transform 1 0 2860 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1607101874
transform 1 0 2868 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_589
timestamp 1607101874
transform 1 0 2876 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1566
timestamp 1607101874
transform 1 0 2972 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1565
timestamp 1607101874
transform -1 0 3036 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_879
timestamp 1607101874
transform -1 0 3068 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_384
timestamp 1607101874
transform 1 0 3068 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_386
timestamp 1607101874
transform 1 0 3100 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_136
timestamp 1607101874
transform 1 0 3132 0 1 1705
box -2 -3 50 103
use INVX1  INVX1_149
timestamp 1607101874
transform -1 0 3196 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1607101874
transform -1 0 3292 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_8
timestamp 1607101874
transform 1 0 3292 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1607101874
transform -1 0 3348 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_621
timestamp 1607101874
transform 1 0 3348 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_6_0
timestamp 1607101874
transform 1 0 3444 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1607101874
transform 1 0 3452 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_977
timestamp 1607101874
transform 1 0 3460 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_978
timestamp 1607101874
transform 1 0 3492 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_489
timestamp 1607101874
transform 1 0 3524 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_11
timestamp 1607101874
transform 1 0 3548 0 1 1705
box -2 -3 50 103
use INVX1  INVX1_16
timestamp 1607101874
transform -1 0 3612 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_609
timestamp 1607101874
transform -1 0 3708 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1607101874
transform 1 0 3708 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_172
timestamp 1607101874
transform 1 0 3804 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_159
timestamp 1607101874
transform -1 0 3868 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_881
timestamp 1607101874
transform 1 0 3868 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_507
timestamp 1607101874
transform 1 0 3900 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_7_0
timestamp 1607101874
transform -1 0 3932 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_7_1
timestamp 1607101874
transform -1 0 3940 0 1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_225
timestamp 1607101874
transform -1 0 3988 0 1 1705
box -2 -3 50 103
use BUFX4  BUFX4_427
timestamp 1607101874
transform 1 0 3988 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1607101874
transform 1 0 4020 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_168
timestamp 1607101874
transform 1 0 4116 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_155
timestamp 1607101874
transform -1 0 4180 0 1 1705
box -2 -3 50 103
use NOR2X1  NOR2X1_451
timestamp 1607101874
transform -1 0 4204 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1051
timestamp 1607101874
transform 1 0 4204 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_264
timestamp 1607101874
transform 1 0 4236 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_880
timestamp 1607101874
transform -1 0 4292 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_867
timestamp 1607101874
transform 1 0 4292 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_27
timestamp 1607101874
transform -1 0 4364 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_868
timestamp 1607101874
transform -1 0 4396 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_8_0
timestamp 1607101874
transform 1 0 4396 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_8_1
timestamp 1607101874
transform 1 0 4404 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1607101874
transform 1 0 4412 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_151
timestamp 1607101874
transform 1 0 4508 0 1 1705
box -2 -3 50 103
use INVX1  INVX1_164
timestamp 1607101874
transform -1 0 4572 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1607101874
transform -1 0 4668 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_638
timestamp 1607101874
transform 1 0 4668 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_24
timestamp 1607101874
transform -1 0 4732 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1607101874
transform -1 0 4828 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_86
timestamp 1607101874
transform 1 0 4828 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_368
timestamp 1607101874
transform -1 0 4884 0 1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_81
timestamp 1607101874
transform -1 0 4956 0 1 1705
box -2 -3 74 103
use FILL  FILL_17_9_0
timestamp 1607101874
transform -1 0 4964 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_9_1
timestamp 1607101874
transform -1 0 4972 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_201
timestamp 1607101874
transform -1 0 4996 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_282
timestamp 1607101874
transform 1 0 4996 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_185
timestamp 1607101874
transform -1 0 5052 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_280
timestamp 1607101874
transform -1 0 5068 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_144
timestamp 1607101874
transform 1 0 5068 0 1 1705
box -2 -3 50 103
use INVX1  INVX1_157
timestamp 1607101874
transform -1 0 5132 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1607101874
transform -1 0 5228 0 1 1705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_98
timestamp 1607101874
transform -1 0 5300 0 1 1705
box -2 -3 74 103
use FILL  FILL_18_1
timestamp 1607101874
transform 1 0 5300 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_824
timestamp 1607101874
transform -1 0 100 0 -1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_122
timestamp 1607101874
transform 1 0 100 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_69
timestamp 1607101874
transform -1 0 156 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_310
timestamp 1607101874
transform 1 0 156 0 -1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_491
timestamp 1607101874
transform 1 0 252 0 -1 1905
box -2 -3 34 103
use AND2X2  AND2X2_53
timestamp 1607101874
transform 1 0 284 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_249
timestamp 1607101874
transform 1 0 316 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_0_0
timestamp 1607101874
transform -1 0 340 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1607101874
transform -1 0 348 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_319
timestamp 1607101874
transform -1 0 396 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_552
timestamp 1607101874
transform -1 0 492 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_395
timestamp 1607101874
transform 1 0 492 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_788
timestamp 1607101874
transform 1 0 540 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_789
timestamp 1607101874
transform 1 0 572 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_270
timestamp 1607101874
transform 1 0 604 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_50
timestamp 1607101874
transform -1 0 684 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_590
timestamp 1607101874
transform 1 0 684 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_494
timestamp 1607101874
transform 1 0 716 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1343
timestamp 1607101874
transform 1 0 748 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1342
timestamp 1607101874
transform -1 0 812 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_205
timestamp 1607101874
transform -1 0 860 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_1_0
timestamp 1607101874
transform -1 0 868 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1607101874
transform -1 0 876 0 -1 1905
box -2 -3 10 103
use BUFX4  BUFX4_187
timestamp 1607101874
transform -1 0 908 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_840
timestamp 1607101874
transform 1 0 908 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_98
timestamp 1607101874
transform 1 0 1004 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_85
timestamp 1607101874
transform -1 0 1068 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_854
timestamp 1607101874
transform 1 0 1068 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_376
timestamp 1607101874
transform 1 0 1100 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_859
timestamp 1607101874
transform -1 0 1164 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_822
timestamp 1607101874
transform 1 0 1164 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_159
timestamp 1607101874
transform 1 0 1260 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_158
timestamp 1607101874
transform -1 0 1324 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1213
timestamp 1607101874
transform 1 0 1324 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_2_0
timestamp 1607101874
transform -1 0 1364 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1607101874
transform -1 0 1372 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_856
timestamp 1607101874
transform -1 0 1404 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_855
timestamp 1607101874
transform -1 0 1436 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_327
timestamp 1607101874
transform 1 0 1436 0 -1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_423
timestamp 1607101874
transform -1 0 1556 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_664
timestamp 1607101874
transform -1 0 1580 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_552
timestamp 1607101874
transform -1 0 1612 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_311
timestamp 1607101874
transform -1 0 1708 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_55
timestamp 1607101874
transform -1 0 1732 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_84
timestamp 1607101874
transform 1 0 1732 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_97
timestamp 1607101874
transform -1 0 1796 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_839
timestamp 1607101874
transform -1 0 1892 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_3_0
timestamp 1607101874
transform 1 0 1892 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1607101874
transform 1 0 1900 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_744
timestamp 1607101874
transform 1 0 1908 0 -1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_272
timestamp 1607101874
transform 1 0 2004 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_332
timestamp 1607101874
transform -1 0 2060 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_59
timestamp 1607101874
transform -1 0 2076 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_736
timestamp 1607101874
transform -1 0 2172 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_830
timestamp 1607101874
transform 1 0 2172 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_362
timestamp 1607101874
transform -1 0 2236 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_122
timestamp 1607101874
transform 1 0 2236 0 -1 1905
box -2 -3 34 103
use XOR2X1  XOR2X1_5
timestamp 1607101874
transform -1 0 2324 0 -1 1905
box -2 -3 58 103
use INVX2  INVX2_4
timestamp 1607101874
transform -1 0 2340 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_547
timestamp 1607101874
transform 1 0 2340 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_4_0
timestamp 1607101874
transform -1 0 2380 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1607101874
transform -1 0 2388 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_548
timestamp 1607101874
transform -1 0 2420 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1607101874
transform 1 0 2420 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_5
timestamp 1607101874
transform -1 0 2460 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_11
timestamp 1607101874
transform 1 0 2460 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_13
timestamp 1607101874
transform 1 0 2484 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_9
timestamp 1607101874
transform -1 0 2524 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1607101874
transform -1 0 2556 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1607101874
transform -1 0 2580 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_4
timestamp 1607101874
transform -1 0 2612 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_9
timestamp 1607101874
transform 1 0 2612 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_23
timestamp 1607101874
transform 1 0 2636 0 -1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_2
timestamp 1607101874
transform -1 0 2684 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1607101874
transform -1 0 2716 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1607101874
transform 1 0 2716 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_353
timestamp 1607101874
transform 1 0 2812 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_352
timestamp 1607101874
transform -1 0 2876 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_5_0
timestamp 1607101874
transform 1 0 2876 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1607101874
transform 1 0 2884 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1607101874
transform 1 0 2892 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_361
timestamp 1607101874
transform 1 0 2988 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_360
timestamp 1607101874
transform -1 0 3052 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_295
timestamp 1607101874
transform -1 0 3076 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_198
timestamp 1607101874
transform 1 0 3076 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_486
timestamp 1607101874
transform 1 0 3100 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_642
timestamp 1607101874
transform 1 0 3124 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1607101874
transform 1 0 3156 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_193
timestamp 1607101874
transform 1 0 3180 0 -1 1905
box -2 -3 50 103
use AOI21X1  AOI21X1_166
timestamp 1607101874
transform 1 0 3228 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_261
timestamp 1607101874
transform 1 0 3260 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1607101874
transform -1 0 3380 0 -1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_427
timestamp 1607101874
transform 1 0 3380 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_981
timestamp 1607101874
transform 1 0 3428 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_350
timestamp 1607101874
transform -1 0 3492 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_605
timestamp 1607101874
transform 1 0 3492 0 -1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_503
timestamp 1607101874
transform 1 0 3588 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1607101874
transform 1 0 3620 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_7
timestamp 1607101874
transform -1 0 3684 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_979
timestamp 1607101874
transform 1 0 3684 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_78
timestamp 1607101874
transform 1 0 3716 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1607101874
transform 1 0 3748 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_4
timestamp 1607101874
transform -1 0 3804 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_980
timestamp 1607101874
transform -1 0 3836 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_7
timestamp 1607101874
transform 1 0 3836 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1607101874
transform -1 0 3892 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_330
timestamp 1607101874
transform 1 0 3892 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_7_0
timestamp 1607101874
transform 1 0 3908 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_7_1
timestamp 1607101874
transform 1 0 3916 0 -1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_387
timestamp 1607101874
transform 1 0 3924 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_352
timestamp 1607101874
transform 1 0 3956 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_347
timestamp 1607101874
transform 1 0 3988 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_884
timestamp 1607101874
transform -1 0 4052 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_36
timestamp 1607101874
transform 1 0 4052 0 -1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_14
timestamp 1607101874
transform 1 0 4084 0 -1 1905
box -2 -3 66 103
use OAI21X1  OAI21X1_869
timestamp 1607101874
transform -1 0 4180 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_351
timestamp 1607101874
transform -1 0 4212 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_293
timestamp 1607101874
transform -1 0 4244 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_10
timestamp 1607101874
transform 1 0 4244 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_15
timestamp 1607101874
transform -1 0 4308 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_608
timestamp 1607101874
transform -1 0 4404 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_150
timestamp 1607101874
transform 1 0 4404 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_8_0
timestamp 1607101874
transform -1 0 4460 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_8_1
timestamp 1607101874
transform -1 0 4468 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_163
timestamp 1607101874
transform -1 0 4484 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_559
timestamp 1607101874
transform 1 0 4484 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_297
timestamp 1607101874
transform 1 0 4508 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_377
timestamp 1607101874
transform 1 0 4540 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_295
timestamp 1607101874
transform 1 0 4564 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_639
timestamp 1607101874
transform -1 0 4628 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_637
timestamp 1607101874
transform 1 0 4628 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_592
timestamp 1607101874
transform 1 0 4660 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1570
timestamp 1607101874
transform 1 0 4756 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_362
timestamp 1607101874
transform -1 0 4812 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_801
timestamp 1607101874
transform 1 0 4812 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_353
timestamp 1607101874
transform -1 0 4876 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_799
timestamp 1607101874
transform -1 0 4908 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_436
timestamp 1607101874
transform -1 0 4932 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_9_0
timestamp 1607101874
transform 1 0 4932 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_9_1
timestamp 1607101874
transform 1 0 4940 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_646
timestamp 1607101874
transform 1 0 4948 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_636
timestamp 1607101874
transform -1 0 5012 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_296
timestamp 1607101874
transform -1 0 5044 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1607101874
transform 1 0 5044 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_14
timestamp 1607101874
transform -1 0 5108 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_154
timestamp 1607101874
transform 1 0 5108 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_86
timestamp 1607101874
transform -1 0 5172 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_2
timestamp 1607101874
transform 1 0 5172 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_6
timestamp 1607101874
transform 1 0 5220 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_9
timestamp 1607101874
transform -1 0 5284 0 -1 1905
box -2 -3 18 103
use FILL  FILL_19_1
timestamp 1607101874
transform -1 0 5292 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_2
timestamp 1607101874
transform -1 0 5300 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_3
timestamp 1607101874
transform -1 0 5308 0 -1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_17
timestamp 1607101874
transform 1 0 4 0 1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_436
timestamp 1607101874
transform 1 0 76 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_550
timestamp 1607101874
transform -1 0 204 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_438
timestamp 1607101874
transform 1 0 204 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_1170
timestamp 1607101874
transform 1 0 220 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1171
timestamp 1607101874
transform 1 0 252 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1172
timestamp 1607101874
transform -1 0 316 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1607101874
transform 1 0 316 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_0_0
timestamp 1607101874
transform 1 0 348 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1607101874
transform 1 0 356 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_589
timestamp 1607101874
transform 1 0 364 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_177
timestamp 1607101874
transform 1 0 396 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_323
timestamp 1607101874
transform 1 0 420 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_322
timestamp 1607101874
transform -1 0 532 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_318
timestamp 1607101874
transform 1 0 532 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_271
timestamp 1607101874
transform -1 0 660 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_819
timestamp 1607101874
transform 1 0 660 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1351
timestamp 1607101874
transform -1 0 788 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1607101874
transform 1 0 788 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_1_0
timestamp 1607101874
transform 1 0 820 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1607101874
transform 1 0 828 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_512
timestamp 1607101874
transform 1 0 836 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_320
timestamp 1607101874
transform 1 0 932 0 1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_382
timestamp 1607101874
transform -1 0 996 0 1 1905
box -2 -3 50 103
use BUFX4  BUFX4_218
timestamp 1607101874
transform -1 0 1028 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_323
timestamp 1607101874
transform 1 0 1028 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1345
timestamp 1607101874
transform 1 0 1124 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1344
timestamp 1607101874
transform -1 0 1188 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1607101874
transform 1 0 1188 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_820
timestamp 1607101874
transform 1 0 1220 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_154
timestamp 1607101874
transform -1 0 1348 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1607101874
transform 1 0 1348 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1607101874
transform 1 0 1356 0 1 1905
box -2 -3 10 103
use AND2X2  AND2X2_34
timestamp 1607101874
transform 1 0 1364 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_759
timestamp 1607101874
transform 1 0 1396 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1356
timestamp 1607101874
transform 1 0 1428 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_321
timestamp 1607101874
transform -1 0 1556 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1357
timestamp 1607101874
transform -1 0 1588 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_682
timestamp 1607101874
transform 1 0 1588 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_550
timestamp 1607101874
transform 1 0 1620 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_662
timestamp 1607101874
transform -1 0 1676 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_422
timestamp 1607101874
transform -1 0 1700 0 1 1905
box -2 -3 26 103
use OAI22X1  OAI22X1_20
timestamp 1607101874
transform -1 0 1740 0 1 1905
box -2 -3 42 103
use BUFX4  BUFX4_388
timestamp 1607101874
transform 1 0 1740 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_52
timestamp 1607101874
transform -1 0 1796 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_116
timestamp 1607101874
transform 1 0 1796 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_51
timestamp 1607101874
transform 1 0 1820 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1122
timestamp 1607101874
transform 1 0 1844 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_3_0
timestamp 1607101874
transform -1 0 1884 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1607101874
transform -1 0 1892 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_178
timestamp 1607101874
transform -1 0 1916 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_130
timestamp 1607101874
transform 1 0 1916 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_541
timestamp 1607101874
transform -1 0 1964 0 1 1905
box -2 -3 26 103
use OAI22X1  OAI22X1_59
timestamp 1607101874
transform 1 0 1964 0 1 1905
box -2 -3 42 103
use MUX2X1  MUX2X1_222
timestamp 1607101874
transform 1 0 2004 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_1127
timestamp 1607101874
transform 1 0 2052 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_13
timestamp 1607101874
transform 1 0 2084 0 1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_760
timestamp 1607101874
transform 1 0 2124 0 1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_85
timestamp 1607101874
transform -1 0 2228 0 1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_432
timestamp 1607101874
transform -1 0 2324 0 1 1905
box -2 -3 98 103
use BUFX4  BUFX4_226
timestamp 1607101874
transform -1 0 2356 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_247
timestamp 1607101874
transform 1 0 2356 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_4_0
timestamp 1607101874
transform 1 0 2388 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1607101874
transform 1 0 2396 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_227
timestamp 1607101874
transform 1 0 2404 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_254
timestamp 1607101874
transform 1 0 2436 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_235
timestamp 1607101874
transform -1 0 2500 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_26
timestamp 1607101874
transform -1 0 2524 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_14
timestamp 1607101874
transform -1 0 2540 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_10
timestamp 1607101874
transform -1 0 2564 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1607101874
transform -1 0 2588 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1607101874
transform -1 0 2612 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_17
timestamp 1607101874
transform -1 0 2636 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_32
timestamp 1607101874
transform -1 0 2660 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_18
timestamp 1607101874
transform 1 0 2660 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1607101874
transform -1 0 2708 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1607101874
transform 1 0 2708 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_2
timestamp 1607101874
transform -1 0 2748 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1607101874
transform 1 0 2748 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_4
timestamp 1607101874
transform 1 0 2772 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_23
timestamp 1607101874
transform -1 0 2820 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_10
timestamp 1607101874
transform 1 0 2820 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1607101874
transform -1 0 2868 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_15
timestamp 1607101874
transform -1 0 2892 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_5_0
timestamp 1607101874
transform 1 0 2892 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1607101874
transform 1 0 2900 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_1558
timestamp 1607101874
transform 1 0 2908 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_585
timestamp 1607101874
transform 1 0 2940 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1557
timestamp 1607101874
transform 1 0 3036 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_974
timestamp 1607101874
transform -1 0 3100 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_276
timestamp 1607101874
transform 1 0 3100 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_641
timestamp 1607101874
transform 1 0 3116 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_975
timestamp 1607101874
transform 1 0 3148 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_487
timestamp 1607101874
transform -1 0 3204 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_488
timestamp 1607101874
transform -1 0 3228 0 1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_27
timestamp 1607101874
transform 1 0 3228 0 1 1905
box -2 -3 42 103
use BUFX4  BUFX4_175
timestamp 1607101874
transform -1 0 3300 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_617
timestamp 1607101874
transform -1 0 3396 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_25
timestamp 1607101874
transform 1 0 3396 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_6_0
timestamp 1607101874
transform -1 0 3420 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1607101874
transform -1 0 3428 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_976
timestamp 1607101874
transform -1 0 3460 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_19
timestamp 1607101874
transform -1 0 3508 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_885
timestamp 1607101874
transform -1 0 3540 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_169
timestamp 1607101874
transform 1 0 3540 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_146
timestamp 1607101874
transform -1 0 3604 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1607101874
transform 1 0 3604 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_428
timestamp 1607101874
transform -1 0 3668 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_601
timestamp 1607101874
transform -1 0 3764 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_620
timestamp 1607101874
transform 1 0 3764 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_429
timestamp 1607101874
transform -1 0 3892 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_7_0
timestamp 1607101874
transform 1 0 3892 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_7_1
timestamp 1607101874
transform 1 0 3900 0 1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_47
timestamp 1607101874
transform 1 0 3908 0 1 1905
box -2 -3 74 103
use OAI21X1  OAI21X1_800
timestamp 1607101874
transform -1 0 4012 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1607101874
transform 1 0 4012 0 1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_18
timestamp 1607101874
transform -1 0 4076 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_993
timestamp 1607101874
transform -1 0 4108 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_616
timestamp 1607101874
transform -1 0 4204 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_593
timestamp 1607101874
transform -1 0 4300 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_363
timestamp 1607101874
transform 1 0 4300 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1571
timestamp 1607101874
transform -1 0 4356 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_209
timestamp 1607101874
transform 1 0 4356 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_8_0
timestamp 1607101874
transform 1 0 4388 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_8_1
timestamp 1607101874
transform 1 0 4396 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1607101874
transform 1 0 4404 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1607101874
transform -1 0 4596 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_90
timestamp 1607101874
transform 1 0 4596 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_372
timestamp 1607101874
transform -1 0 4652 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_344
timestamp 1607101874
transform -1 0 4668 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_360
timestamp 1607101874
transform -1 0 4764 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_803
timestamp 1607101874
transform -1 0 4796 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_802
timestamp 1607101874
transform -1 0 4828 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_202
timestamp 1607101874
transform -1 0 4852 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_647
timestamp 1607101874
transform -1 0 4884 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_279
timestamp 1607101874
transform -1 0 4900 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_9_0
timestamp 1607101874
transform -1 0 4908 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_9_1
timestamp 1607101874
transform -1 0 4916 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_612
timestamp 1607101874
transform -1 0 5012 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_3
timestamp 1607101874
transform 1 0 5012 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1607101874
transform -1 0 5068 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_600
timestamp 1607101874
transform -1 0 5164 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_604
timestamp 1607101874
transform -1 0 5260 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_543
timestamp 1607101874
transform -1 0 5292 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1607101874
transform 1 0 5292 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1607101874
transform 1 0 5300 0 1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_42
timestamp 1607101874
transform 1 0 4 0 -1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_554
timestamp 1607101874
transform 1 0 76 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_439
timestamp 1607101874
transform 1 0 172 0 -1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_397
timestamp 1607101874
transform -1 0 236 0 -1 2105
box -2 -3 50 103
use AOI21X1  AOI21X1_70
timestamp 1607101874
transform 1 0 236 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_123
timestamp 1607101874
transform -1 0 292 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_549
timestamp 1607101874
transform -1 0 324 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_304
timestamp 1607101874
transform 1 0 324 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_0_0
timestamp 1607101874
transform -1 0 356 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1607101874
transform -1 0 364 0 -1 2105
box -2 -3 10 103
use INVX2  INVX2_1
timestamp 1607101874
transform -1 0 380 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_3
timestamp 1607101874
transform 1 0 380 0 -1 2105
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1607101874
transform -1 0 428 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_435
timestamp 1607101874
transform -1 0 524 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_52
timestamp 1607101874
transform -1 0 548 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1607101874
transform 1 0 548 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_13
timestamp 1607101874
transform 1 0 564 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_37
timestamp 1607101874
transform -1 0 612 0 -1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_9
timestamp 1607101874
transform -1 0 668 0 -1 2105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_821
timestamp 1607101874
transform -1 0 764 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_1350
timestamp 1607101874
transform -1 0 796 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_156
timestamp 1607101874
transform -1 0 828 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1607101874
transform -1 0 860 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_1_0
timestamp 1607101874
transform 1 0 860 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1607101874
transform 1 0 868 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_152
timestamp 1607101874
transform 1 0 876 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_8
timestamp 1607101874
transform 1 0 908 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_360
timestamp 1607101874
transform -1 0 948 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_428
timestamp 1607101874
transform 1 0 948 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_313
timestamp 1607101874
transform 1 0 980 0 -1 2105
box -2 -3 98 103
use AND2X2  AND2X2_20
timestamp 1607101874
transform 1 0 1076 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_553
timestamp 1607101874
transform 1 0 1108 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_665
timestamp 1607101874
transform -1 0 1164 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_678
timestamp 1607101874
transform 1 0 1164 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_10
timestamp 1607101874
transform 1 0 1196 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_783
timestamp 1607101874
transform 1 0 1212 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_214
timestamp 1607101874
transform 1 0 1244 0 -1 2105
box -2 -3 50 103
use OAI22X1  OAI22X1_13
timestamp 1607101874
transform 1 0 1292 0 -1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_540
timestamp 1607101874
transform 1 0 1332 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_2_0
timestamp 1607101874
transform 1 0 1356 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1607101874
transform 1 0 1364 0 -1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_282
timestamp 1607101874
transform 1 0 1372 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_677
timestamp 1607101874
transform -1 0 1436 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_329
timestamp 1607101874
transform -1 0 1460 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1119
timestamp 1607101874
transform 1 0 1460 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_56
timestamp 1607101874
transform 1 0 1492 0 -1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_1118
timestamp 1607101874
transform -1 0 1564 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_393
timestamp 1607101874
transform -1 0 1588 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_395
timestamp 1607101874
transform 1 0 1588 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_3
timestamp 1607101874
transform 1 0 1612 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_51
timestamp 1607101874
transform 1 0 1628 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_115
timestamp 1607101874
transform 1 0 1652 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_11
timestamp 1607101874
transform 1 0 1676 0 -1 2105
box -2 -3 18 103
use BUFX4  BUFX4_184
timestamp 1607101874
transform 1 0 1692 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_325
timestamp 1607101874
transform -1 0 1820 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_1348
timestamp 1607101874
transform -1 0 1852 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1349
timestamp 1607101874
transform -1 0 1884 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 2105
box -2 -3 10 103
use INVX2  INVX2_9
timestamp 1607101874
transform 1 0 1900 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_144
timestamp 1607101874
transform 1 0 1916 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1607101874
transform -1 0 1980 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_815
timestamp 1607101874
transform -1 0 2076 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_1352
timestamp 1607101874
transform 1 0 2076 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1353
timestamp 1607101874
transform 1 0 2108 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_319
timestamp 1607101874
transform 1 0 2140 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_325
timestamp 1607101874
transform -1 0 2268 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1607101874
transform 1 0 2268 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_236
timestamp 1607101874
transform -1 0 2332 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_220
timestamp 1607101874
transform -1 0 2364 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_283
timestamp 1607101874
transform 1 0 2364 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_4_0
timestamp 1607101874
transform 1 0 2396 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1607101874
transform 1 0 2404 0 -1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_21
timestamp 1607101874
transform 1 0 2412 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_219
timestamp 1607101874
transform 1 0 2436 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1607101874
transform 1 0 2468 0 -1 2105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_11
timestamp 1607101874
transform -1 0 2564 0 -1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_433
timestamp 1607101874
transform -1 0 2660 0 -1 2105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_8
timestamp 1607101874
transform -1 0 2716 0 -1 2105
box -2 -3 58 103
use NOR2X1  NOR2X1_256
timestamp 1607101874
transform -1 0 2740 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_53
timestamp 1607101874
transform -1 0 2764 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1607101874
transform 1 0 2764 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_271
timestamp 1607101874
transform 1 0 2860 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_5_0
timestamp 1607101874
transform -1 0 2892 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1607101874
transform -1 0 2900 0 -1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_174
timestamp 1607101874
transform -1 0 2932 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_640
timestamp 1607101874
transform -1 0 2964 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_151
timestamp 1607101874
transform -1 0 2980 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1607101874
transform -1 0 3076 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_152
timestamp 1607101874
transform 1 0 3076 0 -1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_138
timestamp 1607101874
transform -1 0 3140 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_139
timestamp 1607101874
transform 1 0 3140 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_973
timestamp 1607101874
transform 1 0 3188 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_229
timestamp 1607101874
transform 1 0 3220 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_278
timestamp 1607101874
transform 1 0 3252 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_192
timestamp 1607101874
transform 1 0 3284 0 -1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_378
timestamp 1607101874
transform 1 0 3332 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_645
timestamp 1607101874
transform 1 0 3356 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_426
timestamp 1607101874
transform -1 0 3420 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_6_0
timestamp 1607101874
transform 1 0 3420 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1607101874
transform 1 0 3428 0 -1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_410
timestamp 1607101874
transform 1 0 3436 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_391
timestamp 1607101874
transform -1 0 3500 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_581
timestamp 1607101874
transform -1 0 3596 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_557
timestamp 1607101874
transform -1 0 3620 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_746
timestamp 1607101874
transform 1 0 3620 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_507
timestamp 1607101874
transform -1 0 3684 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1607101874
transform 1 0 3684 0 -1 2105
box -2 -3 42 103
use OAI22X1  OAI22X1_46
timestamp 1607101874
transform -1 0 3764 0 -1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_300
timestamp 1607101874
transform 1 0 3764 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_246
timestamp 1607101874
transform -1 0 3812 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_805
timestamp 1607101874
transform -1 0 3844 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_804
timestamp 1607101874
transform -1 0 3876 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_71
timestamp 1607101874
transform -1 0 3908 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_7_0
timestamp 1607101874
transform 1 0 3908 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_7_1
timestamp 1607101874
transform 1 0 3916 0 -1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_73
timestamp 1607101874
transform 1 0 3924 0 -1 2105
box -2 -3 74 103
use BUFX4  BUFX4_69
timestamp 1607101874
transform 1 0 3996 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_299
timestamp 1607101874
transform 1 0 4028 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_298
timestamp 1607101874
transform -1 0 4092 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_197
timestamp 1607101874
transform -1 0 4140 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_651
timestamp 1607101874
transform 1 0 4140 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_206
timestamp 1607101874
transform -1 0 4196 0 -1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1607101874
transform -1 0 4236 0 -1 2105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1607101874
transform -1 0 4332 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_429
timestamp 1607101874
transform -1 0 4364 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_430
timestamp 1607101874
transform -1 0 4396 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_650
timestamp 1607101874
transform 1 0 4396 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_8_0
timestamp 1607101874
transform -1 0 4436 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_8_1
timestamp 1607101874
transform -1 0 4444 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_205
timestamp 1607101874
transform -1 0 4468 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_633
timestamp 1607101874
transform 1 0 4468 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_189
timestamp 1607101874
transform 1 0 4500 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_630
timestamp 1607101874
transform 1 0 4548 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1607101874
transform -1 0 4604 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_59
timestamp 1607101874
transform 1 0 4604 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_60
timestamp 1607101874
transform -1 0 4668 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_423
timestamp 1607101874
transform 1 0 4668 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_307
timestamp 1607101874
transform -1 0 4748 0 -1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_683
timestamp 1607101874
transform -1 0 4844 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1607101874
transform -1 0 4940 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_9_0
timestamp 1607101874
transform 1 0 4940 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_9_1
timestamp 1607101874
transform 1 0 4948 0 -1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_194
timestamp 1607101874
transform 1 0 4956 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_195
timestamp 1607101874
transform 1 0 5004 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_648
timestamp 1607101874
transform 1 0 5052 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_635
timestamp 1607101874
transform -1 0 5116 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1607101874
transform -1 0 5212 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_59
timestamp 1607101874
transform -1 0 5244 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_158
timestamp 1607101874
transform 1 0 5244 0 -1 2105
box -2 -3 50 103
use FILL  FILL_21_1
timestamp 1607101874
transform -1 0 5300 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_2
timestamp 1607101874
transform -1 0 5308 0 -1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_64
timestamp 1607101874
transform 1 0 4 0 1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1042
timestamp 1607101874
transform 1 0 76 0 1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_155
timestamp 1607101874
transform 1 0 172 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_244
timestamp 1607101874
transform 1 0 204 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_825
timestamp 1607101874
transform 1 0 228 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_0_0
timestamp 1607101874
transform -1 0 332 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1607101874
transform -1 0 340 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_1340
timestamp 1607101874
transform -1 0 372 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_248
timestamp 1607101874
transform -1 0 388 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_326
timestamp 1607101874
transform -1 0 484 0 1 2105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_36
timestamp 1607101874
transform 1 0 484 0 1 2105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_79
timestamp 1607101874
transform 1 0 556 0 1 2105
box -2 -3 74 103
use INVX8  INVX8_26
timestamp 1607101874
transform -1 0 668 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_1007
timestamp 1607101874
transform -1 0 700 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_395
timestamp 1607101874
transform -1 0 716 0 1 2105
box -2 -3 18 103
use INVX8  INVX8_9
timestamp 1607101874
transform -1 0 756 0 1 2105
box -2 -3 42 103
use INVX2  INVX2_7
timestamp 1607101874
transform 1 0 756 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_303
timestamp 1607101874
transform -1 0 796 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_148
timestamp 1607101874
transform 1 0 796 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1607101874
transform -1 0 860 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_1_0
timestamp 1607101874
transform -1 0 868 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1607101874
transform -1 0 876 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_817
timestamp 1607101874
transform -1 0 972 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_437
timestamp 1607101874
transform 1 0 972 0 1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_361
timestamp 1607101874
transform -1 0 1092 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_362
timestamp 1607101874
transform 1 0 1092 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_516
timestamp 1607101874
transform 1 0 1116 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_242
timestamp 1607101874
transform -1 0 1236 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1021
timestamp 1607101874
transform 1 0 1236 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_139
timestamp 1607101874
transform 1 0 1332 0 1 2105
box -2 -3 18 103
use FILL  FILL_21_2_0
timestamp 1607101874
transform -1 0 1356 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1607101874
transform -1 0 1364 0 1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_126
timestamp 1607101874
transform -1 0 1412 0 1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_1071
timestamp 1607101874
transform 1 0 1412 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_438
timestamp 1607101874
transform 1 0 1444 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_551
timestamp 1607101874
transform 1 0 1540 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_3
timestamp 1607101874
transform 1 0 1572 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_496
timestamp 1607101874
transform -1 0 1612 0 1 2105
box -2 -3 26 103
use INVX2  INVX2_12
timestamp 1607101874
transform -1 0 1628 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_184
timestamp 1607101874
transform 1 0 1628 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1607101874
transform -1 0 1676 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_73
timestamp 1607101874
transform -1 0 1708 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1510
timestamp 1607101874
transform -1 0 1740 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_517
timestamp 1607101874
transform -1 0 1836 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_662
timestamp 1607101874
transform -1 0 1868 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_3_0
timestamp 1607101874
transform 1 0 1868 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1607101874
transform 1 0 1876 0 1 2105
box -2 -3 10 103
use INVX1  INVX1_137
timestamp 1607101874
transform 1 0 1884 0 1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_124
timestamp 1607101874
transform 1 0 1900 0 1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_1010
timestamp 1607101874
transform 1 0 1948 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1019
timestamp 1607101874
transform -1 0 2076 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_59
timestamp 1607101874
transform -1 0 2108 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_258
timestamp 1607101874
transform -1 0 2140 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_256
timestamp 1607101874
transform -1 0 2172 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_242
timestamp 1607101874
transform 1 0 2172 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_225
timestamp 1607101874
transform -1 0 2236 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_185
timestamp 1607101874
transform -1 0 2260 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_311
timestamp 1607101874
transform 1 0 2260 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_688
timestamp 1607101874
transform 1 0 2292 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_267
timestamp 1607101874
transform 1 0 2324 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_241
timestamp 1607101874
transform 1 0 2356 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_4_0
timestamp 1607101874
transform -1 0 2396 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1607101874
transform -1 0 2404 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_271
timestamp 1607101874
transform -1 0 2436 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1607101874
transform 1 0 2436 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1607101874
transform -1 0 2492 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_279
timestamp 1607101874
transform -1 0 2524 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_290
timestamp 1607101874
transform 1 0 2524 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1607101874
transform 1 0 2556 0 1 2105
box -2 -3 18 103
use INVX8  INVX8_30
timestamp 1607101874
transform 1 0 2572 0 1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_14
timestamp 1607101874
transform 1 0 2612 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_287
timestamp 1607101874
transform -1 0 2668 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_266
timestamp 1607101874
transform 1 0 2668 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_264
timestamp 1607101874
transform 1 0 2700 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_284
timestamp 1607101874
transform -1 0 2764 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_18
timestamp 1607101874
transform 1 0 2764 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_265
timestamp 1607101874
transform 1 0 2796 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_197
timestamp 1607101874
transform 1 0 2828 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_5_0
timestamp 1607101874
transform 1 0 2852 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1607101874
transform 1 0 2860 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1607101874
transform 1 0 2868 0 1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_406
timestamp 1607101874
transform 1 0 2964 0 1 2105
box -2 -3 50 103
use INVX1  INVX1_460
timestamp 1607101874
transform -1 0 3028 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_577
timestamp 1607101874
transform 1 0 3028 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_17
timestamp 1607101874
transform 1 0 3124 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_291
timestamp 1607101874
transform -1 0 3188 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_234
timestamp 1607101874
transform 1 0 3188 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_644
timestamp 1607101874
transform 1 0 3220 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_228
timestamp 1607101874
transform -1 0 3284 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_709
timestamp 1607101874
transform 1 0 3284 0 1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_190
timestamp 1607101874
transform -1 0 3364 0 1 2105
box -2 -3 50 103
use BUFX4  BUFX4_245
timestamp 1607101874
transform -1 0 3396 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_6_0
timestamp 1607101874
transform 1 0 3396 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1607101874
transform 1 0 3404 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_281
timestamp 1607101874
transform 1 0 3412 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_222
timestamp 1607101874
transform -1 0 3476 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_223
timestamp 1607101874
transform 1 0 3476 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_231
timestamp 1607101874
transform -1 0 3540 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_277
timestamp 1607101874
transform 1 0 3540 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_289
timestamp 1607101874
transform -1 0 3604 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_238
timestamp 1607101874
transform -1 0 3636 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_240
timestamp 1607101874
transform 1 0 3636 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_352
timestamp 1607101874
transform 1 0 3668 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_345
timestamp 1607101874
transform 1 0 3764 0 1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_311
timestamp 1607101874
transform -1 0 3828 0 1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_914
timestamp 1607101874
transform 1 0 3828 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_275
timestamp 1607101874
transform -1 0 3884 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_229
timestamp 1607101874
transform -1 0 3932 0 1 2105
box -2 -3 50 103
use FILL  FILL_21_7_0
timestamp 1607101874
transform -1 0 3940 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_7_1
timestamp 1607101874
transform -1 0 3948 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_729
timestamp 1607101874
transform -1 0 3980 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1607101874
transform 1 0 3980 0 1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_310
timestamp 1607101874
transform 1 0 4012 0 1 2105
box -2 -3 50 103
use INVX1  INVX1_296
timestamp 1607101874
transform -1 0 4076 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_351
timestamp 1607101874
transform -1 0 4172 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_274
timestamp 1607101874
transform -1 0 4196 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_913
timestamp 1607101874
transform -1 0 4228 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_728
timestamp 1607101874
transform -1 0 4260 0 1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_306
timestamp 1607101874
transform -1 0 4308 0 1 2105
box -2 -3 50 103
use INVX1  INVX1_294
timestamp 1607101874
transform -1 0 4324 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_359
timestamp 1607101874
transform -1 0 4420 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_8_0
timestamp 1607101874
transform -1 0 4428 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_8_1
timestamp 1607101874
transform -1 0 4436 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_568
timestamp 1607101874
transform -1 0 4468 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_452
timestamp 1607101874
transform 1 0 4468 0 1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_309
timestamp 1607101874
transform -1 0 4532 0 1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_350
timestamp 1607101874
transform -1 0 4628 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_629
timestamp 1607101874
transform -1 0 4660 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_281
timestamp 1607101874
transform -1 0 4676 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_421
timestamp 1607101874
transform 1 0 4676 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_422
timestamp 1607101874
transform -1 0 4740 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1607101874
transform 1 0 4740 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_303
timestamp 1607101874
transform 1 0 4836 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_294
timestamp 1607101874
transform 1 0 4868 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_197
timestamp 1607101874
transform -1 0 4924 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_364
timestamp 1607101874
transform 1 0 4924 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_9_0
timestamp 1607101874
transform 1 0 4956 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_9_1
timestamp 1607101874
transform 1 0 4964 0 1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_196
timestamp 1607101874
transform 1 0 4972 0 1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_170
timestamp 1607101874
transform 1 0 5020 0 1 2105
box -2 -3 50 103
use INVX1  INVX1_275
timestamp 1607101874
transform -1 0 5084 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_203
timestamp 1607101874
transform -1 0 5108 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_51
timestamp 1607101874
transform 1 0 5108 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1607101874
transform 1 0 5140 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_291
timestamp 1607101874
transform -1 0 5196 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_346
timestamp 1607101874
transform -1 0 5292 0 1 2105
box -2 -3 98 103
use FILL  FILL_22_1
timestamp 1607101874
transform 1 0 5292 0 1 2105
box -2 -3 10 103
use FILL  FILL_22_2
timestamp 1607101874
transform 1 0 5300 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_542
timestamp 1607101874
transform 1 0 4 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_441
timestamp 1607101874
transform 1 0 100 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_393
timestamp 1607101874
transform -1 0 164 0 -1 2305
box -2 -3 50 103
use NOR2X1  NOR2X1_242
timestamp 1607101874
transform -1 0 188 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_153
timestamp 1607101874
transform -1 0 220 0 -1 2305
box -2 -3 34 103
use AND2X2  AND2X2_55
timestamp 1607101874
transform 1 0 220 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_492
timestamp 1607101874
transform 1 0 252 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1174
timestamp 1607101874
transform 1 0 284 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_0_0
timestamp 1607101874
transform -1 0 324 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1607101874
transform -1 0 332 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_260
timestamp 1607101874
transform -1 0 380 0 -1 2305
box -2 -3 50 103
use AOI21X1  AOI21X1_154
timestamp 1607101874
transform 1 0 380 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_152
timestamp 1607101874
transform 1 0 412 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_241
timestamp 1607101874
transform -1 0 468 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1039
timestamp 1607101874
transform 1 0 468 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_531
timestamp 1607101874
transform 1 0 564 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_261
timestamp 1607101874
transform 1 0 660 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_389
timestamp 1607101874
transform -1 0 724 0 -1 2305
box -2 -3 50 103
use AND2X2  AND2X2_37
timestamp 1607101874
transform 1 0 724 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1006
timestamp 1607101874
transform 1 0 756 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_616
timestamp 1607101874
transform 1 0 788 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_728
timestamp 1607101874
transform -1 0 844 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_1_0
timestamp 1607101874
transform 1 0 844 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1607101874
transform 1 0 852 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_539
timestamp 1607101874
transform 1 0 860 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_243
timestamp 1607101874
transform -1 0 1004 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_254
timestamp 1607101874
transform -1 0 1052 0 -1 2305
box -2 -3 50 103
use AOI21X1  AOI21X1_68
timestamp 1607101874
transform 1 0 1052 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_121
timestamp 1607101874
transform -1 0 1108 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_823
timestamp 1607101874
transform 1 0 1108 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1508
timestamp 1607101874
transform 1 0 1204 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1507
timestamp 1607101874
transform -1 0 1268 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_232
timestamp 1607101874
transform -1 0 1292 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_392
timestamp 1607101874
transform 1 0 1292 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_459
timestamp 1607101874
transform 1 0 1316 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_2_0
timestamp 1607101874
transform 1 0 1348 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1607101874
transform 1 0 1356 0 -1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_342
timestamp 1607101874
transform 1 0 1364 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_605
timestamp 1607101874
transform 1 0 1396 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_182
timestamp 1607101874
transform -1 0 1452 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_281
timestamp 1607101874
transform 1 0 1452 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_239
timestamp 1607101874
transform -1 0 1508 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_309
timestamp 1607101874
transform 1 0 1508 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_308
timestamp 1607101874
transform -1 0 1572 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1025
timestamp 1607101874
transform -1 0 1668 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1509
timestamp 1607101874
transform 1 0 1668 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_304
timestamp 1607101874
transform 1 0 1700 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_305
timestamp 1607101874
transform -1 0 1764 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1023
timestamp 1607101874
transform 1 0 1764 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_283
timestamp 1607101874
transform 1 0 1860 0 -1 2305
box -2 -3 18 103
use FILL  FILL_22_3_0
timestamp 1607101874
transform 1 0 1876 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1607101874
transform 1 0 1884 0 -1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_300
timestamp 1607101874
transform 1 0 1892 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_73
timestamp 1607101874
transform 1 0 1924 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_149
timestamp 1607101874
transform -1 0 1972 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_168
timestamp 1607101874
transform 1 0 1972 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1347
timestamp 1607101874
transform 1 0 1996 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_324
timestamp 1607101874
transform 1 0 2028 0 -1 2305
box -2 -3 98 103
use BUFX4  BUFX4_32
timestamp 1607101874
transform 1 0 2124 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_424
timestamp 1607101874
transform 1 0 2156 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_165
timestamp 1607101874
transform -1 0 2220 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_230
timestamp 1607101874
transform -1 0 2252 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_253
timestamp 1607101874
transform 1 0 2252 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_708
timestamp 1607101874
transform 1 0 2284 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1607101874
transform 1 0 2316 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_11
timestamp 1607101874
transform 1 0 2348 0 -1 2305
box -2 -3 42 103
use FILL  FILL_22_4_0
timestamp 1607101874
transform -1 0 2396 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1607101874
transform -1 0 2404 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_268
timestamp 1607101874
transform -1 0 2436 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_394
timestamp 1607101874
transform -1 0 2468 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_441
timestamp 1607101874
transform 1 0 2468 0 -1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_25
timestamp 1607101874
transform -1 0 2540 0 -1 2305
box -2 -3 42 103
use BUFX4  BUFX4_211
timestamp 1607101874
transform -1 0 2572 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_28
timestamp 1607101874
transform -1 0 2612 0 -1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_101
timestamp 1607101874
transform 1 0 2612 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_38
timestamp 1607101874
transform -1 0 2660 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_393
timestamp 1607101874
transform 1 0 2660 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_171
timestamp 1607101874
transform -1 0 2716 0 -1 2305
box -2 -3 26 103
use OAI22X1  OAI22X1_50
timestamp 1607101874
transform -1 0 2756 0 -1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_218
timestamp 1607101874
transform 1 0 2756 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_248
timestamp 1607101874
transform -1 0 2828 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_396
timestamp 1607101874
transform 1 0 2828 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1175
timestamp 1607101874
transform 1 0 2860 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_5_0
timestamp 1607101874
transform -1 0 2900 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1607101874
transform -1 0 2908 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_51
timestamp 1607101874
transform -1 0 2940 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_279
timestamp 1607101874
transform -1 0 2964 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_50
timestamp 1607101874
transform -1 0 2996 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1607101874
transform -1 0 3028 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_49
timestamp 1607101874
transform 1 0 3028 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1607101874
transform -1 0 3092 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_391
timestamp 1607101874
transform 1 0 3092 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_392
timestamp 1607101874
transform 1 0 3124 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_390
timestamp 1607101874
transform 1 0 3156 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_199
timestamp 1607101874
transform -1 0 3236 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_994
timestamp 1607101874
transform 1 0 3236 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1607101874
transform 1 0 3268 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_213
timestamp 1607101874
transform -1 0 3324 0 -1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_78
timestamp 1607101874
transform 1 0 3324 0 -1 2305
box -2 -3 74 103
use FILL  FILL_22_6_0
timestamp 1607101874
transform -1 0 3404 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1607101874
transform -1 0 3412 0 -1 2305
box -2 -3 10 103
use AND2X2  AND2X2_54
timestamp 1607101874
transform -1 0 3444 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_388
timestamp 1607101874
transform -1 0 3476 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_339
timestamp 1607101874
transform -1 0 3508 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_262
timestamp 1607101874
transform 1 0 3508 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_29
timestamp 1607101874
transform -1 0 3556 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_747
timestamp 1607101874
transform 1 0 3556 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1607101874
transform -1 0 3628 0 -1 2305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_348
timestamp 1607101874
transform 1 0 3628 0 -1 2305
box -2 -3 98 103
use AND2X2  AND2X2_27
timestamp 1607101874
transform 1 0 3724 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_437
timestamp 1607101874
transform 1 0 3756 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_331
timestamp 1607101874
transform -1 0 3876 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_730
timestamp 1607101874
transform -1 0 3908 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_416
timestamp 1607101874
transform -1 0 3932 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_7_0
timestamp 1607101874
transform -1 0 3940 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_7_1
timestamp 1607101874
transform -1 0 3948 0 -1 2305
box -2 -3 10 103
use AND2X2  AND2X2_35
timestamp 1607101874
transform -1 0 3980 0 -1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_28
timestamp 1607101874
transform -1 0 4020 0 -1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_450
timestamp 1607101874
transform 1 0 4020 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_356
timestamp 1607101874
transform 1 0 4044 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1328
timestamp 1607101874
transform 1 0 4140 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1327
timestamp 1607101874
transform -1 0 4204 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_319
timestamp 1607101874
transform 1 0 4204 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1607101874
transform 1 0 4236 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1323
timestamp 1607101874
transform 1 0 4260 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1324
timestamp 1607101874
transform -1 0 4324 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_354
timestamp 1607101874
transform 1 0 4324 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_175
timestamp 1607101874
transform -1 0 4444 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_8_0
timestamp 1607101874
transform -1 0 4452 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_8_1
timestamp 1607101874
transform -1 0 4460 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_567
timestamp 1607101874
transform -1 0 4492 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_257
timestamp 1607101874
transform 1 0 4492 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_256
timestamp 1607101874
transform -1 0 4556 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_30
timestamp 1607101874
transform 1 0 4556 0 -1 2305
box -2 -3 50 103
use INVX1  INVX1_38
timestamp 1607101874
transform -1 0 4620 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_679
timestamp 1607101874
transform -1 0 4716 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_305
timestamp 1607101874
transform 1 0 4716 0 -1 2305
box -2 -3 50 103
use INVX1  INVX1_230
timestamp 1607101874
transform -1 0 4780 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_415
timestamp 1607101874
transform 1 0 4780 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1607101874
transform -1 0 4828 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_20
timestamp 1607101874
transform -1 0 4860 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_676
timestamp 1607101874
transform -1 0 4956 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_9_0
timestamp 1607101874
transform 1 0 4956 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_9_1
timestamp 1607101874
transform 1 0 4964 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_313
timestamp 1607101874
transform 1 0 4972 0 -1 2305
box -2 -3 50 103
use INVX1  INVX1_231
timestamp 1607101874
transform -1 0 5036 0 -1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_96
timestamp 1607101874
transform 1 0 5036 0 -1 2305
box -2 -3 74 103
use NOR2X1  NOR2X1_297
timestamp 1607101874
transform -1 0 5132 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_200
timestamp 1607101874
transform -1 0 5164 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_429
timestamp 1607101874
transform 1 0 5164 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_4
timestamp 1607101874
transform -1 0 5284 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1607101874
transform -1 0 5300 0 -1 2305
box -2 -3 18 103
use FILL  FILL_23_1
timestamp 1607101874
transform -1 0 5308 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_534
timestamp 1607101874
transform 1 0 4 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_440
timestamp 1607101874
transform 1 0 100 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_1173
timestamp 1607101874
transform 1 0 116 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_391
timestamp 1607101874
transform 1 0 148 0 1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1040
timestamp 1607101874
transform 1 0 196 0 1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_493
timestamp 1607101874
transform -1 0 324 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_0_0
timestamp 1607101874
transform 1 0 324 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1607101874
transform 1 0 332 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1041
timestamp 1607101874
transform 1 0 340 0 1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_243
timestamp 1607101874
transform 1 0 436 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_459
timestamp 1607101874
transform 1 0 460 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_520
timestamp 1607101874
transform 1 0 492 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_321
timestamp 1607101874
transform 1 0 516 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1043
timestamp 1607101874
transform 1 0 548 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_657
timestamp 1607101874
transform 1 0 644 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_331
timestamp 1607101874
transform -1 0 700 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1081
timestamp 1607101874
transform -1 0 732 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_658
timestamp 1607101874
transform 1 0 732 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_311
timestamp 1607101874
transform 1 0 764 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1044
timestamp 1607101874
transform 1 0 796 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_1_0
timestamp 1607101874
transform 1 0 892 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1607101874
transform 1 0 900 0 1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_245
timestamp 1607101874
transform 1 0 908 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_323
timestamp 1607101874
transform 1 0 932 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_322
timestamp 1607101874
transform -1 0 996 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1075
timestamp 1607101874
transform 1 0 996 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_535
timestamp 1607101874
transform 1 0 1028 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1522
timestamp 1607101874
transform 1 0 1124 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1521
timestamp 1607101874
transform 1 0 1156 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1498
timestamp 1607101874
transform 1 0 1188 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_503
timestamp 1607101874
transform 1 0 1220 0 1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_389
timestamp 1607101874
transform 1 0 1316 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_2_0
timestamp 1607101874
transform -1 0 1356 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1607101874
transform -1 0 1364 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_891
timestamp 1607101874
transform -1 0 1396 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_386
timestamp 1607101874
transform -1 0 1428 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_216
timestamp 1607101874
transform 1 0 1428 0 1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_79
timestamp 1607101874
transform 1 0 1476 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_76
timestamp 1607101874
transform -1 0 1524 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_327
timestamp 1607101874
transform -1 0 1556 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_182
timestamp 1607101874
transform -1 0 1604 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_606
timestamp 1607101874
transform -1 0 1636 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_15
timestamp 1607101874
transform 1 0 1636 0 1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_201
timestamp 1607101874
transform -1 0 1700 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_221
timestamp 1607101874
transform 1 0 1700 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_77
timestamp 1607101874
transform 1 0 1724 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_120
timestamp 1607101874
transform 1 0 1748 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_371
timestamp 1607101874
transform 1 0 1772 0 1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_320
timestamp 1607101874
transform 1 0 1788 0 1 2305
box -2 -3 50 103
use AOI21X1  AOI21X1_411
timestamp 1607101874
transform 1 0 1836 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_3_0
timestamp 1607101874
transform -1 0 1876 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1607101874
transform -1 0 1884 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_947
timestamp 1607101874
transform -1 0 1916 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_320
timestamp 1607101874
transform -1 0 2012 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1355
timestamp 1607101874
transform 1 0 2012 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1354
timestamp 1607101874
transform -1 0 2076 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1346
timestamp 1607101874
transform 1 0 2076 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_282
timestamp 1607101874
transform -1 0 2132 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_896
timestamp 1607101874
transform 1 0 2132 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_412
timestamp 1607101874
transform -1 0 2196 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_259
timestamp 1607101874
transform -1 0 2228 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_423
timestamp 1607101874
transform -1 0 2260 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_26
timestamp 1607101874
transform 1 0 2260 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_261
timestamp 1607101874
transform -1 0 2332 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_234
timestamp 1607101874
transform 1 0 2332 0 1 2305
box -2 -3 50 103
use FILL  FILL_23_4_0
timestamp 1607101874
transform -1 0 2388 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1607101874
transform -1 0 2396 0 1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_180
timestamp 1607101874
transform -1 0 2444 0 1 2305
box -2 -3 50 103
use BUFX4  BUFX4_244
timestamp 1607101874
transform 1 0 2444 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_27
timestamp 1607101874
transform -1 0 2508 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_29
timestamp 1607101874
transform 1 0 2508 0 1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_89
timestamp 1607101874
transform -1 0 2572 0 1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_223
timestamp 1607101874
transform -1 0 2620 0 1 2305
box -2 -3 50 103
use NAND3X1  NAND3X1_75
timestamp 1607101874
transform -1 0 2652 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_519
timestamp 1607101874
transform -1 0 2676 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_771
timestamp 1607101874
transform 1 0 2676 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_338
timestamp 1607101874
transform -1 0 2740 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1128
timestamp 1607101874
transform 1 0 2740 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_524
timestamp 1607101874
transform -1 0 2796 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_23
timestamp 1607101874
transform -1 0 2836 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_1221
timestamp 1607101874
transform 1 0 2836 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_14
timestamp 1607101874
transform -1 0 2908 0 1 2305
box -2 -3 42 103
use FILL  FILL_23_5_0
timestamp 1607101874
transform 1 0 2908 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1607101874
transform 1 0 2916 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_1082
timestamp 1607101874
transform 1 0 2924 0 1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_48
timestamp 1607101874
transform -1 0 2996 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_413
timestamp 1607101874
transform 1 0 2996 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_425
timestamp 1607101874
transform 1 0 3028 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_25
timestamp 1607101874
transform 1 0 3060 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_950
timestamp 1607101874
transform 1 0 3100 0 1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_42
timestamp 1607101874
transform 1 0 3132 0 1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_28
timestamp 1607101874
transform 1 0 3172 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_283
timestamp 1607101874
transform 1 0 3212 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_17
timestamp 1607101874
transform 1 0 3244 0 1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_191
timestamp 1607101874
transform 1 0 3284 0 1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_317
timestamp 1607101874
transform -1 0 3356 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_907
timestamp 1607101874
transform -1 0 3388 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_908
timestamp 1607101874
transform -1 0 3420 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_6_0
timestamp 1607101874
transform 1 0 3420 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1607101874
transform 1 0 3428 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_317
timestamp 1607101874
transform 1 0 3436 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_18
timestamp 1607101874
transform -1 0 3508 0 1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_33
timestamp 1607101874
transform -1 0 3548 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_461
timestamp 1607101874
transform -1 0 3580 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_255
timestamp 1607101874
transform -1 0 3628 0 1 2305
box -2 -3 50 103
use AOI21X1  AOI21X1_346
timestamp 1607101874
transform 1 0 3628 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_392
timestamp 1607101874
transform 1 0 3660 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_357
timestamp 1607101874
transform 1 0 3692 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_820
timestamp 1607101874
transform -1 0 3756 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_819
timestamp 1607101874
transform 1 0 3756 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_792
timestamp 1607101874
transform -1 0 3820 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_733
timestamp 1607101874
transform 1 0 3820 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_321
timestamp 1607101874
transform -1 0 3884 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_393
timestamp 1607101874
transform -1 0 3916 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_7_0
timestamp 1607101874
transform 1 0 3916 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_7_1
timestamp 1607101874
transform 1 0 3924 0 1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_653
timestamp 1607101874
transform 1 0 3932 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_541
timestamp 1607101874
transform -1 0 3988 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_547
timestamp 1607101874
transform 1 0 3988 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_659
timestamp 1607101874
transform 1 0 4020 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_417
timestamp 1607101874
transform -1 0 4076 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_299
timestamp 1607101874
transform 1 0 4076 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_45
timestamp 1607101874
transform -1 0 4124 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_419
timestamp 1607101874
transform -1 0 4156 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_416
timestamp 1607101874
transform -1 0 4188 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_355
timestamp 1607101874
transform -1 0 4284 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1326
timestamp 1607101874
transform 1 0 4284 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1325
timestamp 1607101874
transform -1 0 4348 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_446
timestamp 1607101874
transform -1 0 4380 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1607101874
transform 1 0 4380 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_3
timestamp 1607101874
transform 1 0 4404 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_8_0
timestamp 1607101874
transform -1 0 4444 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_8_1
timestamp 1607101874
transform -1 0 4452 0 1 2305
box -2 -3 10 103
use BUFX4  BUFX4_418
timestamp 1607101874
transform -1 0 4484 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_660
timestamp 1607101874
transform -1 0 4508 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_548
timestamp 1607101874
transform -1 0 4540 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_332
timestamp 1607101874
transform -1 0 4636 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_194
timestamp 1607101874
transform -1 0 4660 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_45
timestamp 1607101874
transform -1 0 4684 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1607101874
transform -1 0 4716 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_675
timestamp 1607101874
transform -1 0 4812 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_809
timestamp 1607101874
transform -1 0 4844 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_358
timestamp 1607101874
transform -1 0 4940 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_9_0
timestamp 1607101874
transform 1 0 4940 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_9_1
timestamp 1607101874
transform 1 0 4948 0 1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_314
timestamp 1607101874
transform 1 0 4956 0 1 2305
box -2 -3 50 103
use INVX1  INVX1_295
timestamp 1607101874
transform -1 0 5020 0 1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_347
timestamp 1607101874
transform 1 0 5020 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1607101874
transform -1 0 5212 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_1084
timestamp 1607101874
transform 1 0 5212 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_723
timestamp 1607101874
transform 1 0 5244 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1083
timestamp 1607101874
transform -1 0 5308 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_530
timestamp 1607101874
transform 1 0 4 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1520
timestamp 1607101874
transform 1 0 100 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_340
timestamp 1607101874
transform -1 0 156 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1519
timestamp 1607101874
transform -1 0 188 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_538
timestamp 1607101874
transform 1 0 188 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1528
timestamp 1607101874
transform 1 0 284 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1527
timestamp 1607101874
transform -1 0 348 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_0_0
timestamp 1607101874
transform -1 0 356 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1607101874
transform -1 0 364 0 -1 2505
box -2 -3 10 103
use BUFX4  BUFX4_310
timestamp 1607101874
transform -1 0 396 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_445
timestamp 1607101874
transform 1 0 396 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_1260
timestamp 1607101874
transform 1 0 412 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1261
timestamp 1607101874
transform 1 0 444 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_313
timestamp 1607101874
transform 1 0 476 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_156
timestamp 1607101874
transform 1 0 508 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_246
timestamp 1607101874
transform -1 0 564 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_320
timestamp 1607101874
transform 1 0 564 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_382
timestamp 1607101874
transform 1 0 596 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_313
timestamp 1607101874
transform 1 0 620 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_312
timestamp 1607101874
transform 1 0 652 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_381
timestamp 1607101874
transform 1 0 684 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_9
timestamp 1607101874
transform -1 0 748 0 -1 2505
box -2 -3 42 103
use MUX2X1  MUX2X1_215
timestamp 1607101874
transform 1 0 748 0 -1 2505
box -2 -3 50 103
use NAND2X1  NAND2X1_209
timestamp 1607101874
transform -1 0 820 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_659
timestamp 1607101874
transform -1 0 852 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_1_0
timestamp 1607101874
transform 1 0 852 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1607101874
transform 1 0 860 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_888
timestamp 1607101874
transform 1 0 868 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_300
timestamp 1607101874
transform -1 0 932 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_890
timestamp 1607101874
transform -1 0 964 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_889
timestamp 1607101874
transform 1 0 964 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_517
timestamp 1607101874
transform 1 0 996 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_80
timestamp 1607101874
transform 1 0 1020 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1074
timestamp 1607101874
transform 1 0 1052 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1005
timestamp 1607101874
transform 1 0 1084 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1497
timestamp 1607101874
transform 1 0 1180 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1504
timestamp 1607101874
transform 1 0 1212 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1503
timestamp 1607101874
transform 1 0 1244 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_506
timestamp 1607101874
transform 1 0 1276 0 -1 2505
box -2 -3 98 103
use FILL  FILL_24_2_0
timestamp 1607101874
transform 1 0 1372 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1607101874
transform 1 0 1380 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_78
timestamp 1607101874
transform 1 0 1388 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_566
timestamp 1607101874
transform 1 0 1412 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1169
timestamp 1607101874
transform 1 0 1436 0 -1 2505
box -2 -3 34 103
use INVX8  INVX8_25
timestamp 1607101874
transform -1 0 1508 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_469
timestamp 1607101874
transform 1 0 1508 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_357
timestamp 1607101874
transform 1 0 1540 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_186
timestamp 1607101874
transform -1 0 1620 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_664
timestamp 1607101874
transform 1 0 1620 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_312
timestamp 1607101874
transform 1 0 1652 0 -1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_610
timestamp 1607101874
transform 1 0 1748 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_609
timestamp 1607101874
transform 1 0 1780 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_721
timestamp 1607101874
transform -1 0 1836 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1257
timestamp 1607101874
transform -1 0 1868 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_3_0
timestamp 1607101874
transform 1 0 1868 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1607101874
transform 1 0 1876 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_946
timestamp 1607101874
transform 1 0 1884 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_564
timestamp 1607101874
transform 1 0 1916 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1168
timestamp 1607101874
transform 1 0 1940 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_489
timestamp 1607101874
transform 1 0 1972 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_490
timestamp 1607101874
transform -1 0 2036 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_482
timestamp 1607101874
transform 1 0 2036 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_385
timestamp 1607101874
transform -1 0 2084 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_302
timestamp 1607101874
transform -1 0 2116 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1262
timestamp 1607101874
transform 1 0 2116 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_82
timestamp 1607101874
transform -1 0 2180 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_285
timestamp 1607101874
transform -1 0 2212 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_288
timestamp 1607101874
transform -1 0 2244 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_243
timestamp 1607101874
transform -1 0 2276 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_242
timestamp 1607101874
transform 1 0 2276 0 -1 2505
box -2 -3 50 103
use BUFX4  BUFX4_224
timestamp 1607101874
transform 1 0 2324 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_698
timestamp 1607101874
transform -1 0 2388 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_4_0
timestamp 1607101874
transform -1 0 2396 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1607101874
transform -1 0 2404 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_1016
timestamp 1607101874
transform -1 0 2436 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_167
timestamp 1607101874
transform -1 0 2468 0 -1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_38
timestamp 1607101874
transform -1 0 2540 0 -1 2505
box -2 -3 74 103
use NOR2X1  NOR2X1_576
timestamp 1607101874
transform -1 0 2564 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_728
timestamp 1607101874
transform 1 0 2564 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_310
timestamp 1607101874
transform -1 0 2684 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_81
timestamp 1607101874
transform -1 0 2724 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_31
timestamp 1607101874
transform -1 0 2764 0 -1 2505
box -2 -3 42 103
use OAI22X1  OAI22X1_60
timestamp 1607101874
transform -1 0 2804 0 -1 2505
box -2 -3 42 103
use INVX8  INVX8_33
timestamp 1607101874
transform -1 0 2844 0 -1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_397
timestamp 1607101874
transform 1 0 2844 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1200
timestamp 1607101874
transform -1 0 2908 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_5_0
timestamp 1607101874
transform 1 0 2908 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1607101874
transform 1 0 2916 0 -1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_473
timestamp 1607101874
transform 1 0 2924 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_24
timestamp 1607101874
transform -1 0 2988 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_1107
timestamp 1607101874
transform -1 0 3020 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_280
timestamp 1607101874
transform -1 0 3052 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_253
timestamp 1607101874
transform 1 0 3052 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_272
timestamp 1607101874
transform 1 0 3084 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_207
timestamp 1607101874
transform 1 0 3116 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_1263
timestamp 1607101874
transform -1 0 3196 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_391
timestamp 1607101874
transform -1 0 3228 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_548
timestamp 1607101874
transform -1 0 3252 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_600
timestamp 1607101874
transform -1 0 3276 0 -1 2505
box -2 -3 26 103
use INVX4  INVX4_14
timestamp 1607101874
transform -1 0 3300 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_721
timestamp 1607101874
transform -1 0 3332 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_93
timestamp 1607101874
transform 1 0 3332 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_1264
timestamp 1607101874
transform 1 0 3372 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_6_0
timestamp 1607101874
transform 1 0 3404 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1607101874
transform 1 0 3412 0 -1 2505
box -2 -3 10 103
use OAI22X1  OAI22X1_94
timestamp 1607101874
transform 1 0 3420 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_1177
timestamp 1607101874
transform -1 0 3492 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1243
timestamp 1607101874
transform -1 0 3524 0 -1 2505
box -2 -3 34 103
use INVX4  INVX4_13
timestamp 1607101874
transform 1 0 3524 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1176
timestamp 1607101874
transform -1 0 3580 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1152
timestamp 1607101874
transform -1 0 3612 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_732
timestamp 1607101874
transform -1 0 3644 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_298
timestamp 1607101874
transform -1 0 3660 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_1049
timestamp 1607101874
transform -1 0 3692 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_276
timestamp 1607101874
transform -1 0 3716 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_818
timestamp 1607101874
transform -1 0 3748 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1607101874
transform 1 0 3748 0 -1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_316
timestamp 1607101874
transform 1 0 3772 0 -1 2505
box -2 -3 50 103
use INVX1  INVX1_297
timestamp 1607101874
transform -1 0 3836 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_731
timestamp 1607101874
transform 1 0 3836 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1334
timestamp 1607101874
transform -1 0 3900 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1335
timestamp 1607101874
transform -1 0 3932 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_7_0
timestamp 1607101874
transform -1 0 3940 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_7_1
timestamp 1607101874
transform -1 0 3948 0 -1 2505
box -2 -3 10 103
use BUFX4  BUFX4_409
timestamp 1607101874
transform -1 0 3980 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_413
timestamp 1607101874
transform -1 0 4012 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_414
timestamp 1607101874
transform -1 0 4044 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1607101874
transform 1 0 4044 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_320
timestamp 1607101874
transform -1 0 4100 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_49
timestamp 1607101874
transform -1 0 4124 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_373
timestamp 1607101874
transform 1 0 4124 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_789
timestamp 1607101874
transform 1 0 4156 0 -1 2505
box -2 -3 98 103
use OAI22X1  OAI22X1_86
timestamp 1607101874
transform 1 0 4252 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_1242
timestamp 1607101874
transform -1 0 4324 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_272
timestamp 1607101874
transform 1 0 4324 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_24
timestamp 1607101874
transform -1 0 4388 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_811
timestamp 1607101874
transform -1 0 4420 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_8_0
timestamp 1607101874
transform -1 0 4428 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_8_1
timestamp 1607101874
transform -1 0 4436 0 -1 2505
box -2 -3 10 103
use AND2X2  AND2X2_50
timestamp 1607101874
transform -1 0 4468 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_65
timestamp 1607101874
transform -1 0 4508 0 -1 2505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_339
timestamp 1607101874
transform -1 0 4604 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_810
timestamp 1607101874
transform -1 0 4636 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1607101874
transform 1 0 4636 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1607101874
transform -1 0 4692 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_85
timestamp 1607101874
transform 1 0 4692 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_1240
timestamp 1607101874
transform -1 0 4764 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_611
timestamp 1607101874
transform -1 0 4788 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_23
timestamp 1607101874
transform 1 0 4788 0 -1 2505
box -2 -3 42 103
use CLKBUF1  CLKBUF1_87
timestamp 1607101874
transform -1 0 4900 0 -1 2505
box -2 -3 74 103
use OAI21X1  OAI21X1_435
timestamp 1607101874
transform -1 0 4932 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_441
timestamp 1607101874
transform -1 0 4956 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_9_0
timestamp 1607101874
transform -1 0 4964 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_9_1
timestamp 1607101874
transform -1 0 4972 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_684
timestamp 1607101874
transform -1 0 5068 0 -1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_546
timestamp 1607101874
transform 1 0 5068 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_428
timestamp 1607101874
transform 1 0 5100 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_430
timestamp 1607101874
transform 1 0 5196 0 -1 2505
box -2 -3 98 103
use FILL  FILL_25_1
timestamp 1607101874
transform -1 0 5300 0 -1 2505
box -2 -3 10 103
use FILL  FILL_25_2
timestamp 1607101874
transform -1 0 5308 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1038
timestamp 1607101874
transform 1 0 4 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_319
timestamp 1607101874
transform 1 0 100 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_318
timestamp 1607101874
transform -1 0 164 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1037
timestamp 1607101874
transform 1 0 164 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_317
timestamp 1607101874
transform 1 0 260 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_316
timestamp 1607101874
transform -1 0 324 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_407
timestamp 1607101874
transform 1 0 324 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_0_0
timestamp 1607101874
transform 1 0 340 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1607101874
transform 1 0 348 0 1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_352
timestamp 1607101874
transform 1 0 356 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_510
timestamp 1607101874
transform 1 0 380 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_511
timestamp 1607101874
transform 1 0 412 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1079
timestamp 1607101874
transform 1 0 444 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1523
timestamp 1607101874
transform 1 0 476 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1047
timestamp 1607101874
transform 1 0 508 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1035
timestamp 1607101874
transform 1 0 604 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1011
timestamp 1607101874
transform -1 0 796 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_296
timestamp 1607101874
transform -1 0 828 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_297
timestamp 1607101874
transform -1 0 860 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_1_0
timestamp 1607101874
transform 1 0 860 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1607101874
transform 1 0 868 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1013
timestamp 1607101874
transform 1 0 876 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_301
timestamp 1607101874
transform 1 0 972 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_300
timestamp 1607101874
transform -1 0 1036 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_458
timestamp 1607101874
transform -1 0 1068 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_298
timestamp 1607101874
transform 1 0 1068 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_293
timestamp 1607101874
transform 1 0 1100 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_518
timestamp 1607101874
transform -1 0 1156 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_292
timestamp 1607101874
transform -1 0 1188 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_456
timestamp 1607101874
transform 1 0 1188 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_498
timestamp 1607101874
transform 1 0 1220 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1496
timestamp 1607101874
transform 1 0 1316 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_2_0
timestamp 1607101874
transform 1 0 1348 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1607101874
transform 1 0 1356 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_1495
timestamp 1607101874
transform 1 0 1364 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_389
timestamp 1607101874
transform -1 0 1428 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_567
timestamp 1607101874
transform -1 0 1452 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_457
timestamp 1607101874
transform 1 0 1452 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_265
timestamp 1607101874
transform 1 0 1484 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_610
timestamp 1607101874
transform 1 0 1500 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1607101874
transform 1 0 1532 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_294
timestamp 1607101874
transform 1 0 1556 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_295
timestamp 1607101874
transform 1 0 1588 0 1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_184
timestamp 1607101874
transform -1 0 1668 0 1 2505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1006
timestamp 1607101874
transform 1 0 1668 0 1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_722
timestamp 1607101874
transform -1 0 1788 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_510
timestamp 1607101874
transform 1 0 1788 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_3_0
timestamp 1607101874
transform -1 0 1892 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1607101874
transform -1 0 1900 0 1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_35
timestamp 1607101874
transform -1 0 1924 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_565
timestamp 1607101874
transform -1 0 1948 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_509
timestamp 1607101874
transform 1 0 1948 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_965
timestamp 1607101874
transform 1 0 2044 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_422
timestamp 1607101874
transform 1 0 2076 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_56
timestamp 1607101874
transform 1 0 2108 0 1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_16
timestamp 1607101874
transform -1 0 2212 0 1 2505
box -2 -3 74 103
use AOI21X1  AOI21X1_38
timestamp 1607101874
transform 1 0 2212 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_75
timestamp 1607101874
transform -1 0 2268 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_406
timestamp 1607101874
transform 1 0 2268 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_715
timestamp 1607101874
transform -1 0 2388 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_4_0
timestamp 1607101874
transform -1 0 2396 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1607101874
transform -1 0 2404 0 1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_308
timestamp 1607101874
transform -1 0 2428 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_342
timestamp 1607101874
transform -1 0 2452 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_720
timestamp 1607101874
transform 1 0 2452 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_50
timestamp 1607101874
transform 1 0 2548 0 1 2505
box -2 -3 18 103
use MUX2X1  MUX2X1_40
timestamp 1607101874
transform 1 0 2564 0 1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_827
timestamp 1607101874
transform 1 0 2612 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_361
timestamp 1607101874
transform -1 0 2676 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_81
timestamp 1607101874
transform 1 0 2676 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_42
timestamp 1607101874
transform -1 0 2732 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_538
timestamp 1607101874
transform -1 0 2756 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_370
timestamp 1607101874
transform 1 0 2756 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_568
timestamp 1607101874
transform -1 0 2812 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_88
timestamp 1607101874
transform -1 0 2844 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_92
timestamp 1607101874
transform -1 0 2876 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_81
timestamp 1607101874
transform -1 0 2908 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_5_0
timestamp 1607101874
transform -1 0 2916 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1607101874
transform -1 0 2924 0 1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_259
timestamp 1607101874
transform -1 0 2956 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_403
timestamp 1607101874
transform -1 0 2988 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1165
timestamp 1607101874
transform 1 0 2988 0 1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_66
timestamp 1607101874
transform -1 0 3060 0 1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_446
timestamp 1607101874
transform -1 0 3092 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_409
timestamp 1607101874
transform 1 0 3092 0 1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_12
timestamp 1607101874
transform -1 0 3164 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_676
timestamp 1607101874
transform 1 0 3164 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1607101874
transform 1 0 3196 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_170
timestamp 1607101874
transform -1 0 3252 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_286
timestamp 1607101874
transform 1 0 3252 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_275
timestamp 1607101874
transform -1 0 3316 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_270
timestamp 1607101874
transform -1 0 3348 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_239
timestamp 1607101874
transform -1 0 3380 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_282
timestamp 1607101874
transform -1 0 3412 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_6_0
timestamp 1607101874
transform 1 0 3412 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1607101874
transform 1 0 3420 0 1 2505
box -2 -3 10 103
use BUFX4  BUFX4_237
timestamp 1607101874
transform 1 0 3428 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_95
timestamp 1607101874
transform -1 0 3492 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_110
timestamp 1607101874
transform -1 0 3524 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_98
timestamp 1607101874
transform 1 0 3524 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_341
timestamp 1607101874
transform -1 0 3580 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_171
timestamp 1607101874
transform 1 0 3580 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_400
timestamp 1607101874
transform -1 0 3644 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_399
timestamp 1607101874
transform -1 0 3676 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_401
timestamp 1607101874
transform -1 0 3708 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_402
timestamp 1607101874
transform -1 0 3740 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_30
timestamp 1607101874
transform -1 0 3780 0 1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_445
timestamp 1607101874
transform -1 0 3812 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_343
timestamp 1607101874
transform -1 0 3908 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_7_0
timestamp 1607101874
transform -1 0 3916 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_7_1
timestamp 1607101874
transform -1 0 3924 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_335
timestamp 1607101874
transform -1 0 4020 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_190
timestamp 1607101874
transform 1 0 4020 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_415
timestamp 1607101874
transform -1 0 4084 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_411
timestamp 1607101874
transform 1 0 4084 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_102
timestamp 1607101874
transform 1 0 4116 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_273
timestamp 1607101874
transform 1 0 4140 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_313
timestamp 1607101874
transform 1 0 4164 0 1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_73
timestamp 1607101874
transform 1 0 4188 0 1 2505
box -2 -3 50 103
use INVX1  INVX1_83
timestamp 1607101874
transform 1 0 4236 0 1 2505
box -2 -3 18 103
use BUFX4  BUFX4_412
timestamp 1607101874
transform -1 0 4284 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_398
timestamp 1607101874
transform -1 0 4316 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1607101874
transform -1 0 4340 0 1 2505
box -2 -3 26 103
use INVX8  INVX8_18
timestamp 1607101874
transform 1 0 4340 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_44
timestamp 1607101874
transform -1 0 4404 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_410
timestamp 1607101874
transform -1 0 4436 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_8_0
timestamp 1607101874
transform 1 0 4436 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_8_1
timestamp 1607101874
transform 1 0 4444 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_1147
timestamp 1607101874
transform 1 0 4452 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_335
timestamp 1607101874
transform -1 0 4508 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_678
timestamp 1607101874
transform -1 0 4604 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_426
timestamp 1607101874
transform -1 0 4620 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_1241
timestamp 1607101874
transform -1 0 4652 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_680
timestamp 1607101874
transform -1 0 4748 0 1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_656
timestamp 1607101874
transform 1 0 4748 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_544
timestamp 1607101874
transform -1 0 4804 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_674
timestamp 1607101874
transform -1 0 4900 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_436
timestamp 1607101874
transform -1 0 4932 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_9_0
timestamp 1607101874
transform -1 0 4940 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_9_1
timestamp 1607101874
transform -1 0 4948 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1607101874
transform -1 0 5044 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_61
timestamp 1607101874
transform 1 0 5044 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_62
timestamp 1607101874
transform -1 0 5108 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_658
timestamp 1607101874
transform 1 0 5108 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_56
timestamp 1607101874
transform -1 0 5164 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_673
timestamp 1607101874
transform -1 0 5260 0 1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_624
timestamp 1607101874
transform -1 0 5284 0 1 2505
box -2 -3 26 103
use FILL  FILL_26_1
timestamp 1607101874
transform 1 0 5284 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_2
timestamp 1607101874
transform 1 0 5292 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_3
timestamp 1607101874
transform 1 0 5300 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_528
timestamp 1607101874
transform 1 0 4 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1516
timestamp 1607101874
transform 1 0 100 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_244
timestamp 1607101874
transform -1 0 156 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1515
timestamp 1607101874
transform -1 0 188 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_159
timestamp 1607101874
transform -1 0 220 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_249
timestamp 1607101874
transform -1 0 244 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_327
timestamp 1607101874
transform 1 0 244 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_326
timestamp 1607101874
transform -1 0 308 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_0_0
timestamp 1607101874
transform 1 0 308 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1607101874
transform 1 0 316 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1046
timestamp 1607101874
transform 1 0 324 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1524
timestamp 1607101874
transform 1 0 420 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_536
timestamp 1607101874
transform 1 0 452 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_791
timestamp 1607101874
transform -1 0 580 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_344
timestamp 1607101874
transform -1 0 612 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1004
timestamp 1607101874
transform 1 0 612 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_291
timestamp 1607101874
transform 1 0 708 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_459
timestamp 1607101874
transform 1 0 740 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_290
timestamp 1607101874
transform -1 0 796 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_341
timestamp 1607101874
transform 1 0 796 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_240
timestamp 1607101874
transform 1 0 812 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_457
timestamp 1607101874
transform -1 0 860 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_1_0
timestamp 1607101874
transform 1 0 860 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1607101874
transform 1 0 868 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_1500
timestamp 1607101874
transform 1 0 876 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1499
timestamp 1607101874
transform 1 0 908 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_458
timestamp 1607101874
transform 1 0 940 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_504
timestamp 1607101874
transform 1 0 964 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_434
timestamp 1607101874
transform 1 0 1060 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1513
timestamp 1607101874
transform -1 0 1116 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_786
timestamp 1607101874
transform 1 0 1116 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_435
timestamp 1607101874
transform 1 0 1148 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1489
timestamp 1607101874
transform 1 0 1172 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_496
timestamp 1607101874
transform -1 0 1300 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1492
timestamp 1607101874
transform 1 0 1300 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1491
timestamp 1607101874
transform -1 0 1364 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_2_0
timestamp 1607101874
transform 1 0 1364 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1607101874
transform 1 0 1372 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_341
timestamp 1607101874
transform 1 0 1380 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1493
timestamp 1607101874
transform 1 0 1412 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1494
timestamp 1607101874
transform -1 0 1476 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_497
timestamp 1607101874
transform 1 0 1476 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_227
timestamp 1607101874
transform 1 0 1572 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_143
timestamp 1607101874
transform 1 0 1596 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_485
timestamp 1607101874
transform -1 0 1652 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_966
timestamp 1607101874
transform 1 0 1652 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_226
timestamp 1607101874
transform 1 0 1684 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_73
timestamp 1607101874
transform 1 0 1708 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_264
timestamp 1607101874
transform 1 0 1732 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_609
timestamp 1607101874
transform -1 0 1780 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_621
timestamp 1607101874
transform 1 0 1780 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_79
timestamp 1607101874
transform -1 0 1828 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_606
timestamp 1607101874
transform 1 0 1828 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_718
timestamp 1607101874
transform -1 0 1884 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_502
timestamp 1607101874
transform 1 0 1900 0 -1 2705
box -2 -3 98 103
use BUFX4  BUFX4_318
timestamp 1607101874
transform -1 0 2028 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_483
timestamp 1607101874
transform -1 0 2052 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_77
timestamp 1607101874
transform -1 0 2076 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1015
timestamp 1607101874
transform -1 0 2108 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1014
timestamp 1607101874
transform 1 0 2108 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_249
timestamp 1607101874
transform 1 0 2140 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_74
timestamp 1607101874
transform -1 0 2188 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_250
timestamp 1607101874
transform -1 0 2212 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_707
timestamp 1607101874
transform 1 0 2212 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_18
timestamp 1607101874
transform 1 0 2244 0 -1 2705
box -2 -3 42 103
use MUX2X1  MUX2X1_39
timestamp 1607101874
transform 1 0 2284 0 -1 2705
box -2 -3 50 103
use INVX1  INVX1_49
timestamp 1607101874
transform -1 0 2348 0 -1 2705
box -2 -3 18 103
use FILL  FILL_26_4_0
timestamp 1607101874
transform -1 0 2356 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1607101874
transform -1 0 2364 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_719
timestamp 1607101874
transform -1 0 2460 0 -1 2705
box -2 -3 98 103
use BUFX4  BUFX4_365
timestamp 1607101874
transform 1 0 2460 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_724
timestamp 1607101874
transform 1 0 2492 0 -1 2705
box -2 -3 98 103
use BUFX4  BUFX4_89
timestamp 1607101874
transform -1 0 2620 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_77
timestamp 1607101874
transform 1 0 2620 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_74
timestamp 1607101874
transform 1 0 2652 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_33
timestamp 1607101874
transform 1 0 2684 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_91
timestamp 1607101874
transform -1 0 2740 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1607101874
transform -1 0 2756 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_716
timestamp 1607101874
transform 1 0 2756 0 -1 2705
box -2 -3 98 103
use BUFX4  BUFX4_90
timestamp 1607101874
transform -1 0 2884 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_5_0
timestamp 1607101874
transform 1 0 2884 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1607101874
transform 1 0 2892 0 -1 2705
box -2 -3 10 103
use BUFX4  BUFX4_78
timestamp 1607101874
transform 1 0 2900 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_188
timestamp 1607101874
transform -1 0 2964 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_76
timestamp 1607101874
transform -1 0 2996 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_80
timestamp 1607101874
transform 1 0 2996 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_11
timestamp 1607101874
transform -1 0 3060 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_16
timestamp 1607101874
transform 1 0 3060 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_99
timestamp 1607101874
transform 1 0 3092 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1607101874
transform -1 0 3156 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_84
timestamp 1607101874
transform 1 0 3156 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_94
timestamp 1607101874
transform -1 0 3220 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_87
timestamp 1607101874
transform 1 0 3220 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_101
timestamp 1607101874
transform 1 0 3252 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_15
timestamp 1607101874
transform -1 0 3316 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_109
timestamp 1607101874
transform 1 0 3316 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_97
timestamp 1607101874
transform -1 0 3380 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_79
timestamp 1607101874
transform 1 0 3380 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 2705
box -2 -3 10 103
use BUFX4  BUFX4_96
timestamp 1607101874
transform 1 0 3428 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1607101874
transform 1 0 3460 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_107
timestamp 1607101874
transform 1 0 3492 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_316
timestamp 1607101874
transform 1 0 3524 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_103
timestamp 1607101874
transform 1 0 3548 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1607101874
transform -1 0 3612 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_86
timestamp 1607101874
transform 1 0 3612 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1037
timestamp 1607101874
transform -1 0 3676 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_400
timestamp 1607101874
transform -1 0 3692 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_26
timestamp 1607101874
transform -1 0 3724 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_447
timestamp 1607101874
transform -1 0 3756 0 -1 2705
box -2 -3 34 103
use INVX4  INVX4_4
timestamp 1607101874
transform 1 0 3756 0 -1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_249
timestamp 1607101874
transform -1 0 3828 0 -1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_1036
timestamp 1607101874
transform -1 0 3860 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_315
timestamp 1607101874
transform -1 0 3884 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_31
timestamp 1607101874
transform 1 0 3884 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_7_0
timestamp 1607101874
transform 1 0 3916 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_7_1
timestamp 1607101874
transform 1 0 3924 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_108
timestamp 1607101874
transform 1 0 3932 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_801
timestamp 1607101874
transform -1 0 4052 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_88
timestamp 1607101874
transform -1 0 4068 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_797
timestamp 1607101874
transform -1 0 4164 0 -1 2705
box -2 -3 98 103
use MUX2X1  MUX2X1_78
timestamp 1607101874
transform -1 0 4212 0 -1 2705
box -2 -3 50 103
use MUX2X1  MUX2X1_248
timestamp 1607101874
transform 1 0 4212 0 -1 2705
box -2 -3 50 103
use BUFX4  BUFX4_395
timestamp 1607101874
transform 1 0 4260 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_228
timestamp 1607101874
transform -1 0 4340 0 -1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_912
timestamp 1607101874
transform -1 0 4372 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_343
timestamp 1607101874
transform -1 0 4388 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_1336
timestamp 1607101874
transform 1 0 4388 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_8_0
timestamp 1607101874
transform -1 0 4428 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_8_1
timestamp 1607101874
transform -1 0 4436 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_1337
timestamp 1607101874
transform -1 0 4468 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_257
timestamp 1607101874
transform 1 0 4468 0 -1 2705
box -2 -3 50 103
use NOR2X1  NOR2X1_48
timestamp 1607101874
transform 1 0 4516 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1607101874
transform -1 0 4572 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1607101874
transform 1 0 4572 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_298
timestamp 1607101874
transform 1 0 4668 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_22
timestamp 1607101874
transform -1 0 4724 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_302
timestamp 1607101874
transform 1 0 4724 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1148
timestamp 1607101874
transform -1 0 4788 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_610
timestamp 1607101874
transform -1 0 4812 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_57
timestamp 1607101874
transform -1 0 4844 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_58
timestamp 1607101874
transform -1 0 4876 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_440
timestamp 1607101874
transform -1 0 4900 0 -1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_32
timestamp 1607101874
transform 1 0 4900 0 -1 2705
box -2 -3 50 103
use FILL  FILL_26_9_0
timestamp 1607101874
transform -1 0 4956 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_9_1
timestamp 1607101874
transform -1 0 4964 0 -1 2705
box -2 -3 10 103
use INVX1  INVX1_40
timestamp 1607101874
transform -1 0 4980 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_682
timestamp 1607101874
transform -1 0 5076 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_392
timestamp 1607101874
transform -1 0 5092 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_330
timestamp 1607101874
transform -1 0 5188 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_431
timestamp 1607101874
transform 1 0 5188 0 -1 2705
box -2 -3 98 103
use FILL  FILL_27_1
timestamp 1607101874
transform -1 0 5292 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_2
timestamp 1607101874
transform -1 0 5300 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_3
timestamp 1607101874
transform -1 0 5308 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_532
timestamp 1607101874
transform 1 0 4 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_324
timestamp 1607101874
transform 1 0 100 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_790
timestamp 1607101874
transform 1 0 116 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1050
timestamp 1607101874
transform 1 0 148 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1036
timestamp 1607101874
transform 1 0 244 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_0_0
timestamp 1607101874
transform 1 0 340 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1607101874
transform 1 0 348 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_314
timestamp 1607101874
transform 1 0 356 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_315
timestamp 1607101874
transform -1 0 420 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1016
timestamp 1607101874
transform 1 0 420 0 1 2705
box -2 -3 98 103
use AOI21X1  AOI21X1_145
timestamp 1607101874
transform 1 0 516 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_229
timestamp 1607101874
transform 1 0 548 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_288
timestamp 1607101874
transform -1 0 604 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_345
timestamp 1607101874
transform -1 0 636 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_460
timestamp 1607101874
transform 1 0 636 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_336
timestamp 1607101874
transform -1 0 692 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_661
timestamp 1607101874
transform -1 0 724 0 1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_31
timestamp 1607101874
transform 1 0 724 0 1 2705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_1012
timestamp 1607101874
transform 1 0 764 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_1_0
timestamp 1607101874
transform 1 0 860 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1607101874
transform 1 0 868 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_299
timestamp 1607101874
transform 1 0 876 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_298
timestamp 1607101874
transform 1 0 908 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_895
timestamp 1607101874
transform 1 0 940 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_527
timestamp 1607101874
transform 1 0 972 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1514
timestamp 1607101874
transform 1 0 1068 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1013
timestamp 1607101874
transform 1 0 1100 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1490
timestamp 1607101874
transform 1 0 1132 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_495
timestamp 1607101874
transform 1 0 1164 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_505
timestamp 1607101874
transform 1 0 1260 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_2_0
timestamp 1607101874
transform 1 0 1356 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1607101874
transform 1 0 1364 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_303
timestamp 1607101874
transform 1 0 1372 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_302
timestamp 1607101874
transform -1 0 1436 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1502
timestamp 1607101874
transform 1 0 1436 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1501
timestamp 1607101874
transform -1 0 1500 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_484
timestamp 1607101874
transform 1 0 1500 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_222
timestamp 1607101874
transform 1 0 1524 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1254
timestamp 1607101874
transform 1 0 1548 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1010
timestamp 1607101874
transform 1 0 1580 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1253
timestamp 1607101874
transform 1 0 1676 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_155
timestamp 1607101874
transform -1 0 1740 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_185
timestamp 1607101874
transform -1 0 1764 0 1 2705
box -2 -3 26 103
use OAI22X1  OAI22X1_92
timestamp 1607101874
transform 1 0 1764 0 1 2705
box -2 -3 42 103
use BUFX4  BUFX4_366
timestamp 1607101874
transform 1 0 1804 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_605
timestamp 1607101874
transform 1 0 1836 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_3_0
timestamp 1607101874
transform -1 0 1876 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1607101874
transform -1 0 1884 0 1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_717
timestamp 1607101874
transform -1 0 1908 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_501
timestamp 1607101874
transform 1 0 1908 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_834
timestamp 1607101874
transform 1 0 2004 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_290
timestamp 1607101874
transform -1 0 2060 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_390
timestamp 1607101874
transform 1 0 2060 0 1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_219
timestamp 1607101874
transform -1 0 2140 0 1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_833
timestamp 1607101874
transform 1 0 2140 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1607101874
transform -1 0 2196 0 1 2705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_68
timestamp 1607101874
transform -1 0 2268 0 1 2705
box -2 -3 74 103
use OAI21X1  OAI21X1_706
timestamp 1607101874
transform 1 0 2268 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_760
timestamp 1607101874
transform 1 0 2300 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_4_0
timestamp 1607101874
transform 1 0 2396 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1607101874
transform 1 0 2404 0 1 2705
box -2 -3 10 103
use BUFX4  BUFX4_63
timestamp 1607101874
transform 1 0 2412 0 1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_43
timestamp 1607101874
transform -1 0 2492 0 1 2705
box -2 -3 50 103
use NOR2X1  NOR2X1_446
timestamp 1607101874
transform -1 0 2516 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_829
timestamp 1607101874
transform -1 0 2548 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_53
timestamp 1607101874
transform -1 0 2564 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_828
timestamp 1607101874
transform -1 0 2596 0 1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_277
timestamp 1607101874
transform 1 0 2596 0 1 2705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1607101874
transform 1 0 2644 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_346
timestamp 1607101874
transform 1 0 2740 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_915
timestamp 1607101874
transform -1 0 2788 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_255
timestamp 1607101874
transform 1 0 2788 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1607101874
transform -1 0 2844 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_118
timestamp 1607101874
transform -1 0 2876 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_104
timestamp 1607101874
transform -1 0 2908 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1607101874
transform -1 0 2916 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1607101874
transform -1 0 2924 0 1 2705
box -2 -3 10 103
use AOI22X1  AOI22X1_12
timestamp 1607101874
transform -1 0 2964 0 1 2705
box -2 -3 42 103
use BUFX4  BUFX4_91
timestamp 1607101874
transform 1 0 2964 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_75
timestamp 1607101874
transform 1 0 2996 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_116
timestamp 1607101874
transform -1 0 3060 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_100
timestamp 1607101874
transform 1 0 3060 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_105
timestamp 1607101874
transform 1 0 3092 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_117
timestamp 1607101874
transform -1 0 3156 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_390
timestamp 1607101874
transform -1 0 3180 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_285
timestamp 1607101874
transform -1 0 3204 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_270
timestamp 1607101874
transform 1 0 3204 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_112
timestamp 1607101874
transform 1 0 3228 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_83
timestamp 1607101874
transform 1 0 3260 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_20
timestamp 1607101874
transform -1 0 3364 0 1 2705
box -2 -3 74 103
use FILL  FILL_27_6_0
timestamp 1607101874
transform 1 0 3364 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1607101874
transform 1 0 3372 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_809
timestamp 1607101874
transform 1 0 3380 0 1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_113
timestamp 1607101874
transform -1 0 3500 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_64
timestamp 1607101874
transform -1 0 3532 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_792
timestamp 1607101874
transform 1 0 3532 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_85
timestamp 1607101874
transform 1 0 3628 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_805
timestamp 1607101874
transform -1 0 3740 0 1 2705
box -2 -3 98 103
use BUFX4  BUFX4_201
timestamp 1607101874
transform -1 0 3772 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_203
timestamp 1607101874
transform -1 0 3804 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_6
timestamp 1607101874
transform 1 0 3804 0 1 2705
box -2 -3 74 103
use OAI21X1  OAI21X1_139
timestamp 1607101874
transform 1 0 3876 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_7_0
timestamp 1607101874
transform -1 0 3916 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_7_1
timestamp 1607101874
transform -1 0 3924 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_138
timestamp 1607101874
transform -1 0 3956 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_60
timestamp 1607101874
transform 1 0 3956 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_871
timestamp 1607101874
transform 1 0 3988 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_261
timestamp 1607101874
transform -1 0 4044 0 1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_224
timestamp 1607101874
transform -1 0 4092 0 1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_870
timestamp 1607101874
transform -1 0 4124 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_431
timestamp 1607101874
transform -1 0 4156 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_432
timestamp 1607101874
transform -1 0 4188 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_338
timestamp 1607101874
transform -1 0 4204 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_1028
timestamp 1607101874
transform -1 0 4236 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1029
timestamp 1607101874
transform -1 0 4268 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_423
timestamp 1607101874
transform 1 0 4268 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_424
timestamp 1607101874
transform -1 0 4332 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1607101874
transform -1 0 4428 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_8_0
timestamp 1607101874
transform -1 0 4436 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_8_1
timestamp 1607101874
transform -1 0 4444 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_336
timestamp 1607101874
transform -1 0 4540 0 1 2705
box -2 -3 98 103
use MUX2X1  MUX2X1_178
timestamp 1607101874
transform -1 0 4588 0 1 2705
box -2 -3 50 103
use NAND2X1  NAND2X1_196
timestamp 1607101874
transform 1 0 4588 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_201
timestamp 1607101874
transform 1 0 4612 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_570
timestamp 1607101874
transform 1 0 4644 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_571
timestamp 1607101874
transform 1 0 4676 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1607101874
transform 1 0 4708 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_336
timestamp 1607101874
transform 1 0 4740 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_66
timestamp 1607101874
transform -1 0 4796 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_686
timestamp 1607101874
transform -1 0 4892 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_911
timestamp 1607101874
transform -1 0 4924 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_271
timestamp 1607101874
transform 1 0 4924 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_9_0
timestamp 1607101874
transform 1 0 4948 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_9_1
timestamp 1607101874
transform 1 0 4956 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_63
timestamp 1607101874
transform 1 0 4964 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_64
timestamp 1607101874
transform -1 0 5028 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_433
timestamp 1607101874
transform 1 0 5028 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_434
timestamp 1607101874
transform -1 0 5092 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1607101874
transform -1 0 5188 0 1 2705
box -2 -3 98 103
use AOI21X1  AOI21X1_545
timestamp 1607101874
transform 1 0 5188 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_35
timestamp 1607101874
transform -1 0 5236 0 1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_657
timestamp 1607101874
transform 1 0 5236 0 1 2705
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1607101874
transform 1 0 5260 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_409
timestamp 1607101874
transform 1 0 5284 0 1 2705
box -2 -3 18 103
use FILL  FILL_28_1
timestamp 1607101874
transform 1 0 5300 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1045
timestamp 1607101874
transform 1 0 4 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_390
timestamp 1607101874
transform -1 0 148 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_392
timestamp 1607101874
transform -1 0 196 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_1518
timestamp 1607101874
transform 1 0 196 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1517
timestamp 1607101874
transform -1 0 260 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_325
timestamp 1607101874
transform 1 0 260 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_324
timestamp 1607101874
transform -1 0 324 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_408
timestamp 1607101874
transform 1 0 324 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_0_0
timestamp 1607101874
transform 1 0 340 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1607101874
transform 1 0 348 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_385
timestamp 1607101874
transform 1 0 356 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_1080
timestamp 1607101874
transform 1 0 372 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1003
timestamp 1607101874
transform 1 0 404 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_289
timestamp 1607101874
transform -1 0 532 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_383
timestamp 1607101874
transform 1 0 532 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_660
timestamp 1607101874
transform -1 0 588 0 -1 2905
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1607101874
transform -1 0 628 0 -1 2905
box -2 -3 42 103
use AOI21X1  AOI21X1_140
timestamp 1607101874
transform 1 0 628 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_223
timestamp 1607101874
transform 1 0 660 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_515
timestamp 1607101874
transform 1 0 684 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1073
timestamp 1607101874
transform 1 0 708 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_894
timestamp 1607101874
transform 1 0 740 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1048
timestamp 1607101874
transform 1 0 772 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_1_0
timestamp 1607101874
transform 1 0 868 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1607101874
transform 1 0 876 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_615
timestamp 1607101874
transform 1 0 884 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_727
timestamp 1607101874
transform -1 0 940 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_432
timestamp 1607101874
transform 1 0 940 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_604
timestamp 1607101874
transform 1 0 964 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_716
timestamp 1607101874
transform -1 0 1020 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_433
timestamp 1607101874
transform -1 0 1044 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_785
timestamp 1607101874
transform 1 0 1044 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_391
timestamp 1607101874
transform 1 0 1076 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1525
timestamp 1607101874
transform 1 0 1100 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1526
timestamp 1607101874
transform -1 0 1164 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_537
timestamp 1607101874
transform 1 0 1164 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_288
timestamp 1607101874
transform -1 0 1284 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_967
timestamp 1607101874
transform -1 0 1316 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_2_0
timestamp 1607101874
transform 1 0 1316 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1607101874
transform 1 0 1324 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1014
timestamp 1607101874
transform 1 0 1332 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_499
timestamp 1607101874
transform 1 0 1428 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_237
timestamp 1607101874
transform -1 0 1572 0 -1 2905
box -2 -3 50 103
use INVX1  INVX1_219
timestamp 1607101874
transform -1 0 1588 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_756
timestamp 1607101874
transform 1 0 1588 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_66
timestamp 1607101874
transform 1 0 1684 0 -1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_56
timestamp 1607101874
transform -1 0 1748 0 -1 2905
box -2 -3 50 103
use AOI21X1  AOI21X1_41
timestamp 1607101874
transform 1 0 1748 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_80
timestamp 1607101874
transform -1 0 1804 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_727
timestamp 1607101874
transform 1 0 1804 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_3_0
timestamp 1607101874
transform 1 0 1900 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1607101874
transform 1 0 1908 0 -1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_407
timestamp 1607101874
transform 1 0 1916 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_723
timestamp 1607101874
transform 1 0 1940 0 -1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_40
timestamp 1607101874
transform 1 0 2036 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_78
timestamp 1607101874
transform -1 0 2092 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_252
timestamp 1607101874
transform -1 0 2116 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_836
timestamp 1607101874
transform -1 0 2148 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_739
timestamp 1607101874
transform 1 0 2148 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_772
timestamp 1607101874
transform -1 0 2276 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_70
timestamp 1607101874
transform 1 0 2276 0 -1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_60
timestamp 1607101874
transform -1 0 2340 0 -1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_251
timestamp 1607101874
transform -1 0 2364 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_4_0
timestamp 1607101874
transform -1 0 2372 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1607101874
transform -1 0 2380 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_768
timestamp 1607101874
transform -1 0 2476 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1607101874
transform -1 0 2572 0 -1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_639
timestamp 1607101874
transform 1 0 2572 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_527
timestamp 1607101874
transform -1 0 2628 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_388
timestamp 1607101874
transform 1 0 2628 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_348
timestamp 1607101874
transform 1 0 2724 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_916
timestamp 1607101874
transform 1 0 2740 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_917
timestamp 1607101874
transform -1 0 2804 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_471
timestamp 1607101874
transform 1 0 2804 0 -1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_283
timestamp 1607101874
transform 1 0 2828 0 -1 2905
box -2 -3 50 103
use INVX1  INVX1_347
timestamp 1607101874
transform -1 0 2892 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_5_0
timestamp 1607101874
transform -1 0 2900 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1607101874
transform -1 0 2908 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_380
timestamp 1607101874
transform -1 0 3004 0 -1 2905
box -2 -3 98 103
use INVX8  INVX8_6
timestamp 1607101874
transform 1 0 3004 0 -1 2905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1607101874
transform 1 0 3044 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_292
timestamp 1607101874
transform 1 0 3140 0 -1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_295
timestamp 1607101874
transform -1 0 3204 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_113
timestamp 1607101874
transform 1 0 3204 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_725
timestamp 1607101874
transform 1 0 3236 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_63
timestamp 1607101874
transform 1 0 3268 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_112
timestamp 1607101874
transform -1 0 3324 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_253
timestamp 1607101874
transform -1 0 3348 0 -1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_208
timestamp 1607101874
transform -1 0 3396 0 -1 2905
box -2 -3 50 103
use FILL  FILL_28_6_0
timestamp 1607101874
transform 1 0 3396 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1607101874
transform 1 0 3404 0 -1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_209
timestamp 1607101874
transform 1 0 3412 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_111
timestamp 1607101874
transform -1 0 3492 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_106
timestamp 1607101874
transform 1 0 3492 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_840
timestamp 1607101874
transform -1 0 3556 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_369
timestamp 1607101874
transform -1 0 3588 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_75
timestamp 1607101874
transform -1 0 3636 0 -1 2905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_788
timestamp 1607101874
transform -1 0 3732 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_82
timestamp 1607101874
transform 1 0 3732 0 -1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_72
timestamp 1607101874
transform -1 0 3796 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_200
timestamp 1607101874
transform -1 0 3828 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_205
timestamp 1607101874
transform -1 0 3860 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1607101874
transform 1 0 3860 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_7_0
timestamp 1607101874
transform 1 0 3956 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_7_1
timestamp 1607101874
transform 1 0 3964 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_185
timestamp 1607101874
transform 1 0 3972 0 -1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_171
timestamp 1607101874
transform -1 0 4036 0 -1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_260
timestamp 1607101874
transform -1 0 4060 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1607101874
transform -1 0 4156 0 -1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_198
timestamp 1607101874
transform -1 0 4188 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1607101874
transform -1 0 4284 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_69
timestamp 1607101874
transform -1 0 4332 0 -1 2905
box -2 -3 50 103
use INVX1  INVX1_79
timestamp 1607101874
transform -1 0 4348 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_781
timestamp 1607101874
transform -1 0 4444 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_8_0
timestamp 1607101874
transform -1 0 4452 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_8_1
timestamp 1607101874
transform -1 0 4460 0 -1 2905
box -2 -3 10 103
use AND2X2  AND2X2_46
timestamp 1607101874
transform -1 0 4492 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_233
timestamp 1607101874
transform 1 0 4492 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_448
timestamp 1607101874
transform -1 0 4540 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_296
timestamp 1607101874
transform -1 0 4564 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_199
timestamp 1607101874
transform -1 0 4596 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1607101874
transform -1 0 4692 0 -1 2905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_99
timestamp 1607101874
transform 1 0 4692 0 -1 2905
box -2 -3 74 103
use OAI21X1  OAI21X1_992
timestamp 1607101874
transform 1 0 4764 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_240
timestamp 1607101874
transform -1 0 4844 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_989
timestamp 1607101874
transform 1 0 4844 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_297
timestamp 1607101874
transform -1 0 4900 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_462
timestamp 1607101874
transform 1 0 4900 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_9_0
timestamp 1607101874
transform 1 0 4932 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_9_1
timestamp 1607101874
transform 1 0 4940 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_988
timestamp 1607101874
transform 1 0 4948 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_685
timestamp 1607101874
transform -1 0 5076 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_427
timestamp 1607101874
transform 1 0 5076 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1607101874
transform -1 0 5204 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_677
timestamp 1607101874
transform 1 0 5204 0 -1 2905
box -2 -3 98 103
use FILL  FILL_29_1
timestamp 1607101874
transform -1 0 5308 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_540
timestamp 1607101874
transform -1 0 100 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_325
timestamp 1607101874
transform 1 0 100 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_529
timestamp 1607101874
transform 1 0 116 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_508
timestamp 1607101874
transform 1 0 212 0 1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_608
timestamp 1607101874
transform 1 0 308 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_0_0
timestamp 1607101874
transform -1 0 348 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1607101874
transform -1 0 356 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_720
timestamp 1607101874
transform -1 0 380 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_460
timestamp 1607101874
transform 1 0 380 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1007
timestamp 1607101874
transform 1 0 412 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1009
timestamp 1607101874
transform 1 0 508 0 1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_142
timestamp 1607101874
transform 1 0 604 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_225
timestamp 1607101874
transform -1 0 660 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_516
timestamp 1607101874
transform 1 0 660 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_157
timestamp 1607101874
transform 1 0 684 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_451
timestamp 1607101874
transform 1 0 716 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_247
timestamp 1607101874
transform -1 0 772 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_192
timestamp 1607101874
transform -1 0 804 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_1_0
timestamp 1607101874
transform 1 0 804 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1607101874
transform 1 0 812 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_533
timestamp 1607101874
transform 1 0 820 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_72
timestamp 1607101874
transform -1 0 948 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_500
timestamp 1607101874
transform 1 0 948 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_176
timestamp 1607101874
transform -1 0 1076 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_186
timestamp 1607101874
transform -1 0 1100 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_446
timestamp 1607101874
transform -1 0 1116 0 1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_276
timestamp 1607101874
transform -1 0 1164 0 1 2905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1607101874
transform 1 0 1164 0 1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_737
timestamp 1607101874
transform 1 0 1260 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_323
timestamp 1607101874
transform -1 0 1324 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_386
timestamp 1607101874
transform 1 0 1324 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_968
timestamp 1607101874
transform -1 0 1372 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_2_0
timestamp 1607101874
transform 1 0 1372 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1607101874
transform 1 0 1380 0 1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_603
timestamp 1607101874
transform 1 0 1388 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_715
timestamp 1607101874
transform -1 0 1444 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_132
timestamp 1607101874
transform -1 0 1476 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_757
timestamp 1607101874
transform 1 0 1476 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_67
timestamp 1607101874
transform 1 0 1572 0 1 2905
box -2 -3 18 103
use BUFX4  BUFX4_135
timestamp 1607101874
transform 1 0 1588 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1479
timestamp 1607101874
transform 1 0 1620 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1480
timestamp 1607101874
transform -1 0 1684 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_486
timestamp 1607101874
transform -1 0 1780 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_181
timestamp 1607101874
transform 1 0 1780 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_498
timestamp 1607101874
transform 1 0 1812 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_3_0
timestamp 1607101874
transform 1 0 1836 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1607101874
transform 1 0 1844 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_748
timestamp 1607101874
transform 1 0 1852 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_134
timestamp 1607101874
transform -1 0 1980 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_62
timestamp 1607101874
transform 1 0 1980 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_835
timestamp 1607101874
transform 1 0 1996 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_364
timestamp 1607101874
transform 1 0 2028 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_363
timestamp 1607101874
transform -1 0 2092 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1607101874
transform -1 0 2108 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_776
timestamp 1607101874
transform -1 0 2204 0 1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_64
timestamp 1607101874
transform -1 0 2252 0 1 2905
box -2 -3 50 103
use BUFX4  BUFX4_144
timestamp 1607101874
transform 1 0 2252 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_93
timestamp 1607101874
transform 1 0 2284 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_49
timestamp 1607101874
transform -1 0 2340 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_280
timestamp 1607101874
transform 1 0 2340 0 1 2905
box -2 -3 50 103
use FILL  FILL_29_4_0
timestamp 1607101874
transform 1 0 2388 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1607101874
transform 1 0 2396 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_98
timestamp 1607101874
transform 1 0 2404 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_53
timestamp 1607101874
transform -1 0 2460 0 1 2905
box -2 -3 34 103
use INVX8  INVX8_31
timestamp 1607101874
transform -1 0 2500 0 1 2905
box -2 -3 42 103
use AOI21X1  AOI21X1_365
timestamp 1607101874
transform 1 0 2500 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_21
timestamp 1607101874
transform 1 0 2532 0 1 2905
box -2 -3 42 103
use MUX2X1  MUX2X1_281
timestamp 1607101874
transform 1 0 2572 0 1 2905
box -2 -3 50 103
use AOI21X1  AOI21X1_394
timestamp 1607101874
transform -1 0 2652 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_638
timestamp 1607101874
transform -1 0 2676 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_526
timestamp 1607101874
transform -1 0 2708 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1607101874
transform -1 0 2804 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1607101874
transform 1 0 2804 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_5_0
timestamp 1607101874
transform 1 0 2900 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1607101874
transform 1 0 2908 0 1 2905
box -2 -3 10 103
use INVX1  INVX1_227
timestamp 1607101874
transform 1 0 2916 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_174
timestamp 1607101874
transform 1 0 2932 0 1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_177
timestamp 1607101874
transform -1 0 3004 0 1 2905
box -2 -3 50 103
use BUFX4  BUFX4_85
timestamp 1607101874
transform -1 0 3036 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_114
timestamp 1607101874
transform -1 0 3068 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_115
timestamp 1607101874
transform 1 0 3068 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1607101874
transform 1 0 3100 0 1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_535
timestamp 1607101874
transform 1 0 3196 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_647
timestamp 1607101874
transform 1 0 3228 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_229
timestamp 1607101874
transform -1 0 3276 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_808
timestamp 1607101874
transform 1 0 3276 0 1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_564
timestamp 1607101874
transform 1 0 3372 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_6_0
timestamp 1607101874
transform 1 0 3404 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1607101874
transform 1 0 3412 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_173
timestamp 1607101874
transform 1 0 3420 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_93
timestamp 1607101874
transform -1 0 3476 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_102
timestamp 1607101874
transform 1 0 3476 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_108
timestamp 1607101874
transform -1 0 3540 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_82
timestamp 1607101874
transform -1 0 3572 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_182
timestamp 1607101874
transform 1 0 3572 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_777
timestamp 1607101874
transform 1 0 3604 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_75
timestamp 1607101874
transform 1 0 3700 0 1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_65
timestamp 1607101874
transform -1 0 3764 0 1 2905
box -2 -3 50 103
use BUFX4  BUFX4_204
timestamp 1607101874
transform 1 0 3764 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_206
timestamp 1607101874
transform 1 0 3796 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_793
timestamp 1607101874
transform 1 0 3828 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_7_0
timestamp 1607101874
transform 1 0 3924 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_7_1
timestamp 1607101874
transform 1 0 3932 0 1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_57
timestamp 1607101874
transform 1 0 3940 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_104
timestamp 1607101874
transform 1 0 3972 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_202
timestamp 1607101874
transform -1 0 4028 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_312
timestamp 1607101874
transform 1 0 4028 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_207
timestamp 1607101874
transform -1 0 4084 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1607101874
transform -1 0 4108 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_295
timestamp 1607101874
transform -1 0 4132 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_129
timestamp 1607101874
transform 1 0 4132 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_130
timestamp 1607101874
transform -1 0 4196 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_311
timestamp 1607101874
transform -1 0 4220 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_785
timestamp 1607101874
transform -1 0 4316 0 1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_609
timestamp 1607101874
transform 1 0 4316 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1048
timestamp 1607101874
transform -1 0 4372 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1044
timestamp 1607101874
transform -1 0 4404 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1045
timestamp 1607101874
transform 1 0 4404 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_8_0
timestamp 1607101874
transform -1 0 4444 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_8_1
timestamp 1607101874
transform -1 0 4452 0 1 2905
box -2 -3 10 103
use BUFX4  BUFX4_461
timestamp 1607101874
transform -1 0 4484 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1043
timestamp 1607101874
transform -1 0 4516 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_172
timestamp 1607101874
transform 1 0 4516 0 1 2905
box -2 -3 50 103
use INVX1  INVX1_186
timestamp 1607101874
transform -1 0 4580 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1607101874
transform -1 0 4676 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_401
timestamp 1607101874
transform -1 0 4692 0 1 2905
box -2 -3 18 103
use BUFX4  BUFX4_464
timestamp 1607101874
transform 1 0 4692 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_681
timestamp 1607101874
transform 1 0 4724 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_39
timestamp 1607101874
transform 1 0 4820 0 1 2905
box -2 -3 18 103
use MUX2X1  MUX2X1_31
timestamp 1607101874
transform 1 0 4836 0 1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_425
timestamp 1607101874
transform 1 0 4884 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_426
timestamp 1607101874
transform -1 0 4948 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_9_0
timestamp 1607101874
transform -1 0 4956 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_9_1
timestamp 1607101874
transform -1 0 4964 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_296
timestamp 1607101874
transform -1 0 4988 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1607101874
transform -1 0 5084 0 1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_317
timestamp 1607101874
transform 1 0 5084 0 1 2905
box -2 -3 50 103
use NOR2X1  NOR2X1_47
timestamp 1607101874
transform 1 0 5132 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1607101874
transform -1 0 5188 0 1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_51
timestamp 1607101874
transform -1 0 5260 0 1 2905
box -2 -3 74 103
use INVX1  INVX1_181
timestamp 1607101874
transform -1 0 5276 0 1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_512
timestamp 1607101874
transform -1 0 5308 0 1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_60
timestamp 1607101874
transform 1 0 4 0 -1 3105
box -2 -3 74 103
use AOI21X1  AOI21X1_158
timestamp 1607101874
transform 1 0 76 0 -1 3105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_67
timestamp 1607101874
transform 1 0 4 0 1 3105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1049
timestamp 1607101874
transform 1 0 76 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_248
timestamp 1607101874
transform -1 0 132 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_429
timestamp 1607101874
transform -1 0 164 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1607101874
transform 1 0 164 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_228
timestamp 1607101874
transform -1 0 220 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1015
timestamp 1607101874
transform 1 0 172 0 1 3105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_18
timestamp 1607101874
transform 1 0 220 0 -1 3105
box -2 -3 74 103
use AOI21X1  AOI21X1_141
timestamp 1607101874
transform 1 0 292 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_319
timestamp 1607101874
transform -1 0 300 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_0_0
timestamp 1607101874
transform 1 0 300 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_224
timestamp 1607101874
transform -1 0 348 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_0_0
timestamp 1607101874
transform 1 0 348 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1607101874
transform 1 0 356 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1017
timestamp 1607101874
transform 1 0 364 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_0_1
timestamp 1607101874
transform 1 0 308 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1008
timestamp 1607101874
transform 1 0 316 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_507
timestamp 1607101874
transform 1 0 460 0 -1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_146
timestamp 1607101874
transform 1 0 412 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_230
timestamp 1607101874
transform -1 0 468 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_987
timestamp 1607101874
transform 1 0 468 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_719
timestamp 1607101874
transform -1 0 580 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_607
timestamp 1607101874
transform -1 0 612 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_384
timestamp 1607101874
transform 1 0 564 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_265
timestamp 1607101874
transform 1 0 588 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_118
timestamp 1607101874
transform -1 0 636 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_66
timestamp 1607101874
transform -1 0 668 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_811
timestamp 1607101874
transform 1 0 668 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_264
timestamp 1607101874
transform -1 0 652 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_380
timestamp 1607101874
transform -1 0 684 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_331
timestamp 1607101874
transform 1 0 684 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_617
timestamp 1607101874
transform 1 0 764 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_729
timestamp 1607101874
transform -1 0 820 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_374
timestamp 1607101874
transform 1 0 716 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1475
timestamp 1607101874
transform -1 0 780 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1476
timestamp 1607101874
transform -1 0 812 0 1 3105
box -2 -3 34 103
use FILL  FILL_30_1_0
timestamp 1607101874
transform 1 0 820 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_1
timestamp 1607101874
transform 1 0 828 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_541
timestamp 1607101874
transform 1 0 836 0 -1 3105
box -2 -3 98 103
use BUFX4  BUFX4_445
timestamp 1607101874
transform -1 0 844 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_1_0
timestamp 1607101874
transform 1 0 844 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1_1
timestamp 1607101874
transform 1 0 852 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_1465
timestamp 1607101874
transform 1 0 860 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1466
timestamp 1607101874
transform 1 0 892 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1018
timestamp 1607101874
transform 1 0 932 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_479
timestamp 1607101874
transform 1 0 924 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_995
timestamp 1607101874
transform 1 0 1028 0 -1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_147
timestamp 1607101874
transform 1 0 1020 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_231
timestamp 1607101874
transform -1 0 1076 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_252
timestamp 1607101874
transform 1 0 1076 0 1 3105
box -2 -3 18 103
use INVX1  INVX1_284
timestamp 1607101874
transform 1 0 1092 0 1 3105
box -2 -3 18 103
use INVX8  INVX8_24
timestamp 1607101874
transform -1 0 1148 0 1 3105
box -2 -3 42 103
use INVX1  INVX1_135
timestamp 1607101874
transform 1 0 1124 0 -1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_122
timestamp 1607101874
transform -1 0 1188 0 -1 3105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_485
timestamp 1607101874
transform 1 0 1188 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_72
timestamp 1607101874
transform -1 0 1172 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_74
timestamp 1607101874
transform 1 0 1172 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_272
timestamp 1607101874
transform 1 0 1196 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_622
timestamp 1607101874
transform 1 0 1284 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_289
timestamp 1607101874
transform -1 0 1332 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_273
timestamp 1607101874
transform -1 0 1260 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_991
timestamp 1607101874
transform 1 0 1260 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_671
timestamp 1607101874
transform 1 0 1332 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_2_0
timestamp 1607101874
transform 1 0 1364 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_1
timestamp 1607101874
transform 1 0 1372 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_1478
timestamp 1607101874
transform 1 0 1380 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_942
timestamp 1607101874
transform 1 0 1412 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_2_0
timestamp 1607101874
transform 1 0 1356 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_1
timestamp 1607101874
transform 1 0 1364 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_672
timestamp 1607101874
transform 1 0 1372 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_670
timestamp 1607101874
transform 1 0 1404 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1477
timestamp 1607101874
transform -1 0 1476 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_374
timestamp 1607101874
transform 1 0 1476 0 -1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_57
timestamp 1607101874
transform -1 0 1540 0 -1 3105
box -2 -3 50 103
use AOI21X1  AOI21X1_304
timestamp 1607101874
transform 1 0 1436 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1012
timestamp 1607101874
transform 1 0 1468 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_142
timestamp 1607101874
transform 1 0 1500 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_479
timestamp 1607101874
transform 1 0 1540 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_945
timestamp 1607101874
transform 1 0 1564 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1473
timestamp 1607101874
transform 1 0 1596 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_434
timestamp 1607101874
transform -1 0 1564 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1481
timestamp 1607101874
transform 1 0 1564 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1482
timestamp 1607101874
transform -1 0 1628 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_487
timestamp 1607101874
transform 1 0 1628 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1474
timestamp 1607101874
transform 1 0 1660 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_273
timestamp 1607101874
transform 1 0 1692 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1159
timestamp 1607101874
transform 1 0 1628 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_593
timestamp 1607101874
transform 1 0 1660 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_491
timestamp 1607101874
transform -1 0 1788 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_483
timestamp 1607101874
transform -1 0 1820 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_905
timestamp 1607101874
transform -1 0 1852 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_480
timestamp 1607101874
transform 1 0 1788 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_721
timestamp 1607101874
transform 1 0 1812 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_951
timestamp 1607101874
transform 1 0 1852 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_414
timestamp 1607101874
transform 1 0 1900 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_3_0
timestamp 1607101874
transform 1 0 1908 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_1
timestamp 1607101874
transform 1 0 1916 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_996
timestamp 1607101874
transform -1 0 2028 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_51
timestamp 1607101874
transform 1 0 1924 0 1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_41
timestamp 1607101874
transform -1 0 1988 0 1 3105
box -2 -3 50 103
use AOI21X1  AOI21X1_435
timestamp 1607101874
transform 1 0 1988 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_152
timestamp 1607101874
transform -1 0 2052 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_219
timestamp 1607101874
transform 1 0 2028 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_138
timestamp 1607101874
transform -1 0 2084 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_52
timestamp 1607101874
transform -1 0 2132 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_1031
timestamp 1607101874
transform 1 0 2052 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_590
timestamp 1607101874
transform 1 0 2084 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_749
timestamp 1607101874
transform 1 0 2108 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_324
timestamp 1607101874
transform 1 0 2132 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_738
timestamp 1607101874
transform -1 0 2196 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_302
timestamp 1607101874
transform -1 0 2212 0 -1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_387
timestamp 1607101874
transform -1 0 2308 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_63
timestamp 1607101874
transform 1 0 2204 0 1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_53
timestamp 1607101874
transform -1 0 2268 0 1 3105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_379
timestamp 1607101874
transform -1 0 2404 0 -1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_443
timestamp 1607101874
transform 1 0 2268 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_442
timestamp 1607101874
transform 1 0 2300 0 1 3105
box -2 -3 34 103
use FILL  FILL_30_4_0
timestamp 1607101874
transform 1 0 2404 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_1
timestamp 1607101874
transform 1 0 2412 0 -1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_529
timestamp 1607101874
transform 1 0 2420 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1030
timestamp 1607101874
transform 1 0 2332 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_4_0
timestamp 1607101874
transform 1 0 2364 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_4_1
timestamp 1607101874
transform 1 0 2372 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_494
timestamp 1607101874
transform 1 0 2380 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_641
timestamp 1607101874
transform 1 0 2452 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_462
timestamp 1607101874
transform -1 0 2508 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1607101874
transform 1 0 2508 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1488
timestamp 1607101874
transform -1 0 2508 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1487
timestamp 1607101874
transform -1 0 2540 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1607101874
transform -1 0 2564 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1160
timestamp 1607101874
transform -1 0 2596 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_380
timestamp 1607101874
transform 1 0 2596 0 -1 3105
box -2 -3 50 103
use NAND2X1  NAND2X1_41
timestamp 1607101874
transform -1 0 2564 0 1 3105
box -2 -3 26 103
use AND2X2  AND2X2_52
timestamp 1607101874
transform 1 0 2564 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1161
timestamp 1607101874
transform 1 0 2596 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1486
timestamp 1607101874
transform 1 0 2628 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_432
timestamp 1607101874
transform -1 0 2660 0 -1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_490
timestamp 1607101874
transform -1 0 2756 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1485
timestamp 1607101874
transform 1 0 2660 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_493
timestamp 1607101874
transform 1 0 2692 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_38
timestamp 1607101874
transform 1 0 2756 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_953
timestamp 1607101874
transform -1 0 2812 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_952
timestamp 1607101874
transform -1 0 2844 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_41
timestamp 1607101874
transform 1 0 2788 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_212
timestamp 1607101874
transform -1 0 2844 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_926
timestamp 1607101874
transform -1 0 2908 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_401
timestamp 1607101874
transform 1 0 2844 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_280
timestamp 1607101874
transform 1 0 2924 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_5_1
timestamp 1607101874
transform 1 0 2916 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_5_0
timestamp 1607101874
transform 1 0 2908 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_375
timestamp 1607101874
transform -1 0 2924 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_5_1
timestamp 1607101874
transform -1 0 2908 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_0
timestamp 1607101874
transform -1 0 2900 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_489
timestamp 1607101874
transform -1 0 3020 0 -1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_379
timestamp 1607101874
transform 1 0 2844 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_563
timestamp 1607101874
transform 1 0 3020 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_695
timestamp 1607101874
transform 1 0 2956 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_583
timestamp 1607101874
transform -1 0 3012 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1607101874
transform -1 0 3108 0 1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_290
timestamp 1607101874
transform -1 0 3100 0 -1 3105
box -2 -3 50 103
use INVX8  INVX8_29
timestamp 1607101874
transform -1 0 3140 0 -1 3105
box -2 -3 42 103
use NAND2X1  NAND2X1_172
timestamp 1607101874
transform 1 0 3108 0 1 3105
box -2 -3 26 103
use AND2X2  AND2X2_26
timestamp 1607101874
transform 1 0 3132 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_430
timestamp 1607101874
transform 1 0 3140 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_421
timestamp 1607101874
transform 1 0 3172 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1607101874
transform -1 0 3300 0 -1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_235
timestamp 1607101874
transform 1 0 3164 0 1 3105
box -2 -3 50 103
use MUX2X1  MUX2X1_302
timestamp 1607101874
transform 1 0 3212 0 1 3105
box -2 -3 50 103
use INVX1  INVX1_228
timestamp 1607101874
transform 1 0 3300 0 -1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_294
timestamp 1607101874
transform -1 0 3364 0 -1 3105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_363
timestamp 1607101874
transform 1 0 3260 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_838
timestamp 1607101874
transform -1 0 3396 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_6_0
timestamp 1607101874
transform 1 0 3396 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_6_1
timestamp 1607101874
transform 1 0 3404 0 -1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_367
timestamp 1607101874
transform 1 0 3412 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_293
timestamp 1607101874
transform 1 0 3356 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_318
timestamp 1607101874
transform 1 0 3372 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_6_0
timestamp 1607101874
transform 1 0 3404 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_6_1
timestamp 1607101874
transform 1 0 3412 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_727
timestamp 1607101874
transform 1 0 3420 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_842
timestamp 1607101874
transform 1 0 3444 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1607101874
transform -1 0 3572 0 -1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_562
timestamp 1607101874
transform 1 0 3452 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_353
timestamp 1607101874
transform -1 0 3508 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_99
timestamp 1607101874
transform -1 0 3532 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_54
timestamp 1607101874
transform -1 0 3564 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_646
timestamp 1607101874
transform 1 0 3572 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_534
timestamp 1607101874
transform -1 0 3628 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_841
timestamp 1607101874
transform -1 0 3660 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_769
timestamp 1607101874
transform 1 0 3564 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_334
timestamp 1607101874
transform -1 0 3676 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_1035
timestamp 1607101874
transform 1 0 3676 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1034
timestamp 1607101874
transform 1 0 3708 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_444
timestamp 1607101874
transform 1 0 3740 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1032
timestamp 1607101874
transform 1 0 3660 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_502
timestamp 1607101874
transform -1 0 3716 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_501
timestamp 1607101874
transform 1 0 3716 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_87
timestamp 1607101874
transform -1 0 3756 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_804
timestamp 1607101874
transform 1 0 3772 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_796
timestamp 1607101874
transform -1 0 3852 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_136
timestamp 1607101874
transform -1 0 3900 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1607101874
transform -1 0 3932 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_7_0
timestamp 1607101874
transform -1 0 3940 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_7_1
timestamp 1607101874
transform -1 0 3948 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_726
timestamp 1607101874
transform -1 0 3884 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_414
timestamp 1607101874
transform 1 0 3884 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_413
timestamp 1607101874
transform -1 0 3932 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_7_0
timestamp 1607101874
transform -1 0 3940 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_7_1
timestamp 1607101874
transform -1 0 3948 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_1033
timestamp 1607101874
transform -1 0 3980 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_106
timestamp 1607101874
transform 1 0 3980 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_874
timestamp 1607101874
transform -1 0 4036 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_773
timestamp 1607101874
transform -1 0 4132 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_367
timestamp 1607101874
transform -1 0 4044 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_71
timestamp 1607101874
transform 1 0 4132 0 -1 3105
box -2 -3 18 103
use INVX1  INVX1_450
timestamp 1607101874
transform 1 0 4044 0 1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_298
timestamp 1607101874
transform -1 0 4108 0 1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_1105
timestamp 1607101874
transform -1 0 4140 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_312
timestamp 1607101874
transform 1 0 4140 0 1 3105
box -2 -3 50 103
use MUX2X1  MUX2X1_61
timestamp 1607101874
transform -1 0 4196 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_632
timestamp 1607101874
transform 1 0 4196 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_396
timestamp 1607101874
transform -1 0 4260 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_418
timestamp 1607101874
transform -1 0 4204 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_353
timestamp 1607101874
transform -1 0 4300 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1332
timestamp 1607101874
transform 1 0 4260 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1333
timestamp 1607101874
transform -1 0 4324 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_334
timestamp 1607101874
transform 1 0 4324 0 -1 3105
box -2 -3 98 103
use BUFX4  BUFX4_397
timestamp 1607101874
transform 1 0 4300 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_320
timestamp 1607101874
transform 1 0 4332 0 1 3105
box -2 -3 26 103
use FILL  FILL_30_8_0
timestamp 1607101874
transform 1 0 4420 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_8_1
timestamp 1607101874
transform 1 0 4428 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_470
timestamp 1607101874
transform 1 0 4436 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1046
timestamp 1607101874
transform -1 0 4388 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_449
timestamp 1607101874
transform -1 0 4420 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_508
timestamp 1607101874
transform 1 0 4420 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_8_0
timestamp 1607101874
transform 1 0 4444 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_1151
timestamp 1607101874
transform -1 0 4500 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1607101874
transform -1 0 4524 0 -1 3105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_55
timestamp 1607101874
transform 1 0 4524 0 -1 3105
box -2 -3 74 103
use FILL  FILL_31_8_1
timestamp 1607101874
transform 1 0 4452 0 1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_368
timestamp 1607101874
transform 1 0 4460 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_839
timestamp 1607101874
transform -1 0 4524 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_127
timestamp 1607101874
transform 1 0 4524 0 1 3105
box -2 -3 34 103
use OAI22X1  OAI22X1_6
timestamp 1607101874
transform 1 0 4596 0 -1 3105
box -2 -3 42 103
use NOR2X1  NOR2X1_375
timestamp 1607101874
transform -1 0 4660 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_128
timestamp 1607101874
transform -1 0 4588 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_784
timestamp 1607101874
transform -1 0 4684 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1607101874
transform -1 0 4756 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_402
timestamp 1607101874
transform -1 0 4700 0 1 3105
box -2 -3 18 103
use BUFX4  BUFX4_358
timestamp 1607101874
transform -1 0 4732 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_409
timestamp 1607101874
transform -1 0 4764 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_410
timestamp 1607101874
transform -1 0 4788 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_655
timestamp 1607101874
transform -1 0 4884 0 -1 3105
box -2 -3 98 103
use BUFX4  BUFX4_339
timestamp 1607101874
transform 1 0 4764 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_569
timestamp 1607101874
transform 1 0 4796 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_417
timestamp 1607101874
transform 1 0 4828 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1607101874
transform -1 0 4916 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1607101874
transform -1 0 4948 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_9_0
timestamp 1607101874
transform 1 0 4948 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_418
timestamp 1607101874
transform -1 0 4892 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1607101874
transform -1 0 4988 0 1 3105
box -2 -3 98 103
use FILL  FILL_30_9_1
timestamp 1607101874
transform 1 0 4956 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_53
timestamp 1607101874
transform 1 0 4964 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_672
timestamp 1607101874
transform -1 0 5092 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_9_0
timestamp 1607101874
transform 1 0 4988 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_9_1
timestamp 1607101874
transform 1 0 4996 0 1 3105
box -2 -3 10 103
use MUX2X1  MUX2X1_68
timestamp 1607101874
transform 1 0 5004 0 1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_631
timestamp 1607101874
transform -1 0 5084 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_344
timestamp 1607101874
transform -1 0 5188 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1197
timestamp 1607101874
transform -1 0 5116 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_315
timestamp 1607101874
transform 1 0 5116 0 1 3105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_802
timestamp 1607101874
transform 1 0 5188 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_232
timestamp 1607101874
transform -1 0 5180 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_61
timestamp 1607101874
transform 1 0 5180 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_342
timestamp 1607101874
transform 1 0 5212 0 1 3105
box -2 -3 98 103
use FILL  FILL_31_1
timestamp 1607101874
transform -1 0 5292 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_2
timestamp 1607101874
transform -1 0 5300 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_3
timestamp 1607101874
transform -1 0 5308 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1607101874
transform -1 0 100 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_301
timestamp 1607101874
transform 1 0 100 0 -1 3305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_89
timestamp 1607101874
transform 1 0 116 0 -1 3305
box -2 -3 74 103
use OAI21X1  OAI21X1_143
timestamp 1607101874
transform -1 0 220 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_92
timestamp 1607101874
transform -1 0 236 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_813
timestamp 1607101874
transform -1 0 332 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_0_0
timestamp 1607101874
transform 1 0 332 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1607101874
transform 1 0 340 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_412
timestamp 1607101874
transform 1 0 348 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_340
timestamp 1607101874
transform -1 0 476 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_319
timestamp 1607101874
transform -1 0 492 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_484
timestamp 1607101874
transform -1 0 588 0 -1 3305
box -2 -3 98 103
use BUFX4  BUFX4_452
timestamp 1607101874
transform -1 0 620 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1402
timestamp 1607101874
transform -1 0 652 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1403
timestamp 1607101874
transform -1 0 684 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_204
timestamp 1607101874
transform 1 0 684 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_205
timestamp 1607101874
transform -1 0 748 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_889
timestamp 1607101874
transform 1 0 748 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_1_0
timestamp 1607101874
transform 1 0 844 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1607101874
transform 1 0 852 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_431
timestamp 1607101874
transform 1 0 860 0 -1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_245
timestamp 1607101874
transform -1 0 924 0 -1 3305
box -2 -3 50 103
use BUFX4  BUFX4_162
timestamp 1607101874
transform -1 0 956 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_328
timestamp 1607101874
transform 1 0 956 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_370
timestamp 1607101874
transform 1 0 1052 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1341
timestamp 1607101874
transform 1 0 1068 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_231
timestamp 1607101874
transform -1 0 1148 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_1470
timestamp 1607101874
transform 1 0 1148 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_481
timestamp 1607101874
transform 1 0 1180 0 -1 3305
box -2 -3 98 103
use BUFX4  BUFX4_160
timestamp 1607101874
transform 1 0 1276 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1469
timestamp 1607101874
transform -1 0 1340 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_2_0
timestamp 1607101874
transform 1 0 1340 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1607101874
transform 1 0 1348 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_992
timestamp 1607101874
transform 1 0 1356 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_274
timestamp 1607101874
transform -1 0 1484 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_275
timestamp 1607101874
transform -1 0 1516 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_904
timestamp 1607101874
transform -1 0 1548 0 -1 3305
box -2 -3 34 103
use OAI22X1  OAI22X1_35
timestamp 1607101874
transform -1 0 1588 0 -1 3305
box -2 -3 42 103
use NAND2X1  NAND2X1_60
timestamp 1607101874
transform 1 0 1588 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_487
timestamp 1607101874
transform 1 0 1612 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_253
timestamp 1607101874
transform 1 0 1708 0 -1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_378
timestamp 1607101874
transform -1 0 1772 0 -1 3305
box -2 -3 50 103
use AND2X2  AND2X2_23
timestamp 1607101874
transform 1 0 1772 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_595
timestamp 1607101874
transform -1 0 1836 0 -1 3305
box -2 -3 34 103
use INVX8  INVX8_7
timestamp 1607101874
transform -1 0 1876 0 -1 3305
box -2 -3 42 103
use FILL  FILL_32_3_0
timestamp 1607101874
transform 1 0 1876 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1607101874
transform 1 0 1884 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_594
timestamp 1607101874
transform 1 0 1892 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_752
timestamp 1607101874
transform 1 0 1924 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_333
timestamp 1607101874
transform -1 0 2036 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_112
timestamp 1607101874
transform 1 0 2036 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1607101874
transform -1 0 2100 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1607101874
transform 1 0 2100 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_764
timestamp 1607101874
transform -1 0 2228 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_120
timestamp 1607101874
transform -1 0 2260 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1607101874
transform 1 0 2260 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_113
timestamp 1607101874
transform 1 0 2292 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_753
timestamp 1607101874
transform -1 0 2420 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_4_0
timestamp 1607101874
transform 1 0 2420 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1607101874
transform 1 0 2428 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_906
timestamp 1607101874
transform 1 0 2436 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1085
timestamp 1607101874
transform 1 0 2468 0 -1 3305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_54
timestamp 1607101874
transform -1 0 2572 0 -1 3305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_13
timestamp 1607101874
transform -1 0 2644 0 -1 3305
box -2 -3 74 103
use NOR2X1  NOR2X1_180
timestamp 1607101874
transform 1 0 2644 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_402
timestamp 1607101874
transform 1 0 2668 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_40
timestamp 1607101874
transform 1 0 2700 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_464
timestamp 1607101874
transform -1 0 2756 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_258
timestamp 1607101874
transform 1 0 2756 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_931
timestamp 1607101874
transform 1 0 2804 0 -1 3305
box -2 -3 34 103
use OAI22X1  OAI22X1_38
timestamp 1607101874
transform -1 0 2876 0 -1 3305
box -2 -3 42 103
use FILL  FILL_32_5_0
timestamp 1607101874
transform 1 0 2876 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1607101874
transform 1 0 2884 0 -1 3305
box -2 -3 10 103
use MUX2X1  MUX2X1_181
timestamp 1607101874
transform 1 0 2892 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_928
timestamp 1607101874
transform -1 0 2972 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1607101874
transform -1 0 2996 0 -1 3305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_65
timestamp 1607101874
transform -1 0 3068 0 -1 3305
box -2 -3 74 103
use BUFX4  BUFX4_449
timestamp 1607101874
transform 1 0 3068 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_927
timestamp 1607101874
transform -1 0 3132 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1607101874
transform 1 0 3132 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_539
timestamp 1607101874
transform 1 0 3228 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_651
timestamp 1607101874
transform -1 0 3284 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_371
timestamp 1607101874
transform -1 0 3380 0 -1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_412
timestamp 1607101874
transform -1 0 3404 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_6_0
timestamp 1607101874
transform -1 0 3412 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_6_1
timestamp 1607101874
transform -1 0 3420 0 -1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_96
timestamp 1607101874
transform -1 0 3444 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_533
timestamp 1607101874
transform 1 0 3444 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1607101874
transform 1 0 3476 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_765
timestamp 1607101874
transform 1 0 3572 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_122
timestamp 1607101874
transform 1 0 3668 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1607101874
transform -1 0 3732 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_366
timestamp 1607101874
transform 1 0 3732 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_77
timestamp 1607101874
transform -1 0 3812 0 -1 3305
box -2 -3 50 103
use BUFX4  BUFX4_316
timestamp 1607101874
transform 1 0 3812 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1607101874
transform 1 0 3844 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1316
timestamp 1607101874
transform 1 0 3876 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_7_0
timestamp 1607101874
transform -1 0 3916 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_7_1
timestamp 1607101874
transform -1 0 3924 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_375
timestamp 1607101874
transform -1 0 4020 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1317
timestamp 1607101874
transform -1 0 4052 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_654
timestamp 1607101874
transform -1 0 4084 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_798
timestamp 1607101874
transform 1 0 4084 0 -1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_581
timestamp 1607101874
transform -1 0 4204 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_89
timestamp 1607101874
transform 1 0 4204 0 -1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_79
timestamp 1607101874
transform -1 0 4268 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_1199
timestamp 1607101874
transform -1 0 4300 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1329
timestamp 1607101874
transform 1 0 4300 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1330
timestamp 1607101874
transform -1 0 4364 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_357
timestamp 1607101874
transform -1 0 4460 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_8_0
timestamp 1607101874
transform -1 0 4468 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_8_1
timestamp 1607101874
transform -1 0 4476 0 -1 3305
box -2 -3 10 103
use OAI22X1  OAI22X1_71
timestamp 1607101874
transform -1 0 4516 0 -1 3305
box -2 -3 42 103
use NAND2X1  NAND2X1_26
timestamp 1607101874
transform 1 0 4516 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1607101874
transform 1 0 4540 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_135
timestamp 1607101874
transform -1 0 4604 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_803
timestamp 1607101874
transform -1 0 4700 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_783
timestamp 1607101874
transform 1 0 4700 0 -1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_298
timestamp 1607101874
transform 1 0 4796 0 -1 3305
box -2 -3 26 103
use BUFX4  BUFX4_58
timestamp 1607101874
transform -1 0 4852 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_653
timestamp 1607101874
transform -1 0 4884 0 -1 3305
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1607101874
transform 1 0 4884 0 -1 3305
box -2 -3 42 103
use NOR2X1  NOR2X1_379
timestamp 1607101874
transform -1 0 4948 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_9_0
timestamp 1607101874
transform -1 0 4956 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_9_1
timestamp 1607101874
transform -1 0 4964 0 -1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_582
timestamp 1607101874
transform -1 0 4988 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_78
timestamp 1607101874
transform -1 0 5004 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_780
timestamp 1607101874
transform -1 0 5100 0 -1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_114
timestamp 1607101874
transform 1 0 5100 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_65
timestamp 1607101874
transform -1 0 5156 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_376
timestamp 1607101874
transform -1 0 5180 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_40
timestamp 1607101874
transform 1 0 5180 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_667
timestamp 1607101874
transform -1 0 5300 0 -1 3305
box -2 -3 98 103
use FILL  FILL_33_1
timestamp 1607101874
transform -1 0 5308 0 -1 3305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_74
timestamp 1607101874
transform 1 0 4 0 1 3305
box -2 -3 74 103
use OAI21X1  OAI21X1_1289
timestamp 1607101874
transform -1 0 108 0 1 3305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_7
timestamp 1607101874
transform 1 0 108 0 1 3305
box -2 -3 74 103
use NAND2X1  NAND2X1_356
timestamp 1607101874
transform 1 0 180 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_50
timestamp 1607101874
transform -1 0 228 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_989
timestamp 1607101874
transform 1 0 228 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_0_0
timestamp 1607101874
transform 1 0 324 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_0_1
timestamp 1607101874
transform 1 0 332 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_269
timestamp 1607101874
transform 1 0 340 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_268
timestamp 1607101874
transform -1 0 404 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_482
timestamp 1607101874
transform 1 0 404 0 1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_579
timestamp 1607101874
transform 1 0 500 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_691
timestamp 1607101874
transform 1 0 532 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1471
timestamp 1607101874
transform -1 0 588 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1607101874
transform 1 0 588 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_470
timestamp 1607101874
transform 1 0 620 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1607101874
transform 1 0 644 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_163
timestamp 1607101874
transform -1 0 764 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_905
timestamp 1607101874
transform 1 0 764 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_1_0
timestamp 1607101874
transform 1 0 860 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_1_1
timestamp 1607101874
transform 1 0 868 0 1 3305
box -2 -3 10 103
use AOI21X1  AOI21X1_101
timestamp 1607101874
transform 1 0 876 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_166
timestamp 1607101874
transform 1 0 908 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_164
timestamp 1607101874
transform -1 0 964 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_267
timestamp 1607101874
transform 1 0 964 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_266
timestamp 1607101874
transform 1 0 996 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_988
timestamp 1607101874
transform 1 0 1028 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_357
timestamp 1607101874
transform -1 0 1148 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_405
timestamp 1607101874
transform 1 0 1148 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_999
timestamp 1607101874
transform 1 0 1164 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_281
timestamp 1607101874
transform 1 0 1260 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_280
timestamp 1607101874
transform -1 0 1324 0 1 3305
box -2 -3 34 103
use AND2X2  AND2X2_25
timestamp 1607101874
transform 1 0 1324 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_2_0
timestamp 1607101874
transform 1 0 1356 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_2_1
timestamp 1607101874
transform 1 0 1364 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_994
timestamp 1607101874
transform 1 0 1372 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_279
timestamp 1607101874
transform 1 0 1468 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_278
timestamp 1607101874
transform -1 0 1532 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_286
timestamp 1607101874
transform -1 0 1564 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_469
timestamp 1607101874
transform 1 0 1564 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_163
timestamp 1607101874
transform 1 0 1588 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_276
timestamp 1607101874
transform 1 0 1620 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1607101874
transform -1 0 1684 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_993
timestamp 1607101874
transform 1 0 1684 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1065
timestamp 1607101874
transform 1 0 1780 0 1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_455
timestamp 1607101874
transform 1 0 1812 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_3_0
timestamp 1607101874
transform 1 0 1844 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_3_1
timestamp 1607101874
transform 1 0 1852 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_717
timestamp 1607101874
transform 1 0 1860 0 1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_39
timestamp 1607101874
transform 1 0 1956 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_76
timestamp 1607101874
transform -1 0 2012 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_376
timestamp 1607101874
transform 1 0 2012 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1017
timestamp 1607101874
transform 1 0 2044 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_345
timestamp 1607101874
transform -1 0 2108 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_79
timestamp 1607101874
transform -1 0 2140 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_314
timestamp 1607101874
transform -1 0 2164 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_161
timestamp 1607101874
transform 1 0 2164 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_761
timestamp 1607101874
transform -1 0 2292 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_94
timestamp 1607101874
transform 1 0 2292 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_50
timestamp 1607101874
transform -1 0 2348 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_4_0
timestamp 1607101874
transform 1 0 2348 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_4_1
timestamp 1607101874
transform 1 0 2356 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_389
timestamp 1607101874
transform 1 0 2364 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_410
timestamp 1607101874
transform 1 0 2460 0 1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_282
timestamp 1607101874
transform 1 0 2476 0 1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_268
timestamp 1607101874
transform 1 0 2524 0 1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_588
timestamp 1607101874
transform 1 0 2620 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_700
timestamp 1607101874
transform -1 0 2676 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_929
timestamp 1607101874
transform -1 0 2708 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_355
timestamp 1607101874
transform 1 0 2708 0 1 3305
box -2 -3 50 103
use INVX1  INVX1_358
timestamp 1607101874
transform -1 0 2772 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1607101874
transform 1 0 2772 0 1 3305
box -2 -3 98 103
use AND2X2  AND2X2_40
timestamp 1607101874
transform -1 0 2900 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_5_0
timestamp 1607101874
transform 1 0 2900 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_5_1
timestamp 1607101874
transform 1 0 2908 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1607101874
transform 1 0 2916 0 1 3305
box -2 -3 98 103
use AND2X2  AND2X2_39
timestamp 1607101874
transform -1 0 3044 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_347
timestamp 1607101874
transform 1 0 3044 0 1 3305
box -2 -3 50 103
use INVX1  INVX1_356
timestamp 1607101874
transform -1 0 3108 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1607101874
transform -1 0 3204 0 1 3305
box -2 -3 98 103
use INVX8  INVX8_17
timestamp 1607101874
transform 1 0 3204 0 1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_1307
timestamp 1607101874
transform 1 0 3244 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1607101874
transform 1 0 3276 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_324
timestamp 1607101874
transform -1 0 3340 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1306
timestamp 1607101874
transform -1 0 3372 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_6_0
timestamp 1607101874
transform 1 0 3372 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_6_1
timestamp 1607101874
transform 1 0 3380 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1607101874
transform 1 0 3388 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_448
timestamp 1607101874
transform 1 0 3484 0 1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_293
timestamp 1607101874
transform -1 0 3548 0 1 3305
box -2 -3 50 103
use NOR2X1  NOR2X1_645
timestamp 1607101874
transform -1 0 3572 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1099
timestamp 1607101874
transform -1 0 3604 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_527
timestamp 1607101874
transform -1 0 3628 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_52
timestamp 1607101874
transform -1 0 3660 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_528
timestamp 1607101874
transform 1 0 3660 0 1 3305
box -2 -3 26 103
use OAI22X1  OAI22X1_51
timestamp 1607101874
transform 1 0 3684 0 1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_1098
timestamp 1607101874
transform -1 0 3756 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_837
timestamp 1607101874
transform 1 0 3756 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_318
timestamp 1607101874
transform 1 0 3788 0 1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_1338
timestamp 1607101874
transform 1 0 3836 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1339
timestamp 1607101874
transform -1 0 3900 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1312
timestamp 1607101874
transform -1 0 3932 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_7_0
timestamp 1607101874
transform -1 0 3940 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_7_1
timestamp 1607101874
transform -1 0 3948 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_1313
timestamp 1607101874
transform -1 0 3980 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1607101874
transform -1 0 4076 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_27
timestamp 1607101874
transform -1 0 4100 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_471
timestamp 1607101874
transform 1 0 4100 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_26
timestamp 1607101874
transform 1 0 4132 0 1 3305
box -2 -3 50 103
use INVX1  INVX1_34
timestamp 1607101874
transform -1 0 4196 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_663
timestamp 1607101874
transform -1 0 4292 0 1 3305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_58
timestamp 1607101874
transform -1 0 4364 0 1 3305
box -2 -3 74 103
use OAI21X1  OAI21X1_132
timestamp 1607101874
transform 1 0 4364 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1607101874
transform 1 0 4396 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_8_0
timestamp 1607101874
transform -1 0 4436 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_8_1
timestamp 1607101874
transform -1 0 4444 0 1 3305
box -2 -3 10 103
use INVX8  INVX8_10
timestamp 1607101874
transform -1 0 4484 0 1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_1198
timestamp 1607101874
transform -1 0 4516 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1607101874
transform -1 0 4548 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_141
timestamp 1607101874
transform -1 0 4580 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1607101874
transform 1 0 4580 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_126
timestamp 1607101874
transform -1 0 4644 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_719
timestamp 1607101874
transform 1 0 4644 0 1 3305
box -2 -3 34 103
use OAI22X1  OAI22X1_19
timestamp 1607101874
transform -1 0 4716 0 1 3305
box -2 -3 42 103
use NOR2X1  NOR2X1_409
timestamp 1607101874
transform -1 0 4740 0 1 3305
box -2 -3 26 103
use MUX2X1  MUX2X1_67
timestamp 1607101874
transform 1 0 4740 0 1 3305
box -2 -3 50 103
use INVX1  INVX1_77
timestamp 1607101874
transform -1 0 4804 0 1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_410
timestamp 1607101874
transform -1 0 4828 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_103
timestamp 1607101874
transform -1 0 4852 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_56
timestamp 1607101874
transform -1 0 4884 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_791
timestamp 1607101874
transform -1 0 4980 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_9_0
timestamp 1607101874
transform -1 0 4988 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_9_1
timestamp 1607101874
transform -1 0 4996 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_810
timestamp 1607101874
transform -1 0 5092 0 1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_76
timestamp 1607101874
transform 1 0 5092 0 1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_795
timestamp 1607101874
transform -1 0 5236 0 1 3305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_77
timestamp 1607101874
transform -1 0 5308 0 1 3305
box -2 -3 74 103
use BUFX4  BUFX4_4
timestamp 1607101874
transform 1 0 4 0 -1 3505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_44
timestamp 1607101874
transform 1 0 36 0 -1 3505
box -2 -3 74 103
use NAND2X1  NAND2X1_353
timestamp 1607101874
transform -1 0 132 0 -1 3505
box -2 -3 26 103
use INVX8  INVX8_3
timestamp 1607101874
transform -1 0 172 0 -1 3505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_480
timestamp 1607101874
transform 1 0 172 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1468
timestamp 1607101874
transform -1 0 300 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1467
timestamp 1607101874
transform -1 0 332 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_0_0
timestamp 1607101874
transform 1 0 332 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_0_1
timestamp 1607101874
transform 1 0 340 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_492
timestamp 1607101874
transform 1 0 348 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1472
timestamp 1607101874
transform 1 0 444 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_778
timestamp 1607101874
transform -1 0 508 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1484
timestamp 1607101874
transform 1 0 508 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1483
timestamp 1607101874
transform -1 0 572 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_431
timestamp 1607101874
transform 1 0 572 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1000
timestamp 1607101874
transform -1 0 692 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_283
timestamp 1607101874
transform -1 0 724 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_878
timestamp 1607101874
transform 1 0 724 0 -1 3505
box -2 -3 98 103
use NOR2X1  NOR2X1_153
timestamp 1607101874
transform 1 0 820 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_1_0
timestamp 1607101874
transform 1 0 844 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_1_1
timestamp 1607101874
transform 1 0 852 0 -1 3505
box -2 -3 10 103
use BUFX4  BUFX4_335
timestamp 1607101874
transform 1 0 860 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_447
timestamp 1607101874
transform 1 0 892 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_270
timestamp 1607101874
transform 1 0 916 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_271
timestamp 1607101874
transform -1 0 980 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_990
timestamp 1607101874
transform 1 0 980 0 -1 3505
box -2 -3 98 103
use BUFX4  BUFX4_174
timestamp 1607101874
transform 1 0 1076 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_893
timestamp 1607101874
transform 1 0 1108 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_212
timestamp 1607101874
transform 1 0 1204 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_213
timestamp 1607101874
transform -1 0 1268 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_846
timestamp 1607101874
transform 1 0 1268 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1607101874
transform 1 0 1300 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_2_0
timestamp 1607101874
transform 1 0 1396 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_2_1
timestamp 1607101874
transform 1 0 1404 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1002
timestamp 1607101874
transform 1 0 1412 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_287
timestamp 1607101874
transform 1 0 1508 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1607101874
transform -1 0 1564 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_285
timestamp 1607101874
transform -1 0 1596 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_615
timestamp 1607101874
transform 1 0 1596 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1001
timestamp 1607101874
transform 1 0 1620 0 -1 3505
box -2 -3 98 103
use AND2X2  AND2X2_47
timestamp 1607101874
transform 1 0 1716 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1607101874
transform 1 0 1748 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1067
timestamp 1607101874
transform 1 0 1772 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_246
timestamp 1607101874
transform -1 0 1852 0 -1 3505
box -2 -3 50 103
use AOI21X1  AOI21X1_111
timestamp 1607101874
transform 1 0 1852 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_181
timestamp 1607101874
transform 1 0 1900 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_935
timestamp 1607101874
transform 1 0 1924 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_221
timestamp 1607101874
transform 1 0 2020 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_937
timestamp 1607101874
transform 1 0 2044 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_65
timestamp 1607101874
transform -1 0 2164 0 -1 3505
box -2 -3 26 103
use MUX2X1  MUX2X1_107
timestamp 1607101874
transform -1 0 2212 0 -1 3505
box -2 -3 50 103
use INVX1  INVX1_120
timestamp 1607101874
transform -1 0 2228 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_929
timestamp 1607101874
transform -1 0 2324 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_66
timestamp 1607101874
transform 1 0 2324 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_64
timestamp 1607101874
transform 1 0 2348 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_118
timestamp 1607101874
transform -1 0 2388 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_4_0
timestamp 1607101874
transform -1 0 2396 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_4_1
timestamp 1607101874
transform -1 0 2404 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_925
timestamp 1607101874
transform -1 0 2500 0 -1 3505
box -2 -3 98 103
use NOR2X1  NOR2X1_169
timestamp 1607101874
transform -1 0 2524 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1607101874
transform 1 0 2524 0 -1 3505
box -2 -3 98 103
use INVX1  INVX1_359
timestamp 1607101874
transform 1 0 2620 0 -1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_352
timestamp 1607101874
transform -1 0 2684 0 -1 3505
box -2 -3 50 103
use OAI21X1  OAI21X1_930
timestamp 1607101874
transform 1 0 2684 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1607101874
transform 1 0 2716 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1435
timestamp 1607101874
transform 1 0 2812 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1434
timestamp 1607101874
transform -1 0 2876 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1426
timestamp 1607101874
transform 1 0 2876 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_5_0
timestamp 1607101874
transform -1 0 2916 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_5_1
timestamp 1607101874
transform -1 0 2924 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1427
timestamp 1607101874
transform -1 0 2956 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_349
timestamp 1607101874
transform -1 0 3004 0 -1 3505
box -2 -3 50 103
use INVX1  INVX1_308
timestamp 1607101874
transform -1 0 3020 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1607101874
transform -1 0 3116 0 -1 3505
box -2 -3 98 103
use BUFX4  BUFX4_66
timestamp 1607101874
transform -1 0 3148 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_328
timestamp 1607101874
transform -1 0 3172 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_53
timestamp 1607101874
transform -1 0 3204 0 -1 3505
box -2 -3 34 103
use OAI22X1  OAI22X1_36
timestamp 1607101874
transform -1 0 3244 0 -1 3505
box -2 -3 42 103
use MUX2X1  MUX2X1_291
timestamp 1607101874
transform 1 0 3244 0 -1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1607101874
transform 1 0 3292 0 -1 3505
box -2 -3 98 103
use INVX1  INVX1_291
timestamp 1607101874
transform 1 0 3388 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_6_0
timestamp 1607101874
transform 1 0 3404 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_6_1
timestamp 1607101874
transform 1 0 3412 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_724
timestamp 1607101874
transform 1 0 3420 0 -1 3505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_22
timestamp 1607101874
transform -1 0 3524 0 -1 3505
box -2 -3 74 103
use NAND2X1  NAND2X1_68
timestamp 1607101874
transform -1 0 3548 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_468
timestamp 1607101874
transform 1 0 3548 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_70
timestamp 1607101874
transform 1 0 3572 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_537
timestamp 1607101874
transform 1 0 3596 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_649
timestamp 1607101874
transform -1 0 3652 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1607101874
transform -1 0 3748 0 -1 3505
box -2 -3 98 103
use BUFX4  BUFX4_37
timestamp 1607101874
transform 1 0 3748 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1607101874
transform 1 0 3780 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_133
timestamp 1607101874
transform -1 0 3836 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_90
timestamp 1607101874
transform -1 0 3852 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_453
timestamp 1607101874
transform -1 0 3868 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_337
timestamp 1607101874
transform 1 0 3868 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_7_0
timestamp 1607101874
transform -1 0 3972 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_7_1
timestamp 1607101874
transform -1 0 3980 0 -1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_529
timestamp 1607101874
transform -1 0 4004 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_371
timestamp 1607101874
transform 1 0 4004 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_542
timestamp 1607101874
transform 1 0 4036 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_654
timestamp 1607101874
transform -1 0 4092 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_349
timestamp 1607101874
transform -1 0 4188 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_333
timestamp 1607101874
transform 1 0 4188 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1106
timestamp 1607101874
transform -1 0 4244 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1607101874
transform 1 0 4244 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_105
timestamp 1607101874
transform -1 0 4300 0 -1 3505
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1607101874
transform 1 0 4300 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_470
timestamp 1607101874
transform 1 0 4324 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_786
timestamp 1607101874
transform 1 0 4356 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_8_0
timestamp 1607101874
transform 1 0 4452 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_8_1
timestamp 1607101874
transform 1 0 4460 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1189
timestamp 1607101874
transform 1 0 4468 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_806
timestamp 1607101874
transform -1 0 4596 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_717
timestamp 1607101874
transform -1 0 4628 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_212
timestamp 1607101874
transform -1 0 4660 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_226
timestamp 1607101874
transform 1 0 4660 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_720
timestamp 1607101874
transform -1 0 4716 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_790
timestamp 1607101874
transform -1 0 4812 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_779
timestamp 1607101874
transform -1 0 4908 0 -1 3505
box -2 -3 98 103
use BUFX4  BUFX4_460
timestamp 1607101874
transform 1 0 4908 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_9_0
timestamp 1607101874
transform -1 0 4948 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_9_1
timestamp 1607101874
transform -1 0 4956 0 -1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_380
timestamp 1607101874
transform -1 0 4980 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_406
timestamp 1607101874
transform 1 0 4980 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_405
timestamp 1607101874
transform -1 0 5044 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1607101874
transform -1 0 5140 0 -1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_166
timestamp 1607101874
transform 1 0 5140 0 -1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1607101874
transform -1 0 5284 0 -1 3505
box -2 -3 98 103
use FILL  FILL_35_1
timestamp 1607101874
transform -1 0 5292 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_2
timestamp 1607101874
transform -1 0 5300 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_3
timestamp 1607101874
transform -1 0 5308 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_997
timestamp 1607101874
transform -1 0 100 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_136
timestamp 1607101874
transform 1 0 100 0 1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_123
timestamp 1607101874
transform -1 0 164 0 1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_488
timestamp 1607101874
transform 1 0 164 0 1 3505
box -2 -3 98 103
use BUFX4  BUFX4_422
timestamp 1607101874
transform 1 0 260 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_602
timestamp 1607101874
transform 1 0 292 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_714
timestamp 1607101874
transform -1 0 348 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_0_0
timestamp 1607101874
transform 1 0 348 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_0_1
timestamp 1607101874
transform 1 0 356 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_779
timestamp 1607101874
transform 1 0 364 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_881
timestamp 1607101874
transform 1 0 396 0 1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_93
timestamp 1607101874
transform 1 0 492 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_156
timestamp 1607101874
transform -1 0 548 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_780
timestamp 1607101874
transform -1 0 580 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_247
timestamp 1607101874
transform -1 0 628 0 1 3505
box -2 -3 50 103
use INVX8  INVX8_14
timestamp 1607101874
transform -1 0 668 0 1 3505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_892
timestamp 1607101874
transform 1 0 668 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_210
timestamp 1607101874
transform 1 0 764 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_211
timestamp 1607101874
transform -1 0 828 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_448
timestamp 1607101874
transform -1 0 852 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_1_0
timestamp 1607101874
transform 1 0 852 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_1_1
timestamp 1607101874
transform 1 0 860 0 1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_152
timestamp 1607101874
transform 1 0 868 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_90
timestamp 1607101874
transform -1 0 924 0 1 3505
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1607101874
transform 1 0 924 0 1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_845
timestamp 1607101874
transform 1 0 964 0 1 3505
box -2 -3 34 103
use OAI22X1  OAI22X1_26
timestamp 1607101874
transform -1 0 1036 0 1 3505
box -2 -3 42 103
use NOR2X1  NOR2X1_585
timestamp 1607101874
transform 1 0 1036 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_900
timestamp 1607101874
transform 1 0 1060 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_255
timestamp 1607101874
transform -1 0 1180 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_219
timestamp 1607101874
transform 1 0 1180 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_218
timestamp 1607101874
transform -1 0 1244 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_887
timestamp 1607101874
transform 1 0 1244 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1411
timestamp 1607101874
transform 1 0 1340 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_2_0
timestamp 1607101874
transform -1 0 1380 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_2_1
timestamp 1607101874
transform -1 0 1388 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1410
timestamp 1607101874
transform -1 0 1420 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_201
timestamp 1607101874
transform 1 0 1420 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_281
timestamp 1607101874
transform -1 0 1476 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_218
timestamp 1607101874
transform -1 0 1500 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1246
timestamp 1607101874
transform 1 0 1500 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_616
timestamp 1607101874
transform 1 0 1532 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_284
timestamp 1607101874
transform 1 0 1556 0 1 3505
box -2 -3 34 103
use OAI22X1  OAI22X1_88
timestamp 1607101874
transform -1 0 1628 0 1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_1066
timestamp 1607101874
transform 1 0 1628 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_998
timestamp 1607101874
transform 1 0 1660 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1247
timestamp 1607101874
transform 1 0 1756 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_220
timestamp 1607101874
transform 1 0 1788 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_139
timestamp 1607101874
transform -1 0 1844 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_3_0
timestamp 1607101874
transform 1 0 1844 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_3_1
timestamp 1607101874
transform 1 0 1852 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_725
timestamp 1607101874
transform 1 0 1860 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_54
timestamp 1607101874
transform 1 0 1956 0 1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_44
timestamp 1607101874
transform -1 0 2020 0 1 3505
box -2 -3 50 103
use AOI21X1  AOI21X1_436
timestamp 1607101874
transform 1 0 2020 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_112
timestamp 1607101874
transform 1 0 2052 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_182
timestamp 1607101874
transform -1 0 2108 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1018
timestamp 1607101874
transform -1 0 2140 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_432
timestamp 1607101874
transform 1 0 2140 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_998
timestamp 1607101874
transform -1 0 2204 0 1 3505
box -2 -3 34 103
use OAI22X1  OAI22X1_43
timestamp 1607101874
transform -1 0 2244 0 1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_1000
timestamp 1607101874
transform -1 0 2276 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_999
timestamp 1607101874
transform -1 0 2308 0 1 3505
box -2 -3 34 103
use AND2X2  AND2X2_43
timestamp 1607101874
transform -1 0 2340 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_105
timestamp 1607101874
transform 1 0 2340 0 1 3505
box -2 -3 50 103
use FILL  FILL_35_4_0
timestamp 1607101874
transform 1 0 2388 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_4_1
timestamp 1607101874
transform 1 0 2396 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_909
timestamp 1607101874
transform 1 0 2404 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_112
timestamp 1607101874
transform 1 0 2500 0 1 3505
box -2 -3 18 103
use BUFX4  BUFX4_35
timestamp 1607101874
transform 1 0 2516 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_997
timestamp 1607101874
transform -1 0 2580 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_996
timestamp 1607101874
transform 1 0 2580 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1318
timestamp 1607101874
transform 1 0 2612 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1319
timestamp 1607101874
transform -1 0 2676 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_365
timestamp 1607101874
transform -1 0 2692 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_376
timestamp 1607101874
transform -1 0 2788 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1425
timestamp 1607101874
transform 1 0 2788 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1424
timestamp 1607101874
transform 1 0 2820 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_5_0
timestamp 1607101874
transform 1 0 2852 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_5_1
timestamp 1607101874
transform 1 0 2860 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1607101874
transform 1 0 2868 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1248
timestamp 1607101874
transform 1 0 2964 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_330
timestamp 1607101874
transform 1 0 2996 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_752
timestamp 1607101874
transform 1 0 3028 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_374
timestamp 1607101874
transform -1 0 3156 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1314
timestamp 1607101874
transform -1 0 3188 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1315
timestamp 1607101874
transform -1 0 3220 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_463
timestamp 1607101874
transform 1 0 3220 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_435
timestamp 1607101874
transform -1 0 3260 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_474
timestamp 1607101874
transform -1 0 3356 0 1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_374
timestamp 1607101874
transform -1 0 3404 0 1 3505
box -2 -3 50 103
use FILL  FILL_35_6_0
timestamp 1607101874
transform 1 0 3404 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_6_1
timestamp 1607101874
transform 1 0 3412 0 1 3505
box -2 -3 10 103
use AOI22X1  AOI22X1_32
timestamp 1607101874
transform 1 0 3420 0 1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_1069
timestamp 1607101874
transform -1 0 3492 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_121
timestamp 1607101874
transform 1 0 3492 0 1 3505
box -2 -3 50 103
use INVX1  INVX1_134
timestamp 1607101874
transform -1 0 3556 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_981
timestamp 1607101874
transform -1 0 3652 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_228
timestamp 1607101874
transform 1 0 3652 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_781
timestamp 1607101874
transform 1 0 3676 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_430
timestamp 1607101874
transform 1 0 3708 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_782
timestamp 1607101874
transform 1 0 3732 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_800
timestamp 1607101874
transform 1 0 3764 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_345
timestamp 1607101874
transform 1 0 3860 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_7_0
timestamp 1607101874
transform -1 0 3964 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_7_1
timestamp 1607101874
transform -1 0 3972 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1096
timestamp 1607101874
transform -1 0 4004 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1095
timestamp 1607101874
transform -1 0 4036 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1097
timestamp 1607101874
transform -1 0 4068 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_526
timestamp 1607101874
transform -1 0 4092 0 1 3505
box -2 -3 26 103
use OAI22X1  OAI22X1_52
timestamp 1607101874
transform 1 0 4092 0 1 3505
box -2 -3 42 103
use BUFX4  BUFX4_158
timestamp 1607101874
transform -1 0 4164 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_578
timestamp 1607101874
transform 1 0 4164 0 1 3505
box -2 -3 26 103
use OAI22X1  OAI22X1_72
timestamp 1607101874
transform 1 0 4188 0 1 3505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_794
timestamp 1607101874
transform 1 0 4228 0 1 3505
box -2 -3 98 103
use NOR2X1  NOR2X1_411
timestamp 1607101874
transform -1 0 4348 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1104
timestamp 1607101874
transform -1 0 4380 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_316
timestamp 1607101874
transform -1 0 4412 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_8_0
timestamp 1607101874
transform -1 0 4420 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_8_1
timestamp 1607101874
transform -1 0 4428 0 1 3505
box -2 -3 10 103
use MUX2X1  MUX2X1_308
timestamp 1607101874
transform -1 0 4476 0 1 3505
box -2 -3 50 103
use OAI21X1  OAI21X1_1191
timestamp 1607101874
transform 1 0 4476 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1190
timestamp 1607101874
transform 1 0 4508 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_718
timestamp 1607101874
transform -1 0 4572 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_497
timestamp 1607101874
transform -1 0 4604 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_315
timestamp 1607101874
transform -1 0 4636 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_70
timestamp 1607101874
transform 1 0 4636 0 1 3505
box -2 -3 50 103
use INVX1  INVX1_84
timestamp 1607101874
transform -1 0 4700 0 1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_74
timestamp 1607101874
transform -1 0 4748 0 1 3505
box -2 -3 50 103
use MUX2X1  MUX2X1_71
timestamp 1607101874
transform 1 0 4748 0 1 3505
box -2 -3 50 103
use INVX1  INVX1_81
timestamp 1607101874
transform -1 0 4812 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_787
timestamp 1607101874
transform -1 0 4908 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_652
timestamp 1607101874
transform -1 0 4940 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_9_0
timestamp 1607101874
transform -1 0 4948 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_9_1
timestamp 1607101874
transform -1 0 4956 0 1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_525
timestamp 1607101874
transform -1 0 4980 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_549
timestamp 1607101874
transform 1 0 4980 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_661
timestamp 1607101874
transform 1 0 5012 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_333
timestamp 1607101874
transform -1 0 5132 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_716
timestamp 1607101874
transform -1 0 5164 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_290
timestamp 1607101874
transform -1 0 5180 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_807
timestamp 1607101874
transform -1 0 5276 0 1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_62
timestamp 1607101874
transform 1 0 5276 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_211
timestamp 1607101874
transform 1 0 4 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_109
timestamp 1607101874
transform 1 0 36 0 -1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_304
timestamp 1607101874
transform 1 0 60 0 -1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_115
timestamp 1607101874
transform -1 0 108 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_449
timestamp 1607101874
transform 1 0 108 0 -1 3705
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1607101874
transform 1 0 140 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_207
timestamp 1607101874
transform 1 0 172 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_209
timestamp 1607101874
transform 1 0 204 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_320
timestamp 1607101874
transform -1 0 268 0 -1 3705
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1607101874
transform -1 0 308 0 -1 3705
box -2 -3 42 103
use FILL  FILL_36_0_0
timestamp 1607101874
transform 1 0 308 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_0_1
timestamp 1607101874
transform 1 0 316 0 -1 3705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_33
timestamp 1607101874
transform 1 0 324 0 -1 3705
box -2 -3 74 103
use INVX2  INVX2_15
timestamp 1607101874
transform 1 0 396 0 -1 3705
box -2 -3 18 103
use AOI21X1  AOI21X1_97
timestamp 1607101874
transform 1 0 412 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_161
timestamp 1607101874
transform -1 0 468 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_411
timestamp 1607101874
transform -1 0 564 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_310
timestamp 1607101874
transform 1 0 564 0 -1 3705
box -2 -3 18 103
use MUX2X1  MUX2X1_341
timestamp 1607101874
transform -1 0 628 0 -1 3705
box -2 -3 50 103
use AOI21X1  AOI21X1_573
timestamp 1607101874
transform 1 0 628 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_685
timestamp 1607101874
transform -1 0 684 0 -1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_232
timestamp 1607101874
transform -1 0 732 0 -1 3705
box -2 -3 50 103
use NOR2X1  NOR2X1_160
timestamp 1607101874
transform -1 0 756 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_96
timestamp 1607101874
transform -1 0 788 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_896
timestamp 1607101874
transform 1 0 788 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_1_0
timestamp 1607101874
transform -1 0 892 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_1_1
timestamp 1607101874
transform -1 0 900 0 -1 3705
box -2 -3 10 103
use BUFX4  BUFX4_405
timestamp 1607101874
transform -1 0 932 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1408
timestamp 1607101874
transform -1 0 964 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_94
timestamp 1607101874
transform 1 0 964 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_157
timestamp 1607101874
transform -1 0 1020 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_882
timestamp 1607101874
transform 1 0 1020 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_944
timestamp 1607101874
transform 1 0 1116 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1204
timestamp 1607101874
transform 1 0 1148 0 -1 3705
box -2 -3 34 103
use OAI22X1  OAI22X1_73
timestamp 1607101874
transform -1 0 1220 0 -1 3705
box -2 -3 42 103
use NOR2X1  NOR2X1_586
timestamp 1607101874
transform -1 0 1244 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_333
timestamp 1607101874
transform 1 0 1244 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_754
timestamp 1607101874
transform 1 0 1276 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_890
timestamp 1607101874
transform -1 0 1404 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_2_0
timestamp 1607101874
transform 1 0 1404 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_2_1
timestamp 1607101874
transform 1 0 1412 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_207
timestamp 1607101874
transform 1 0 1420 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_206
timestamp 1607101874
transform -1 0 1484 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_200
timestamp 1607101874
transform -1 0 1516 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_404
timestamp 1607101874
transform -1 0 1548 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_59
timestamp 1607101874
transform -1 0 1572 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_220
timestamp 1607101874
transform 1 0 1572 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_221
timestamp 1607101874
transform -1 0 1636 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_847
timestamp 1607101874
transform -1 0 1668 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_901
timestamp 1607101874
transform -1 0 1764 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_397
timestamp 1607101874
transform 1 0 1764 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_1011
timestamp 1607101874
transform 1 0 1780 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_307
timestamp 1607101874
transform 1 0 1812 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_410
timestamp 1607101874
transform -1 0 1868 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_3_0
timestamp 1607101874
transform -1 0 1876 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_3_1
timestamp 1607101874
transform -1 0 1884 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_943
timestamp 1607101874
transform -1 0 1916 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1205
timestamp 1607101874
transform -1 0 1948 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1607101874
transform -1 0 1980 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_151
timestamp 1607101874
transform -1 0 2004 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_89
timestamp 1607101874
transform -1 0 2036 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_694
timestamp 1607101874
transform -1 0 2068 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_288
timestamp 1607101874
transform -1 0 2084 0 -1 3705
box -2 -3 18 103
use AOI22X1  AOI22X1_22
timestamp 1607101874
transform 1 0 2084 0 -1 3705
box -2 -3 42 103
use AOI21X1  AOI21X1_375
timestamp 1607101874
transform 1 0 2124 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_168
timestamp 1607101874
transform -1 0 2188 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_921
timestamp 1607101874
transform 1 0 2188 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_911
timestamp 1607101874
transform 1 0 2284 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_4_0
timestamp 1607101874
transform -1 0 2388 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_4_1
timestamp 1607101874
transform -1 0 2396 0 -1 3705
box -2 -3 10 103
use NAND2X1  NAND2X1_63
timestamp 1607101874
transform -1 0 2420 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_697
timestamp 1607101874
transform -1 0 2452 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_695
timestamp 1607101874
transform 1 0 2452 0 -1 3705
box -2 -3 34 103
use OAI22X1  OAI22X1_15
timestamp 1607101874
transform -1 0 2524 0 -1 3705
box -2 -3 42 103
use OAI21X1  OAI21X1_696
timestamp 1607101874
transform -1 0 2556 0 -1 3705
box -2 -3 34 103
use AND2X2  AND2X2_42
timestamp 1607101874
transform -1 0 2588 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_99
timestamp 1607101874
transform -1 0 2636 0 -1 3705
box -2 -3 50 103
use NOR2X1  NOR2X1_398
timestamp 1607101874
transform -1 0 2660 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_937
timestamp 1607101874
transform -1 0 2692 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_565
timestamp 1607101874
transform 1 0 2692 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_367
timestamp 1607101874
transform 1 0 2724 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_566
timestamp 1607101874
transform -1 0 2780 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_581
timestamp 1607101874
transform 1 0 2780 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_693
timestamp 1607101874
transform -1 0 2836 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1163
timestamp 1607101874
transform -1 0 2868 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1164
timestamp 1607101874
transform 1 0 2868 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_5_0
timestamp 1607101874
transform 1 0 2900 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_5_1
timestamp 1607101874
transform 1 0 2908 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1162
timestamp 1607101874
transform 1 0 2916 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_332
timestamp 1607101874
transform 1 0 2948 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_331
timestamp 1607101874
transform -1 0 3012 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_751
timestamp 1607101874
transform -1 0 3044 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_343
timestamp 1607101874
transform 1 0 3044 0 -1 3705
box -2 -3 50 103
use INVX1  INVX1_307
timestamp 1607101874
transform -1 0 3108 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_407
timestamp 1607101874
transform -1 0 3204 0 -1 3705
box -2 -3 98 103
use OAI22X1  OAI22X1_91
timestamp 1607101874
transform 1 0 3204 0 -1 3705
box -2 -3 42 103
use BUFX4  BUFX4_123
timestamp 1607101874
transform -1 0 3276 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_377
timestamp 1607101874
transform -1 0 3308 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_675
timestamp 1607101874
transform -1 0 3340 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_433
timestamp 1607101874
transform -1 0 3356 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_470
timestamp 1607101874
transform -1 0 3452 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_6_0
timestamp 1607101874
transform -1 0 3460 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_6_1
timestamp 1607101874
transform -1 0 3468 0 -1 3705
box -2 -3 10 103
use MUX2X1  MUX2X1_371
timestamp 1607101874
transform -1 0 3516 0 -1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_71
timestamp 1607101874
transform 1 0 3516 0 -1 3705
box -2 -3 26 103
use AND2X2  AND2X2_48
timestamp 1607101874
transform -1 0 3572 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_166
timestamp 1607101874
transform 1 0 3572 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_457
timestamp 1607101874
transform -1 0 3636 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1070
timestamp 1607101874
transform -1 0 3668 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_975
timestamp 1607101874
transform 1 0 3668 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_305
timestamp 1607101874
transform 1 0 3764 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_901
timestamp 1607101874
transform -1 0 3828 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_673
timestamp 1607101874
transform -1 0 3860 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_754
timestamp 1607101874
transform 1 0 3860 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_7_0
timestamp 1607101874
transform 1 0 3956 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_7_1
timestamp 1607101874
transform 1 0 3964 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_116
timestamp 1607101874
transform 1 0 3972 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1607101874
transform 1 0 4004 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_343
timestamp 1607101874
transform 1 0 4036 0 -1 3705
box -2 -3 26 103
use BUFX4  BUFX4_33
timestamp 1607101874
transform 1 0 4060 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_54
timestamp 1607101874
transform 1 0 4092 0 -1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_1192
timestamp 1607101874
transform -1 0 4172 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1103
timestamp 1607101874
transform -1 0 4204 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_456
timestamp 1607101874
transform -1 0 4236 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1068
timestamp 1607101874
transform -1 0 4268 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_261
timestamp 1607101874
transform 1 0 4268 0 -1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_345
timestamp 1607101874
transform -1 0 4340 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1196
timestamp 1607101874
transform -1 0 4372 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_579
timestamp 1607101874
transform -1 0 4396 0 -1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_208
timestamp 1607101874
transform -1 0 4420 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_417
timestamp 1607101874
transform -1 0 4436 0 -1 3705
box -2 -3 18 103
use FILL  FILL_36_8_0
timestamp 1607101874
transform 1 0 4436 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_8_1
timestamp 1607101874
transform 1 0 4444 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_361
timestamp 1607101874
transform 1 0 4452 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_130
timestamp 1607101874
transform -1 0 4580 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_443
timestamp 1607101874
transform -1 0 4612 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_450
timestamp 1607101874
transform -1 0 4644 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_577
timestamp 1607101874
transform -1 0 4668 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_80
timestamp 1607101874
transform -1 0 4684 0 -1 3705
box -2 -3 18 103
use BUFX4  BUFX4_425
timestamp 1607101874
transform 1 0 4684 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_782
timestamp 1607101874
transform -1 0 4812 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_258
timestamp 1607101874
transform -1 0 4844 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_463
timestamp 1607101874
transform 1 0 4844 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_873
timestamp 1607101874
transform 1 0 4876 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_9_0
timestamp 1607101874
transform -1 0 4916 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_9_1
timestamp 1607101874
transform -1 0 4924 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1607101874
transform -1 0 5020 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_414
timestamp 1607101874
transform 1 0 5020 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_413
timestamp 1607101874
transform -1 0 5084 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1607101874
transform 1 0 5084 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_44
timestamp 1607101874
transform -1 0 5148 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_659
timestamp 1607101874
transform -1 0 5244 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_193
timestamp 1607101874
transform -1 0 5276 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_655
timestamp 1607101874
transform 1 0 5276 0 -1 3705
box -2 -3 26 103
use FILL  FILL_37_1
timestamp 1607101874
transform -1 0 5308 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_448
timestamp 1607101874
transform 1 0 4 0 1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1607101874
transform 1 0 36 0 1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_22
timestamp 1607101874
transform 1 0 68 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_460
timestamp 1607101874
transform 1 0 100 0 1 3705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_3
timestamp 1607101874
transform -1 0 204 0 1 3705
box -2 -3 74 103
use AND2X2  AND2X2_4
timestamp 1607101874
transform 1 0 204 0 1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1607101874
transform -1 0 268 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_539
timestamp 1607101874
transform 1 0 268 0 1 3705
box -2 -3 34 103
use OR2X2  OR2X2_3
timestamp 1607101874
transform 1 0 300 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_0_0
timestamp 1607101874
transform 1 0 332 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_0_1
timestamp 1607101874
transform 1 0 340 0 1 3705
box -2 -3 10 103
use NOR2X1  NOR2X1_307
timestamp 1607101874
transform 1 0 348 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_110
timestamp 1607101874
transform 1 0 372 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1607101874
transform 1 0 396 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_208
timestamp 1607101874
transform 1 0 420 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1607101874
transform 1 0 452 0 1 3705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_71
timestamp 1607101874
transform 1 0 484 0 1 3705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_897
timestamp 1607101874
transform 1 0 556 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1607101874
transform 1 0 652 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_904
timestamp 1607101874
transform 1 0 748 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_1_0
timestamp 1607101874
transform 1 0 844 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_1_1
timestamp 1607101874
transform 1 0 852 0 1 3705
box -2 -3 10 103
use AOI21X1  AOI21X1_100
timestamp 1607101874
transform 1 0 860 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1607101874
transform 1 0 892 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1409
timestamp 1607101874
transform 1 0 916 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1607101874
transform 1 0 948 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_309
timestamp 1607101874
transform 1 0 1044 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1607101874
transform 1 0 1060 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_1397
timestamp 1607101874
transform -1 0 1188 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1114
timestamp 1607101874
transform -1 0 1220 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1396
timestamp 1607101874
transform -1 0 1252 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_415
timestamp 1607101874
transform -1 0 1348 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_2_0
timestamp 1607101874
transform 1 0 1348 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_2_1
timestamp 1607101874
transform 1 0 1356 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1417
timestamp 1607101874
transform 1 0 1364 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1416
timestamp 1607101874
transform -1 0 1428 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_194
timestamp 1607101874
transform 1 0 1428 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_195
timestamp 1607101874
transform -1 0 1492 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_884
timestamp 1607101874
transform 1 0 1492 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_844
timestamp 1607101874
transform 1 0 1588 0 1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_371
timestamp 1607101874
transform -1 0 1652 0 1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_372
timestamp 1607101874
transform -1 0 1684 0 1 3705
box -2 -3 34 103
use INVX8  INVX8_21
timestamp 1607101874
transform -1 0 1724 0 1 3705
box -2 -3 42 103
use NOR2X1  NOR2X1_587
timestamp 1607101874
transform -1 0 1748 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_885
timestamp 1607101874
transform -1 0 1844 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_197
timestamp 1607101874
transform 1 0 1844 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_3_0
timestamp 1607101874
transform -1 0 1884 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_3_1
timestamp 1607101874
transform -1 0 1892 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_196
timestamp 1607101874
transform -1 0 1924 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_198
timestamp 1607101874
transform 1 0 1924 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_199
timestamp 1607101874
transform 1 0 1956 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_886
timestamp 1607101874
transform -1 0 2084 0 1 3705
box -2 -3 98 103
use OAI22X1  OAI22X1_75
timestamp 1607101874
transform 1 0 2084 0 1 3705
box -2 -3 42 103
use NOR2X1  NOR2X1_150
timestamp 1607101874
transform -1 0 2148 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_877
timestamp 1607101874
transform -1 0 2244 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_346
timestamp 1607101874
transform -1 0 2268 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_107
timestamp 1607101874
transform 1 0 2268 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_175
timestamp 1607101874
transform 1 0 2300 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_431
timestamp 1607101874
transform 1 0 2324 0 1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_310
timestamp 1607101874
transform 1 0 2356 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_4_0
timestamp 1607101874
transform -1 0 2396 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_4_1
timestamp 1607101874
transform -1 0 2404 0 1 3705
box -2 -3 10 103
use AOI21X1  AOI21X1_309
timestamp 1607101874
transform -1 0 2436 0 1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_204
timestamp 1607101874
transform -1 0 2484 0 1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_256
timestamp 1607101874
transform 1 0 2484 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_103
timestamp 1607101874
transform 1 0 2508 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_170
timestamp 1607101874
transform 1 0 2540 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_224
timestamp 1607101874
transform -1 0 2596 0 1 3705
box -2 -3 34 103
use INVX8  INVX8_22
timestamp 1607101874
transform 1 0 2596 0 1 3705
box -2 -3 42 103
use BUFX4  BUFX4_140
timestamp 1607101874
transform 1 0 2636 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_139
timestamp 1607101874
transform 1 0 2668 0 1 3705
box -2 -3 34 103
use AOI22X1  AOI22X1_20
timestamp 1607101874
transform -1 0 2740 0 1 3705
box -2 -3 42 103
use NAND2X1  NAND2X1_231
timestamp 1607101874
transform 1 0 2740 0 1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_177
timestamp 1607101874
transform -1 0 2788 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_236
timestamp 1607101874
transform 1 0 2788 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_237
timestamp 1607101874
transform -1 0 2852 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_5_0
timestamp 1607101874
transform -1 0 2860 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_5_1
timestamp 1607101874
transform -1 0 2868 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_933
timestamp 1607101874
transform -1 0 2964 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_488
timestamp 1607101874
transform -1 0 2996 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_328
timestamp 1607101874
transform -1 0 3028 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_232
timestamp 1607101874
transform -1 0 3052 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1607101874
transform -1 0 3148 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_938
timestamp 1607101874
transform 1 0 3148 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_477
timestamp 1607101874
transform -1 0 3204 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_604
timestamp 1607101874
transform 1 0 3204 0 1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_279
timestamp 1607101874
transform 1 0 3236 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_466
timestamp 1607101874
transform -1 0 3364 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_278
timestamp 1607101874
transform 1 0 3364 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_710
timestamp 1607101874
transform 1 0 3396 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_6_0
timestamp 1607101874
transform -1 0 3428 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_6_1
timestamp 1607101874
transform -1 0 3436 0 1 3705
box -2 -3 10 103
use AOI21X1  AOI21X1_598
timestamp 1607101874
transform -1 0 3468 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_603
timestamp 1607101874
transform -1 0 3500 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1607101874
transform -1 0 3524 0 1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_202
timestamp 1607101874
transform -1 0 3548 0 1 3705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_15
timestamp 1607101874
transform 1 0 3548 0 1 3705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_985
timestamp 1607101874
transform -1 0 3716 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_128
timestamp 1607101874
transform 1 0 3716 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_206
timestamp 1607101874
transform -1 0 3772 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_241
timestamp 1607101874
transform 1 0 3772 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_751
timestamp 1607101874
transform 1 0 3796 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_110
timestamp 1607101874
transform 1 0 3892 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_7_0
timestamp 1607101874
transform -1 0 3932 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_7_1
timestamp 1607101874
transform -1 0 3940 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_109
timestamp 1607101874
transform -1 0 3972 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_614
timestamp 1607101874
transform 1 0 3972 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_468
timestamp 1607101874
transform -1 0 4028 0 1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_118
timestamp 1607101874
transform 1 0 4028 0 1 3705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_750
timestamp 1607101874
transform 1 0 4076 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_64
timestamp 1607101874
transform -1 0 4188 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_420
timestamp 1607101874
transform -1 0 4220 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_973
timestamp 1607101874
transform 1 0 4220 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_132
timestamp 1607101874
transform -1 0 4332 0 1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_123
timestamp 1607101874
transform 1 0 4332 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1607101874
transform 1 0 4364 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_8_0
timestamp 1607101874
transform -1 0 4404 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_8_1
timestamp 1607101874
transform -1 0 4412 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_766
timestamp 1607101874
transform -1 0 4508 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_977
timestamp 1607101874
transform -1 0 4604 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_1047
timestamp 1607101874
transform 1 0 4604 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_292
timestamp 1607101874
transform 1 0 4636 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_195
timestamp 1607101874
transform 1 0 4660 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_658
timestamp 1607101874
transform 1 0 4692 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_42
timestamp 1607101874
transform 1 0 4788 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_41
timestamp 1607101874
transform -1 0 4852 0 1 3705
box -2 -3 34 103
use AND2X2  AND2X2_36
timestamp 1607101874
transform 1 0 4852 0 1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_382
timestamp 1607101874
transform -1 0 4916 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_407
timestamp 1607101874
transform 1 0 4916 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_9_0
timestamp 1607101874
transform -1 0 4956 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_9_1
timestamp 1607101874
transform -1 0 4964 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_408
timestamp 1607101874
transform -1 0 4996 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1607101874
transform -1 0 5092 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_415
timestamp 1607101874
transform -1 0 5124 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1607101874
transform 1 0 5124 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_428
timestamp 1607101874
transform -1 0 5188 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1607101874
transform -1 0 5284 0 1 3705
box -2 -3 98 103
use NOR2X1  NOR2X1_290
timestamp 1607101874
transform -1 0 5308 0 1 3705
box -2 -3 26 103
use NOR3X1  NOR3X1_5
timestamp 1607101874
transform -1 0 68 0 -1 3905
box -2 -3 66 103
use OAI21X1  OAI21X1_481
timestamp 1607101874
transform 1 0 68 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_452
timestamp 1607101874
transform -1 0 132 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_459
timestamp 1607101874
transform -1 0 164 0 -1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_210
timestamp 1607101874
transform 1 0 164 0 -1 3905
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1607101874
transform 1 0 196 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_456
timestamp 1607101874
transform 1 0 228 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_108
timestamp 1607101874
transform 1 0 260 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_457
timestamp 1607101874
transform -1 0 316 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_0_0
timestamp 1607101874
transform -1 0 324 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_0_1
timestamp 1607101874
transform -1 0 332 0 -1 3905
box -2 -3 10 103
use MUX2X1  MUX2X1_175
timestamp 1607101874
transform -1 0 380 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_450
timestamp 1607101874
transform 1 0 380 0 -1 3905
box -2 -3 34 103
use AOI22X1  AOI22X1_3
timestamp 1607101874
transform -1 0 452 0 -1 3905
box -2 -3 42 103
use NAND3X1  NAND3X1_15
timestamp 1607101874
transform 1 0 452 0 -1 3905
box -2 -3 34 103
use AND2X2  AND2X2_5
timestamp 1607101874
transform 1 0 484 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_306
timestamp 1607101874
transform 1 0 516 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_117
timestamp 1607101874
transform -1 0 564 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_215
timestamp 1607101874
transform 1 0 564 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1607101874
transform -1 0 692 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_463
timestamp 1607101874
transform 1 0 692 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1607101874
transform 1 0 724 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_1_0
timestamp 1607101874
transform 1 0 820 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_1_1
timestamp 1607101874
transform 1 0 828 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_410
timestamp 1607101874
transform 1 0 836 0 -1 3905
box -2 -3 98 103
use AOI21X1  AOI21X1_578
timestamp 1607101874
transform 1 0 932 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_690
timestamp 1607101874
transform 1 0 964 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_233
timestamp 1607101874
transform -1 0 1012 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_73
timestamp 1607101874
transform -1 0 1044 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_753
timestamp 1607101874
transform -1 0 1076 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_534
timestamp 1607101874
transform 1 0 1076 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_571
timestamp 1607101874
transform 1 0 1100 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_683
timestamp 1607101874
transform -1 0 1156 0 -1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_533
timestamp 1607101874
transform -1 0 1180 0 -1 3905
box -2 -3 26 103
use OAI22X1  OAI22X1_53
timestamp 1607101874
transform 1 0 1180 0 -1 3905
box -2 -3 42 103
use AOI21X1  AOI21X1_334
timestamp 1607101874
transform -1 0 1252 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_888
timestamp 1607101874
transform -1 0 1348 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_2_0
timestamp 1607101874
transform 1 0 1348 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_2_1
timestamp 1607101874
transform 1 0 1356 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_203
timestamp 1607101874
transform 1 0 1364 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_202
timestamp 1607101874
transform -1 0 1428 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_758
timestamp 1607101874
transform -1 0 1460 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_335
timestamp 1607101874
transform 1 0 1460 0 -1 3905
box -2 -3 18 103
use BUFX4  BUFX4_143
timestamp 1607101874
transform -1 0 1508 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_269
timestamp 1607101874
transform 1 0 1508 0 -1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_701
timestamp 1607101874
transform -1 0 1628 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_589
timestamp 1607101874
transform -1 0 1660 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_532
timestamp 1607101874
transform 1 0 1660 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_219
timestamp 1607101874
transform 1 0 1684 0 -1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_230
timestamp 1607101874
transform 1 0 1708 0 -1 3905
box -2 -3 50 103
use NOR2X1  NOR2X1_535
timestamp 1607101874
transform -1 0 1780 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_119
timestamp 1607101874
transform -1 0 1812 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_579
timestamp 1607101874
transform 1 0 1812 0 -1 3905
box -2 -3 34 103
use INVX8  INVX8_4
timestamp 1607101874
transform -1 0 1884 0 -1 3905
box -2 -3 42 103
use FILL  FILL_38_3_0
timestamp 1607101874
transform 1 0 1884 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_3_1
timestamp 1607101874
transform 1 0 1892 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1208
timestamp 1607101874
transform 1 0 1900 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1117
timestamp 1607101874
transform 1 0 1932 0 -1 3905
box -2 -3 34 103
use OAI22X1  OAI22X1_55
timestamp 1607101874
transform 1 0 1964 0 -1 3905
box -2 -3 42 103
use BUFX4  BUFX4_68
timestamp 1607101874
transform 1 0 2004 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1187
timestamp 1607101874
transform 1 0 2036 0 -1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_496
timestamp 1607101874
transform -1 0 2100 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1188
timestamp 1607101874
transform 1 0 2100 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_584
timestamp 1607101874
transform 1 0 2132 0 -1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_729
timestamp 1607101874
transform -1 0 2252 0 -1 3905
box -2 -3 98 103
use AOI21X1  AOI21X1_43
timestamp 1607101874
transform 1 0 2252 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_82
timestamp 1607101874
transform 1 0 2284 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_145
timestamp 1607101874
transform 1 0 2308 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_225
timestamp 1607101874
transform 1 0 2340 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_4_0
timestamp 1607101874
transform 1 0 2372 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_4_1
timestamp 1607101874
transform 1 0 2380 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_915
timestamp 1607101874
transform 1 0 2388 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_232
timestamp 1607101874
transform -1 0 2516 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_917
timestamp 1607101874
transform 1 0 2516 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_228
timestamp 1607101874
transform -1 0 2644 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1607101874
transform -1 0 2676 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1607101874
transform 1 0 2676 0 -1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_329
timestamp 1607101874
transform 1 0 2708 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_372
timestamp 1607101874
transform -1 0 2836 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_363
timestamp 1607101874
transform 1 0 2836 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1322
timestamp 1607101874
transform -1 0 2884 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_5_0
timestamp 1607101874
transform 1 0 2884 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_5_1
timestamp 1607101874
transform 1 0 2892 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_936
timestamp 1607101874
transform 1 0 2900 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1607101874
transform 1 0 2932 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_364
timestamp 1607101874
transform 1 0 3028 0 -1 3905
box -2 -3 18 103
use MUX2X1  MUX2X1_292
timestamp 1607101874
transform -1 0 3092 0 -1 3905
box -2 -3 50 103
use NOR2X1  NOR2X1_90
timestamp 1607101874
transform -1 0 3116 0 -1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_344
timestamp 1607101874
transform 1 0 3116 0 -1 3905
box -2 -3 50 103
use INVX1  INVX1_357
timestamp 1607101874
transform -1 0 3180 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_408
timestamp 1607101874
transform -1 0 3276 0 -1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_67
timestamp 1607101874
transform 1 0 3276 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_55
timestamp 1607101874
transform 1 0 3300 0 -1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_306
timestamp 1607101874
transform 1 0 3332 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_674
timestamp 1607101874
transform -1 0 3396 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_133
timestamp 1607101874
transform -1 0 3412 0 -1 3905
box -2 -3 18 103
use FILL  FILL_38_6_0
timestamp 1607101874
transform -1 0 3420 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_6_1
timestamp 1607101874
transform -1 0 3428 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_979
timestamp 1607101874
transform -1 0 3524 0 -1 3905
box -2 -3 98 103
use MUX2X1  MUX2X1_120
timestamp 1607101874
transform 1 0 3524 0 -1 3905
box -2 -3 50 103
use NAND2X1  NAND2X1_69
timestamp 1607101874
transform 1 0 3572 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_126
timestamp 1607101874
transform 1 0 3596 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_177
timestamp 1607101874
transform -1 0 3660 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_216
timestamp 1607101874
transform 1 0 3660 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_136
timestamp 1607101874
transform -1 0 3716 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_54
timestamp 1607101874
transform 1 0 3716 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1607101874
transform -1 0 3844 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1308
timestamp 1607101874
transform -1 0 3876 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1309
timestamp 1607101874
transform -1 0 3908 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_7_0
timestamp 1607101874
transform 1 0 3908 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_7_1
timestamp 1607101874
transform 1 0 3916 0 -1 3905
box -2 -3 10 103
use BUFX4  BUFX4_25
timestamp 1607101874
transform 1 0 3924 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_224
timestamp 1607101874
transform 1 0 3956 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_131
timestamp 1607101874
transform -1 0 3996 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_971
timestamp 1607101874
transform -1 0 4092 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1331
timestamp 1607101874
transform 1 0 4092 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_355
timestamp 1607101874
transform -1 0 4148 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_415
timestamp 1607101874
transform -1 0 4164 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_341
timestamp 1607101874
transform -1 0 4260 0 -1 3905
box -2 -3 98 103
use MUX2X1  MUX2X1_119
timestamp 1607101874
transform -1 0 4308 0 -1 3905
box -2 -3 50 103
use AOI21X1  AOI21X1_313
timestamp 1607101874
transform 1 0 4308 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1193
timestamp 1607101874
transform 1 0 4340 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_344
timestamp 1607101874
transform -1 0 4396 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_715
timestamp 1607101874
transform -1 0 4428 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_8_0
timestamp 1607101874
transform 1 0 4428 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_8_1
timestamp 1607101874
transform 1 0 4436 0 -1 3905
box -2 -3 10 103
use NOR2X1  NOR2X1_95
timestamp 1607101874
transform 1 0 4444 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_51
timestamp 1607101874
transform -1 0 4500 0 -1 3905
box -2 -3 34 103
use OAI22X1  OAI22X1_70
timestamp 1607101874
transform 1 0 4500 0 -1 3905
box -2 -3 42 103
use MUX2X1  MUX2X1_168
timestamp 1607101874
transform 1 0 4540 0 -1 3905
box -2 -3 50 103
use INVX1  INVX1_182
timestamp 1607101874
transform -1 0 4604 0 -1 3905
box -2 -3 18 103
use NOR2X1  NOR2X1_439
timestamp 1607101874
transform 1 0 4604 0 -1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1607101874
transform -1 0 4724 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_412
timestamp 1607101874
transform 1 0 4724 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1607101874
transform 1 0 4756 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_411
timestamp 1607101874
transform 1 0 4852 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_608
timestamp 1607101874
transform 1 0 4884 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_481
timestamp 1607101874
transform 1 0 4908 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_9_0
timestamp 1607101874
transform 1 0 4940 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_9_1
timestamp 1607101874
transform 1 0 4948 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1150
timestamp 1607101874
transform 1 0 4956 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1239
timestamp 1607101874
transform 1 0 4988 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_338
timestamp 1607101874
transform 1 0 5020 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1607101874
transform -1 0 5148 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_416
timestamp 1607101874
transform -1 0 5180 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_107
timestamp 1607101874
transform -1 0 5204 0 -1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_799
timestamp 1607101874
transform -1 0 5300 0 -1 3905
box -2 -3 98 103
use FILL  FILL_39_1
timestamp 1607101874
transform -1 0 5308 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_476
timestamp 1607101874
transform -1 0 36 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_308
timestamp 1607101874
transform -1 0 60 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_223
timestamp 1607101874
transform -1 0 92 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_339
timestamp 1607101874
transform -1 0 116 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_472
timestamp 1607101874
transform 1 0 116 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_473
timestamp 1607101874
transform -1 0 180 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_194
timestamp 1607101874
transform 1 0 180 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_195
timestamp 1607101874
transform 1 0 196 0 1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_32
timestamp 1607101874
transform -1 0 244 0 1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_36
timestamp 1607101874
transform 1 0 244 0 1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1607101874
transform -1 0 308 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1607101874
transform -1 0 332 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_0_0
timestamp 1607101874
transform -1 0 340 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_0_1
timestamp 1607101874
transform -1 0 348 0 1 3905
box -2 -3 10 103
use NAND3X1  NAND3X1_20
timestamp 1607101874
transform -1 0 380 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_458
timestamp 1607101874
transform 1 0 380 0 1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1607101874
transform -1 0 444 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1607101874
transform 1 0 444 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_464
timestamp 1607101874
transform 1 0 476 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_310
timestamp 1607101874
transform -1 0 532 0 1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_305
timestamp 1607101874
transform -1 0 556 0 1 3905
box -2 -3 26 103
use NAND3X1  NAND3X1_25
timestamp 1607101874
transform -1 0 588 0 1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1607101874
transform -1 0 620 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_465
timestamp 1607101874
transform -1 0 652 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_454
timestamp 1607101874
transform 1 0 652 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_193
timestamp 1607101874
transform 1 0 684 0 1 3905
box -2 -3 18 103
use AOI21X1  AOI21X1_214
timestamp 1607101874
transform 1 0 700 0 1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_576
timestamp 1607101874
transform 1 0 732 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_688
timestamp 1607101874
transform 1 0 764 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_575
timestamp 1607101874
transform 1 0 788 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_687
timestamp 1607101874
transform 1 0 820 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_1_0
timestamp 1607101874
transform 1 0 844 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_1_1
timestamp 1607101874
transform 1 0 852 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1607101874
transform 1 0 860 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1405
timestamp 1607101874
transform 1 0 956 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1404
timestamp 1607101874
transform -1 0 1020 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1401
timestamp 1607101874
transform 1 0 1020 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1400
timestamp 1607101874
transform 1 0 1052 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1607101874
transform 1 0 1084 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1607101874
transform 1 0 1180 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1407
timestamp 1607101874
transform 1 0 1276 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1406
timestamp 1607101874
transform -1 0 1340 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_403
timestamp 1607101874
transform -1 0 1372 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_2_0
timestamp 1607101874
transform 1 0 1372 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_2_1
timestamp 1607101874
transform 1 0 1380 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_757
timestamp 1607101874
transform 1 0 1388 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_234
timestamp 1607101874
transform -1 0 1444 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_387
timestamp 1607101874
transform -1 0 1476 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_407
timestamp 1607101874
transform -1 0 1508 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1398
timestamp 1607101874
transform 1 0 1508 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_421
timestamp 1607101874
transform 1 0 1540 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1607101874
transform 1 0 1564 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1395
timestamp 1607101874
transform 1 0 1660 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1394
timestamp 1607101874
transform -1 0 1724 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_406
timestamp 1607101874
transform -1 0 1756 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1419
timestamp 1607101874
transform 1 0 1756 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1418
timestamp 1607101874
transform -1 0 1820 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_416
timestamp 1607101874
transform -1 0 1916 0 1 3905
box -2 -3 98 103
use FILL  FILL_39_3_0
timestamp 1607101874
transform 1 0 1916 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_3_1
timestamp 1607101874
transform 1 0 1924 0 1 3905
box -2 -3 10 103
use NOR2X1  NOR2X1_158
timestamp 1607101874
transform 1 0 1932 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_474
timestamp 1607101874
transform 1 0 1956 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1110
timestamp 1607101874
transform -1 0 2020 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1112
timestamp 1607101874
transform -1 0 2052 0 1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_475
timestamp 1607101874
transform 1 0 2052 0 1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_356
timestamp 1607101874
transform 1 0 2084 0 1 3905
box -2 -3 50 103
use BUFX4  BUFX4_216
timestamp 1607101874
transform 1 0 2132 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1111
timestamp 1607101874
transform -1 0 2196 0 1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_265
timestamp 1607101874
transform 1 0 2196 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_265
timestamp 1607101874
transform -1 0 2324 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1437
timestamp 1607101874
transform 1 0 2324 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1436
timestamp 1607101874
transform -1 0 2388 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_4_0
timestamp 1607101874
transform -1 0 2396 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_4_1
timestamp 1607101874
transform -1 0 2404 0 1 3905
box -2 -3 10 103
use AOI21X1  AOI21X1_266
timestamp 1607101874
transform -1 0 2436 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_931
timestamp 1607101874
transform -1 0 2532 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_233
timestamp 1607101874
transform -1 0 2564 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_173
timestamp 1607101874
transform -1 0 2588 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1607101874
transform 1 0 2588 0 1 3905
box -2 -3 98 103
use INVX1  INVX1_305
timestamp 1607101874
transform 1 0 2684 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1607101874
transform -1 0 2796 0 1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_697
timestamp 1607101874
transform 1 0 2796 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_585
timestamp 1607101874
transform -1 0 2852 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_354
timestamp 1607101874
transform -1 0 2876 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_383
timestamp 1607101874
transform 1 0 2876 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_5_0
timestamp 1607101874
transform 1 0 2908 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_5_1
timestamp 1607101874
transform 1 0 2916 0 1 3905
box -2 -3 10 103
use BUFX4  BUFX4_384
timestamp 1607101874
transform 1 0 2924 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_445
timestamp 1607101874
transform 1 0 2956 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_359
timestamp 1607101874
transform 1 0 3052 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1455
timestamp 1607101874
transform -1 0 3108 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_380
timestamp 1607101874
transform 1 0 3108 0 1 3905
box -2 -3 18 103
use AOI21X1  AOI21X1_407
timestamp 1607101874
transform -1 0 3156 0 1 3905
box -2 -3 34 103
use OAI22X1  OAI22X1_39
timestamp 1607101874
transform 1 0 3156 0 1 3905
box -2 -3 42 103
use NOR2X1  NOR2X1_91
timestamp 1607101874
transform -1 0 3220 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1607101874
transform -1 0 3316 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1311
timestamp 1607101874
transform 1 0 3316 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1310
timestamp 1607101874
transform -1 0 3380 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1320
timestamp 1607101874
transform 1 0 3380 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_6_0
timestamp 1607101874
transform -1 0 3420 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_6_1
timestamp 1607101874
transform -1 0 3428 0 1 3905
box -2 -3 10 103
use NOR2X1  NOR2X1_210
timestamp 1607101874
transform -1 0 3452 0 1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_213
timestamp 1607101874
transform 1 0 3452 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_417
timestamp 1607101874
transform 1 0 3476 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_958
timestamp 1607101874
transform -1 0 3540 0 1 3905
box -2 -3 34 103
use INVX8  INVX8_23
timestamp 1607101874
transform 1 0 3540 0 1 3905
box -2 -3 42 103
use AOI21X1  AOI21X1_420
timestamp 1607101874
transform -1 0 3612 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_959
timestamp 1607101874
transform 1 0 3612 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_186
timestamp 1607101874
transform -1 0 3668 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1457
timestamp 1607101874
transform 1 0 3668 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1458
timestamp 1607101874
transform -1 0 3732 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_455
timestamp 1607101874
transform -1 0 3828 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_444
timestamp 1607101874
transform 1 0 3828 0 1 3905
box -2 -3 98 103
use FILL  FILL_39_7_0
timestamp 1607101874
transform 1 0 3924 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_7_1
timestamp 1607101874
transform 1 0 3932 0 1 3905
box -2 -3 10 103
use AOI21X1  AOI21X1_590
timestamp 1607101874
transform 1 0 3940 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_702
timestamp 1607101874
transform -1 0 3996 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_240
timestamp 1607101874
transform 1 0 3996 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_70
timestamp 1607101874
transform 1 0 4020 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_530
timestamp 1607101874
transform -1 0 4076 0 1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_51
timestamp 1607101874
transform 1 0 4076 0 1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_747
timestamp 1607101874
transform 1 0 4124 0 1 3905
box -2 -3 98 103
use INVX1  INVX1_61
timestamp 1607101874
transform 1 0 4220 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_710
timestamp 1607101874
transform 1 0 4236 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_471
timestamp 1607101874
transform -1 0 4300 0 1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_206
timestamp 1607101874
transform 1 0 4300 0 1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_117
timestamp 1607101874
transform 1 0 4348 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_762
timestamp 1607101874
transform -1 0 4476 0 1 3905
box -2 -3 98 103
use FILL  FILL_39_8_0
timestamp 1607101874
transform -1 0 4484 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_8_1
timestamp 1607101874
transform -1 0 4492 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1195
timestamp 1607101874
transform -1 0 4524 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1607101874
transform 1 0 4524 0 1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_39
timestamp 1607101874
transform -1 0 4644 0 1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_58
timestamp 1607101874
transform 1 0 4644 0 1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_656
timestamp 1607101874
transform 1 0 4692 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_38
timestamp 1607101874
transform 1 0 4788 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_37
timestamp 1607101874
transform -1 0 4852 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_438
timestamp 1607101874
transform 1 0 4852 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_808
timestamp 1607101874
transform 1 0 4876 0 1 3905
box -2 -3 34 103
use AND2X2  AND2X2_51
timestamp 1607101874
transform 1 0 4908 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_9_0
timestamp 1607101874
transform 1 0 4940 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_9_1
timestamp 1607101874
transform 1 0 4948 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_40
timestamp 1607101874
transform 1 0 4956 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_39
timestamp 1607101874
transform 1 0 4988 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_657
timestamp 1607101874
transform 1 0 5020 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1237
timestamp 1607101874
transform -1 0 5148 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_806
timestamp 1607101874
transform -1 0 5180 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1607101874
transform 1 0 5180 0 1 3905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_100
timestamp 1607101874
transform -1 0 5284 0 1 3905
box -2 -3 74 103
use FILL  FILL_40_1
timestamp 1607101874
transform 1 0 5284 0 1 3905
box -2 -3 10 103
use FILL  FILL_40_2
timestamp 1607101874
transform 1 0 5292 0 1 3905
box -2 -3 10 103
use FILL  FILL_40_3
timestamp 1607101874
transform 1 0 5300 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_424
timestamp 1607101874
transform -1 0 100 0 -1 4105
box -2 -3 98 103
use XOR2X1  XOR2X1_1
timestamp 1607101874
transform -1 0 156 0 -1 4105
box -2 -3 58 103
use NAND2X1  NAND2X1_132
timestamp 1607101874
transform -1 0 180 0 -1 4105
box -2 -3 26 103
use NOR3X1  NOR3X1_4
timestamp 1607101874
transform 1 0 180 0 -1 4105
box -2 -3 66 103
use INVX4  INVX4_8
timestamp 1607101874
transform 1 0 244 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_130
timestamp 1607101874
transform -1 0 292 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_19
timestamp 1607101874
transform -1 0 324 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_0_0
timestamp 1607101874
transform -1 0 332 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_0_1
timestamp 1607101874
transform -1 0 340 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_487
timestamp 1607101874
transform -1 0 372 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_318
timestamp 1607101874
transform -1 0 396 0 -1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_311
timestamp 1607101874
transform 1 0 396 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_124
timestamp 1607101874
transform -1 0 444 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_24
timestamp 1607101874
transform -1 0 476 0 -1 4105
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1607101874
transform 1 0 476 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_214
timestamp 1607101874
transform 1 0 508 0 -1 4105
box -2 -3 18 103
use AOI21X1  AOI21X1_221
timestamp 1607101874
transform 1 0 524 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_220
timestamp 1607101874
transform -1 0 588 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_126
timestamp 1607101874
transform -1 0 612 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_119
timestamp 1607101874
transform 1 0 612 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_31
timestamp 1607101874
transform 1 0 636 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_113
timestamp 1607101874
transform 1 0 668 0 -1 4105
box -2 -3 26 103
use INVX4  INVX4_7
timestamp 1607101874
transform -1 0 716 0 -1 4105
box -2 -3 26 103
use INVX2  INVX2_14
timestamp 1607101874
transform -1 0 732 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_419
timestamp 1607101874
transform -1 0 828 0 -1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_356
timestamp 1607101874
transform -1 0 852 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_1_0
timestamp 1607101874
transform -1 0 860 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_1_1
timestamp 1607101874
transform -1 0 868 0 -1 4105
box -2 -3 10 103
use INVX1  INVX1_192
timestamp 1607101874
transform -1 0 884 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_545
timestamp 1607101874
transform -1 0 916 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_546
timestamp 1607101874
transform 1 0 916 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_420
timestamp 1607101874
transform -1 0 1044 0 -1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1607101874
transform -1 0 1140 0 -1 4105
box -2 -3 98 103
use AOI21X1  AOI21X1_572
timestamp 1607101874
transform 1 0 1140 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_684
timestamp 1607101874
transform -1 0 1196 0 -1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1607101874
transform 1 0 1196 0 -1 4105
box -2 -3 98 103
use AOI21X1  AOI21X1_95
timestamp 1607101874
transform 1 0 1292 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_159
timestamp 1607101874
transform -1 0 1348 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_2_0
timestamp 1607101874
transform 1 0 1348 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_2_1
timestamp 1607101874
transform 1 0 1356 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_755
timestamp 1607101874
transform 1 0 1364 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_756
timestamp 1607101874
transform 1 0 1396 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_216
timestamp 1607101874
transform 1 0 1428 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1392
timestamp 1607101874
transform 1 0 1452 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1393
timestamp 1607101874
transform -1 0 1516 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_570
timestamp 1607101874
transform 1 0 1516 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_682
timestamp 1607101874
transform -1 0 1572 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1399
timestamp 1607101874
transform -1 0 1604 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1607101874
transform -1 0 1700 0 -1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_370
timestamp 1607101874
transform -1 0 1724 0 -1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_247
timestamp 1607101874
transform 1 0 1724 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_371
timestamp 1607101874
transform 1 0 1756 0 -1 4105
box -2 -3 26 103
use OAI22X1  OAI22X1_74
timestamp 1607101874
transform 1 0 1780 0 -1 4105
box -2 -3 42 103
use OAI21X1  OAI21X1_1207
timestamp 1607101874
transform -1 0 1852 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_588
timestamp 1607101874
transform -1 0 1876 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_3_0
timestamp 1607101874
transform -1 0 1884 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_3_1
timestamp 1607101874
transform -1 0 1892 0 -1 4105
box -2 -3 10 103
use BUFX4  BUFX4_148
timestamp 1607101874
transform -1 0 1924 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_692
timestamp 1607101874
transform -1 0 1956 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_202
timestamp 1607101874
transform -1 0 2004 0 -1 4105
box -2 -3 50 103
use INVX1  INVX1_421
timestamp 1607101874
transform -1 0 2020 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1607101874
transform -1 0 2116 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_580
timestamp 1607101874
transform 1 0 2116 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_203
timestamp 1607101874
transform -1 0 2196 0 -1 4105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_726
timestamp 1607101874
transform 1 0 2196 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_55
timestamp 1607101874
transform 1 0 2292 0 -1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_45
timestamp 1607101874
transform 1 0 2308 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_995
timestamp 1607101874
transform 1 0 2356 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_4_0
timestamp 1607101874
transform 1 0 2388 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_4_1
timestamp 1607101874
transform 1 0 2396 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1203
timestamp 1607101874
transform 1 0 2404 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1202
timestamp 1607101874
transform -1 0 2468 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_934
timestamp 1607101874
transform 1 0 2468 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_239
timestamp 1607101874
transform 1 0 2564 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_238
timestamp 1607101874
transform -1 0 2628 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_138
timestamp 1607101874
transform -1 0 2660 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_141
timestamp 1607101874
transform 1 0 2660 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_351
timestamp 1607101874
transform -1 0 2740 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_748
timestamp 1607101874
transform -1 0 2772 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1432
timestamp 1607101874
transform 1 0 2772 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1433
timestamp 1607101874
transform -1 0 2836 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1607101874
transform 1 0 2836 0 -1 4105
box -2 -3 98 103
use FILL  FILL_40_5_0
timestamp 1607101874
transform -1 0 2940 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_5_1
timestamp 1607101874
transform -1 0 2948 0 -1 4105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_39
timestamp 1607101874
transform -1 0 3020 0 -1 4105
box -2 -3 74 103
use BUFX4  BUFX4_317
timestamp 1607101874
transform 1 0 3020 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_358
timestamp 1607101874
transform 1 0 3052 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1454
timestamp 1607101874
transform -1 0 3108 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_443
timestamp 1607101874
transform 1 0 3108 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_258
timestamp 1607101874
transform 1 0 3204 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_601
timestamp 1607101874
transform 1 0 3220 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_276
timestamp 1607101874
transform 1 0 3252 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_600
timestamp 1607101874
transform 1 0 3284 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_172
timestamp 1607101874
transform -1 0 3348 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1321
timestamp 1607101874
transform 1 0 3348 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_6_0
timestamp 1607101874
transform 1 0 3380 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_6_1
timestamp 1607101874
transform 1 0 3388 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_377
timestamp 1607101874
transform 1 0 3396 0 -1 4105
box -2 -3 98 103
use AOI21X1  AOI21X1_134
timestamp 1607101874
transform 1 0 3492 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_292
timestamp 1607101874
transform -1 0 3620 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1451
timestamp 1607101874
transform 1 0 3620 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1450
timestamp 1607101874
transform -1 0 3684 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_962
timestamp 1607101874
transform -1 0 3716 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_419
timestamp 1607101874
transform 1 0 3716 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_961
timestamp 1607101874
transform -1 0 3780 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_471
timestamp 1607101874
transform 1 0 3780 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_256
timestamp 1607101874
transform 1 0 3876 0 -1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_360
timestamp 1607101874
transform 1 0 3892 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_7_0
timestamp 1607101874
transform -1 0 3924 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_7_1
timestamp 1607101874
transform -1 0 3932 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1456
timestamp 1607101874
transform -1 0 3964 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_315
timestamp 1607101874
transform 1 0 3964 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_372
timestamp 1607101874
transform -1 0 4044 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_597
timestamp 1607101874
transform 1 0 4044 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_213
timestamp 1607101874
transform -1 0 4124 0 -1 4105
box -2 -3 50 103
use NAND2X1  NAND2X1_337
timestamp 1607101874
transform 1 0 4124 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_775
timestamp 1607101874
transform 1 0 4148 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_212
timestamp 1607101874
transform 1 0 4180 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_598
timestamp 1607101874
transform 1 0 4228 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1158
timestamp 1607101874
transform -1 0 4292 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_147
timestamp 1607101874
transform 1 0 4292 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_203
timestamp 1607101874
transform -1 0 4348 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_118
timestamp 1607101874
transform 1 0 4348 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_126
timestamp 1607101874
transform -1 0 4412 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_8_0
timestamp 1607101874
transform 1 0 4412 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_8_1
timestamp 1607101874
transform 1 0 4420 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_763
timestamp 1607101874
transform 1 0 4428 0 -1 4105
box -2 -3 98 103
use BUFX4  BUFX4_444
timestamp 1607101874
transform -1 0 4556 0 -1 4105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_46
timestamp 1607101874
transform -1 0 4628 0 -1 4105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_452
timestamp 1607101874
transform -1 0 4724 0 -1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_774
timestamp 1607101874
transform -1 0 4820 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_68
timestamp 1607101874
transform -1 0 4836 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_758
timestamp 1607101874
transform -1 0 4932 0 -1 4105
box -2 -3 98 103
use FILL  FILL_40_9_0
timestamp 1607101874
transform -1 0 4940 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_9_1
timestamp 1607101874
transform -1 0 4948 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_662
timestamp 1607101874
transform -1 0 5044 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_50
timestamp 1607101874
transform 1 0 5044 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1607101874
transform -1 0 5108 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_419
timestamp 1607101874
transform 1 0 5108 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_420
timestamp 1607101874
transform -1 0 5172 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_162
timestamp 1607101874
transform -1 0 5188 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1607101874
transform -1 0 5284 0 -1 4105
box -2 -3 98 103
use FILL  FILL_41_1
timestamp 1607101874
transform -1 0 5292 0 -1 4105
box -2 -3 10 103
use FILL  FILL_41_2
timestamp 1607101874
transform -1 0 5300 0 -1 4105
box -2 -3 10 103
use FILL  FILL_41_3
timestamp 1607101874
transform -1 0 5308 0 -1 4105
box -2 -3 10 103
use NAND2X1  NAND2X1_160
timestamp 1607101874
transform 1 0 4 0 1 4105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_5
timestamp 1607101874
transform -1 0 84 0 1 4105
box -2 -3 58 103
use OAI21X1  OAI21X1_485
timestamp 1607101874
transform -1 0 116 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1607101874
transform 1 0 116 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_315
timestamp 1607101874
transform 1 0 140 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_479
timestamp 1607101874
transform 1 0 164 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_196
timestamp 1607101874
transform 1 0 196 0 1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_57
timestamp 1607101874
transform 1 0 212 0 1 4105
box -2 -3 34 103
use INVX2  INVX2_18
timestamp 1607101874
transform -1 0 260 0 1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_326
timestamp 1607101874
transform 1 0 260 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_488
timestamp 1607101874
transform 1 0 284 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_201
timestamp 1607101874
transform -1 0 332 0 1 4105
box -2 -3 18 103
use FILL  FILL_41_0_0
timestamp 1607101874
transform 1 0 332 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_0_1
timestamp 1607101874
transform 1 0 340 0 1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_489
timestamp 1607101874
transform 1 0 348 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_402
timestamp 1607101874
transform 1 0 380 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_474
timestamp 1607101874
transform -1 0 508 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1607101874
transform 1 0 508 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_351
timestamp 1607101874
transform -1 0 564 0 1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_37
timestamp 1607101874
transform -1 0 596 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1607101874
transform -1 0 628 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_190
timestamp 1607101874
transform -1 0 644 0 1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_16
timestamp 1607101874
transform -1 0 676 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_471
timestamp 1607101874
transform -1 0 708 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_451
timestamp 1607101874
transform 1 0 708 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1607101874
transform 1 0 740 0 1 4105
box -2 -3 26 103
use NOR3X1  NOR3X1_6
timestamp 1607101874
transform 1 0 764 0 1 4105
box -2 -3 66 103
use NOR2X1  NOR2X1_350
timestamp 1607101874
transform 1 0 828 0 1 4105
box -2 -3 26 103
use FILL  FILL_41_1_0
timestamp 1607101874
transform 1 0 852 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_1_1
timestamp 1607101874
transform 1 0 860 0 1 4105
box -2 -3 10 103
use NAND2X1  NAND2X1_168
timestamp 1607101874
transform 1 0 868 0 1 4105
box -2 -3 26 103
use OR2X2  OR2X2_7
timestamp 1607101874
transform 1 0 892 0 1 4105
box -2 -3 34 103
use XOR2X1  XOR2X1_4
timestamp 1607101874
transform -1 0 980 0 1 4105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_418
timestamp 1607101874
transform -1 0 1076 0 1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_891
timestamp 1607101874
transform 1 0 1076 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_209
timestamp 1607101874
transform 1 0 1172 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_208
timestamp 1607101874
transform -1 0 1236 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1413
timestamp 1607101874
transform 1 0 1236 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1412
timestamp 1607101874
transform -1 0 1300 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_895
timestamp 1607101874
transform 1 0 1300 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_2_0
timestamp 1607101874
transform 1 0 1396 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_2_1
timestamp 1607101874
transform 1 0 1404 0 1 4105
box -2 -3 10 103
use INVX1  INVX1_285
timestamp 1607101874
transform 1 0 1412 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_689
timestamp 1607101874
transform 1 0 1428 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1390
timestamp 1607101874
transform 1 0 1460 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1391
timestamp 1607101874
transform -1 0 1524 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_335
timestamp 1607101874
transform -1 0 1556 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_311
timestamp 1607101874
transform -1 0 1572 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1607101874
transform -1 0 1668 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_582
timestamp 1607101874
transform -1 0 1700 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1607101874
transform -1 0 1796 0 1 4105
box -2 -3 98 103
use BUFX4  BUFX4_408
timestamp 1607101874
transform 1 0 1796 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_843
timestamp 1607101874
transform -1 0 1860 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_3_0
timestamp 1607101874
transform 1 0 1860 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_3_1
timestamp 1607101874
transform 1 0 1868 0 1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_214
timestamp 1607101874
transform 1 0 1876 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_215
timestamp 1607101874
transform 1 0 1908 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_894
timestamp 1607101874
transform 1 0 1940 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_287
timestamp 1607101874
transform -1 0 2052 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_192
timestamp 1607101874
transform 1 0 2052 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_193
timestamp 1607101874
transform 1 0 2084 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_262
timestamp 1607101874
transform -1 0 2148 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_201
timestamp 1607101874
transform -1 0 2196 0 1 4105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_883
timestamp 1607101874
transform -1 0 2292 0 1 4105
box -2 -3 98 103
use BUFX4  BUFX4_367
timestamp 1607101874
transform -1 0 2324 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_106
timestamp 1607101874
transform 1 0 2324 0 1 4105
box -2 -3 50 103
use INVX1  INVX1_119
timestamp 1607101874
transform -1 0 2388 0 1 4105
box -2 -3 18 103
use FILL  FILL_41_4_0
timestamp 1607101874
transform 1 0 2388 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_4_1
timestamp 1607101874
transform 1 0 2396 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_926
timestamp 1607101874
transform 1 0 2404 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1201
timestamp 1607101874
transform 1 0 2500 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_498
timestamp 1607101874
transform -1 0 2564 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_465
timestamp 1607101874
transform -1 0 2596 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_850
timestamp 1607101874
transform -1 0 2628 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_235
timestamp 1607101874
transform 1 0 2628 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_234
timestamp 1607101874
transform -1 0 2692 0 1 4105
box -2 -3 34 103
use AND2X2  AND2X2_32
timestamp 1607101874
transform -1 0 2724 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_226
timestamp 1607101874
transform 1 0 2724 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_750
timestamp 1607101874
transform -1 0 2788 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1607101874
transform -1 0 2820 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_916
timestamp 1607101874
transform -1 0 2916 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_5_0
timestamp 1607101874
transform 1 0 2916 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_5_1
timestamp 1607101874
transform 1 0 2924 0 1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1431
timestamp 1607101874
transform 1 0 2932 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1430
timestamp 1607101874
transform -1 0 2996 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_306
timestamp 1607101874
transform 1 0 2996 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_749
timestamp 1607101874
transform 1 0 3012 0 1 4105
box -2 -3 34 103
use INVX8  INVX8_32
timestamp 1607101874
transform -1 0 3084 0 1 4105
box -2 -3 42 103
use OAI21X1  OAI21X1_848
timestamp 1607101874
transform -1 0 3116 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_98
timestamp 1607101874
transform 1 0 3116 0 1 4105
box -2 -3 50 103
use INVX1  INVX1_111
timestamp 1607101874
transform -1 0 3180 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_908
timestamp 1607101874
transform -1 0 3276 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_939
timestamp 1607101874
transform 1 0 3276 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_408
timestamp 1607101874
transform -1 0 3340 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1607101874
transform -1 0 3436 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_6_0
timestamp 1607101874
transform 1 0 3436 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_6_1
timestamp 1607101874
transform 1 0 3444 0 1 4105
box -2 -3 10 103
use NOR2X1  NOR2X1_648
timestamp 1607101874
transform 1 0 3452 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_536
timestamp 1607101874
transform -1 0 3508 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_214
timestamp 1607101874
transform -1 0 3532 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_983
timestamp 1607101874
transform 1 0 3532 0 1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_461
timestamp 1607101874
transform 1 0 3628 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_382
timestamp 1607101874
transform 1 0 3724 0 1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_367
timestamp 1607101874
transform -1 0 3788 0 1 4105
box -2 -3 50 103
use NOR2X1  NOR2X1_196
timestamp 1607101874
transform -1 0 3812 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_457
timestamp 1607101874
transform -1 0 3908 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_7_0
timestamp 1607101874
transform 1 0 3908 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_7_1
timestamp 1607101874
transform 1 0 3916 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_446
timestamp 1607101874
transform 1 0 3924 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_428
timestamp 1607101874
transform 1 0 4020 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1154
timestamp 1607101874
transform 1 0 4036 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_484
timestamp 1607101874
transform -1 0 4100 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1155
timestamp 1607101874
transform 1 0 4100 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_318
timestamp 1607101874
transform 1 0 4132 0 1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_368
timestamp 1607101874
transform 1 0 4148 0 1 4105
box -2 -3 50 103
use AOI21X1  AOI21X1_486
timestamp 1607101874
transform -1 0 4228 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_430
timestamp 1607101874
transform -1 0 4244 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_462
timestamp 1607101874
transform -1 0 4340 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_777
timestamp 1607101874
transform -1 0 4372 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_972
timestamp 1607101874
transform -1 0 4468 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_8_0
timestamp 1607101874
transform 1 0 4468 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_8_1
timestamp 1607101874
transform 1 0 4476 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_472
timestamp 1607101874
transform 1 0 4484 0 1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_712
timestamp 1607101874
transform 1 0 4580 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_600
timestamp 1607101874
transform -1 0 4636 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_237
timestamp 1607101874
transform 1 0 4636 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_704
timestamp 1607101874
transform 1 0 4660 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_592
timestamp 1607101874
transform -1 0 4716 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1245
timestamp 1607101874
transform -1 0 4748 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_72
timestamp 1607101874
transform 1 0 4748 0 1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_62
timestamp 1607101874
transform 1 0 4764 0 1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_711
timestamp 1607101874
transform 1 0 4812 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1607101874
transform 1 0 4844 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_92
timestamp 1607101874
transform -1 0 4900 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_225
timestamp 1607101874
transform -1 0 4924 0 1 4105
box -2 -3 26 103
use FILL  FILL_41_9_0
timestamp 1607101874
transform -1 0 4932 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_9_1
timestamp 1607101874
transform -1 0 4940 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_759
timestamp 1607101874
transform -1 0 5036 0 1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_982
timestamp 1607101874
transform 1 0 5036 0 1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_212
timestamp 1607101874
transform 1 0 5132 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_133
timestamp 1607101874
transform -1 0 5188 0 1 4105
box -2 -3 34 103
use OAI22X1  OAI22X1_41
timestamp 1607101874
transform 1 0 5188 0 1 4105
box -2 -3 42 103
use BUFX4  BUFX4_62
timestamp 1607101874
transform 1 0 5228 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_48
timestamp 1607101874
transform 1 0 5260 0 1 4105
box -2 -3 34 103
use FILL  FILL_42_1
timestamp 1607101874
transform 1 0 5292 0 1 4105
box -2 -3 10 103
use FILL  FILL_42_2
timestamp 1607101874
transform 1 0 5300 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_425
timestamp 1607101874
transform -1 0 100 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_531
timestamp 1607101874
transform -1 0 132 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1607101874
transform -1 0 148 0 -1 4305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_3
timestamp 1607101874
transform -1 0 204 0 -1 4305
box -2 -3 58 103
use NOR2X1  NOR2X1_303
timestamp 1607101874
transform 1 0 204 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_107
timestamp 1607101874
transform 1 0 228 0 -1 4305
box -2 -3 26 103
use XOR2X1  XOR2X1_2
timestamp 1607101874
transform 1 0 252 0 -1 4305
box -2 -3 58 103
use AND2X2  AND2X2_13
timestamp 1607101874
transform 1 0 308 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_0_0
timestamp 1607101874
transform 1 0 340 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_0_1
timestamp 1607101874
transform 1 0 348 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_519
timestamp 1607101874
transform 1 0 356 0 -1 4305
box -2 -3 34 103
use INVX2  INVX2_19
timestamp 1607101874
transform 1 0 388 0 -1 4305
box -2 -3 18 103
use NOR2X1  NOR2X1_316
timestamp 1607101874
transform -1 0 428 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_317
timestamp 1607101874
transform 1 0 428 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_477
timestamp 1607101874
transform 1 0 452 0 -1 4305
box -2 -3 34 103
use AND2X2  AND2X2_8
timestamp 1607101874
transform 1 0 484 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_224
timestamp 1607101874
transform -1 0 548 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_127
timestamp 1607101874
transform -1 0 572 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_189
timestamp 1607101874
transform 1 0 572 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_213
timestamp 1607101874
transform 1 0 588 0 -1 4305
box -2 -3 18 103
use OAI22X1  OAI22X1_3
timestamp 1607101874
transform 1 0 604 0 -1 4305
box -2 -3 42 103
use AOI21X1  AOI21X1_246
timestamp 1607101874
transform -1 0 676 0 -1 4305
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1607101874
transform 1 0 676 0 -1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_540
timestamp 1607101874
transform -1 0 748 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_466
timestamp 1607101874
transform 1 0 748 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1607101874
transform -1 0 804 0 -1 4305
box -2 -3 26 103
use MUX2X1  MUX2X1_174
timestamp 1607101874
transform 1 0 804 0 -1 4305
box -2 -3 50 103
use FILL  FILL_42_1_0
timestamp 1607101874
transform 1 0 852 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_1_1
timestamp 1607101874
transform 1 0 860 0 -1 4305
box -2 -3 10 103
use NAND3X1  NAND3X1_38
timestamp 1607101874
transform 1 0 868 0 -1 4305
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1607101874
transform -1 0 932 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_309
timestamp 1607101874
transform 1 0 932 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_469
timestamp 1607101874
transform -1 0 988 0 -1 4305
box -2 -3 34 103
use NOR3X1  NOR3X1_2
timestamp 1607101874
transform -1 0 1052 0 -1 4305
box -2 -3 66 103
use INVX1  INVX1_215
timestamp 1607101874
transform 1 0 1052 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_70
timestamp 1607101874
transform 1 0 1068 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_355
timestamp 1607101874
transform 1 0 1100 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_166
timestamp 1607101874
transform -1 0 1148 0 -1 4305
box -2 -3 26 103
use AND2X2  AND2X2_16
timestamp 1607101874
transform 1 0 1148 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_218
timestamp 1607101874
transform 1 0 1180 0 -1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1607101874
transform 1 0 1196 0 -1 4305
box -2 -3 98 103
use AOI21X1  AOI21X1_580
timestamp 1607101874
transform 1 0 1292 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_692
timestamp 1607101874
transform -1 0 1348 0 -1 4305
box -2 -3 26 103
use FILL  FILL_42_2_0
timestamp 1607101874
transform 1 0 1348 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_2_1
timestamp 1607101874
transform 1 0 1356 0 -1 4305
box -2 -3 10 103
use BUFX4  BUFX4_436
timestamp 1607101874
transform 1 0 1364 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_537
timestamp 1607101874
transform 1 0 1396 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_536
timestamp 1607101874
transform -1 0 1444 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1115
timestamp 1607101874
transform 1 0 1444 0 -1 4305
box -2 -3 34 103
use OAI22X1  OAI22X1_54
timestamp 1607101874
transform -1 0 1516 0 -1 4305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1607101874
transform 1 0 1516 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_583
timestamp 1607101874
transform 1 0 1612 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_264
timestamp 1607101874
transform 1 0 1644 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1116
timestamp 1607101874
transform -1 0 1708 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_589
timestamp 1607101874
transform 1 0 1708 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1415
timestamp 1607101874
transform 1 0 1732 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1414
timestamp 1607101874
transform 1 0 1764 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_578
timestamp 1607101874
transform -1 0 1828 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_222
timestamp 1607101874
transform 1 0 1828 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_3_0
timestamp 1607101874
transform 1 0 1860 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_3_1
timestamp 1607101874
transform 1 0 1868 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_386
timestamp 1607101874
transform 1 0 1876 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_552
timestamp 1607101874
transform -1 0 2004 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_279
timestamp 1607101874
transform -1 0 2052 0 -1 4305
box -2 -3 50 103
use INVX1  INVX1_221
timestamp 1607101874
transform 1 0 2052 0 -1 4305
box -2 -3 18 103
use AOI21X1  AOI21X1_248
timestamp 1607101874
transform 1 0 2068 0 -1 4305
box -2 -3 34 103
use BUFX4  BUFX4_437
timestamp 1607101874
transform 1 0 2100 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_338
timestamp 1607101874
transform 1 0 2132 0 -1 4305
box -2 -3 50 103
use NAND3X1  NAND3X1_71
timestamp 1607101874
transform -1 0 2212 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_369
timestamp 1607101874
transform -1 0 2228 0 -1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1607101874
transform 1 0 2228 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1108
timestamp 1607101874
transform 1 0 2324 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1109
timestamp 1607101874
transform 1 0 2356 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_4_0
timestamp 1607101874
transform -1 0 2396 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_4_1
timestamp 1607101874
transform -1 0 2404 0 -1 4305
box -2 -3 10 103
use AOI21X1  AOI21X1_473
timestamp 1607101874
transform -1 0 2436 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_334
timestamp 1607101874
transform -1 0 2460 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1211
timestamp 1607101874
transform 1 0 2460 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1607101874
transform 1 0 2492 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_693
timestamp 1607101874
transform -1 0 2548 0 -1 4305
box -2 -3 34 103
use AND2X2  AND2X2_33
timestamp 1607101874
transform -1 0 2580 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_932
timestamp 1607101874
transform -1 0 2676 0 -1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1607101874
transform 1 0 2676 0 -1 4305
box -2 -3 98 103
use AOI21X1  AOI21X1_260
timestamp 1607101874
transform 1 0 2772 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1423
timestamp 1607101874
transform 1 0 2804 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1422
timestamp 1607101874
transform -1 0 2868 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_234
timestamp 1607101874
transform 1 0 2868 0 -1 4305
box -2 -3 18 103
use FILL  FILL_42_5_0
timestamp 1607101874
transform 1 0 2884 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_5_1
timestamp 1607101874
transform 1 0 2892 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_572
timestamp 1607101874
transform 1 0 2900 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1607101874
transform -1 0 2964 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_237
timestamp 1607101874
transform -1 0 2980 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_231
timestamp 1607101874
transform 1 0 2980 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1607101874
transform 1 0 3012 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_918
timestamp 1607101874
transform 1 0 3044 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_442
timestamp 1607101874
transform 1 0 3140 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_1210
timestamp 1607101874
transform 1 0 3156 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_500
timestamp 1607101874
transform -1 0 3220 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_176
timestamp 1607101874
transform 1 0 3220 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_108
timestamp 1607101874
transform -1 0 3276 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_459
timestamp 1607101874
transform 1 0 3276 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_260
timestamp 1607101874
transform 1 0 3372 0 -1 4305
box -2 -3 18 103
use FILL  FILL_42_6_0
timestamp 1607101874
transform -1 0 3396 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_6_1
timestamp 1607101874
transform -1 0 3404 0 -1 4305
box -2 -3 10 103
use MUX2X1  MUX2X1_365
timestamp 1607101874
transform -1 0 3452 0 -1 4305
box -2 -3 50 103
use MUX2X1  MUX2X1_264
timestamp 1607101874
transform -1 0 3500 0 -1 4305
box -2 -3 50 103
use BUFX4  BUFX4_210
timestamp 1607101874
transform -1 0 3532 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_191
timestamp 1607101874
transform 1 0 3532 0 -1 4305
box -2 -3 26 103
use BUFX4  BUFX4_61
timestamp 1607101874
transform 1 0 3556 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1250
timestamp 1607101874
transform 1 0 3588 0 -1 4305
box -2 -3 34 103
use OAI22X1  OAI22X1_89
timestamp 1607101874
transform -1 0 3660 0 -1 4305
box -2 -3 42 103
use BUFX4  BUFX4_431
timestamp 1607101874
transform -1 0 3692 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1461
timestamp 1607101874
transform 1 0 3692 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1462
timestamp 1607101874
transform 1 0 3724 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1449
timestamp 1607101874
transform 1 0 3756 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1448
timestamp 1607101874
transform 1 0 3788 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1064
timestamp 1607101874
transform -1 0 3852 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_291
timestamp 1607101874
transform 1 0 3852 0 -1 4305
box -2 -3 98 103
use FILL  FILL_42_7_0
timestamp 1607101874
transform -1 0 3956 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_7_1
timestamp 1607101874
transform -1 0 3964 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_942
timestamp 1607101874
transform -1 0 4060 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_126
timestamp 1607101874
transform 1 0 4060 0 -1 4305
box -2 -3 18 103
use MUX2X1  MUX2X1_113
timestamp 1607101874
transform -1 0 4124 0 -1 4305
box -2 -3 50 103
use BUFX4  BUFX4_60
timestamp 1607101874
transform -1 0 4156 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1157
timestamp 1607101874
transform 1 0 4156 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_774
timestamp 1607101874
transform -1 0 4220 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_903
timestamp 1607101874
transform -1 0 4252 0 -1 4305
box -2 -3 34 103
use OAI22X1  OAI22X1_34
timestamp 1607101874
transform 1 0 4252 0 -1 4305
box -2 -3 42 103
use NOR2X1  NOR2X1_466
timestamp 1607101874
transform -1 0 4316 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_429
timestamp 1607101874
transform -1 0 4340 0 -1 4305
box -2 -3 26 103
use OAI22X1  OAI22X1_22
timestamp 1607101874
transform 1 0 4340 0 -1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_776
timestamp 1607101874
transform -1 0 4412 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_428
timestamp 1607101874
transform 1 0 4412 0 -1 4305
box -2 -3 26 103
use FILL  FILL_42_8_0
timestamp 1607101874
transform -1 0 4444 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_8_1
timestamp 1607101874
transform -1 0 4452 0 -1 4305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_50
timestamp 1607101874
transform -1 0 4524 0 -1 4305
box -2 -3 74 103
use NOR2X1  NOR2X1_613
timestamp 1607101874
transform 1 0 4524 0 -1 4305
box -2 -3 26 103
use OAI22X1  OAI22X1_87
timestamp 1607101874
transform 1 0 4548 0 -1 4305
box -2 -3 42 103
use AOI21X1  AOI21X1_596
timestamp 1607101874
transform 1 0 4588 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_708
timestamp 1607101874
transform 1 0 4620 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_476
timestamp 1607101874
transform -1 0 4740 0 -1 4305
box -2 -3 98 103
use MUX2X1  MUX2X1_55
timestamp 1607101874
transform 1 0 4740 0 -1 4305
box -2 -3 50 103
use INVX1  INVX1_65
timestamp 1607101874
transform 1 0 4788 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_955
timestamp 1607101874
transform -1 0 4836 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_612
timestamp 1607101874
transform -1 0 4860 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_974
timestamp 1607101874
transform -1 0 4956 0 -1 4305
box -2 -3 98 103
use FILL  FILL_42_9_0
timestamp 1607101874
transform 1 0 4956 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_9_1
timestamp 1607101874
transform 1 0 4964 0 -1 4305
box -2 -3 10 103
use NOR2X1  NOR2X1_204
timestamp 1607101874
transform 1 0 4972 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_127
timestamp 1607101874
transform -1 0 5028 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_991
timestamp 1607101874
transform -1 0 5060 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_495
timestamp 1607101874
transform -1 0 5084 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_42
timestamp 1607101874
transform 1 0 5084 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1607101874
transform -1 0 5140 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_990
timestamp 1607101874
transform 1 0 5140 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1607101874
transform 1 0 5172 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_661
timestamp 1607101874
transform -1 0 5300 0 -1 4305
box -2 -3 98 103
use FILL  FILL_43_1
timestamp 1607101874
transform -1 0 5308 0 -1 4305
box -2 -3 10 103
use NAND2X1  NAND2X1_121
timestamp 1607101874
transform -1 0 28 0 1 4305
box -2 -3 26 103
use INVX2  INVX2_23
timestamp 1607101874
transform 1 0 28 0 1 4305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_2
timestamp 1607101874
transform -1 0 100 0 1 4305
box -2 -3 58 103
use NAND2X1  NAND2X1_138
timestamp 1607101874
transform 1 0 100 0 1 4305
box -2 -3 26 103
use AND2X2  AND2X2_9
timestamp 1607101874
transform 1 0 124 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_342
timestamp 1607101874
transform 1 0 156 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_157
timestamp 1607101874
transform 1 0 180 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_226
timestamp 1607101874
transform 1 0 204 0 1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_40
timestamp 1607101874
transform 1 0 236 0 1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1607101874
transform 1 0 268 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1607101874
transform 1 0 300 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_0_0
timestamp 1607101874
transform -1 0 332 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_0_1
timestamp 1607101874
transform -1 0 340 0 1 4305
box -2 -3 10 103
use AOI22X1  AOI22X1_7
timestamp 1607101874
transform -1 0 380 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_520
timestamp 1607101874
transform -1 0 412 0 1 4305
box -2 -3 34 103
use XOR2X1  XOR2X1_3
timestamp 1607101874
transform 1 0 412 0 1 4305
box -2 -3 58 103
use NOR2X1  NOR2X1_337
timestamp 1607101874
transform -1 0 492 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_483
timestamp 1607101874
transform -1 0 524 0 1 4305
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1607101874
transform -1 0 540 0 1 4305
box -2 -3 18 103
use NOR2X1  NOR2X1_319
timestamp 1607101874
transform 1 0 540 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_165
timestamp 1607101874
transform 1 0 564 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_541
timestamp 1607101874
transform 1 0 588 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_352
timestamp 1607101874
transform 1 0 620 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_542
timestamp 1607101874
transform -1 0 676 0 1 4305
box -2 -3 34 103
use INVX4  INVX4_6
timestamp 1607101874
transform 1 0 676 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_353
timestamp 1607101874
transform -1 0 724 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_543
timestamp 1607101874
transform 1 0 724 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_307
timestamp 1607101874
transform -1 0 788 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_470
timestamp 1607101874
transform -1 0 820 0 1 4305
box -2 -3 34 103
use INVX2  INVX2_13
timestamp 1607101874
transform 1 0 820 0 1 4305
box -2 -3 18 103
use FILL  FILL_43_1_0
timestamp 1607101874
transform -1 0 844 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_1_1
timestamp 1607101874
transform -1 0 852 0 1 4305
box -2 -3 10 103
use NOR3X1  NOR3X1_7
timestamp 1607101874
transform -1 0 916 0 1 4305
box -2 -3 66 103
use NAND3X1  NAND3X1_29
timestamp 1607101874
transform -1 0 948 0 1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1607101874
transform 1 0 948 0 1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_205
timestamp 1607101874
transform -1 0 1012 0 1 4305
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1607101874
transform 1 0 1012 0 1 4305
box -2 -3 66 103
use NAND2X1  NAND2X1_169
timestamp 1607101874
transform -1 0 1100 0 1 4305
box -2 -3 26 103
use NAND3X1  NAND3X1_13
timestamp 1607101874
transform -1 0 1132 0 1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1607101874
transform 1 0 1132 0 1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_69
timestamp 1607101874
transform -1 0 1196 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1607101874
transform -1 0 1220 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_544
timestamp 1607101874
transform -1 0 1252 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_217
timestamp 1607101874
transform -1 0 1268 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_413
timestamp 1607101874
transform 1 0 1268 0 1 4305
box -2 -3 98 103
use FILL  FILL_43_2_0
timestamp 1607101874
transform 1 0 1364 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_2_1
timestamp 1607101874
transform 1 0 1372 0 1 4305
box -2 -3 10 103
use AOI21X1  AOI21X1_577
timestamp 1607101874
transform 1 0 1380 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_689
timestamp 1607101874
transform -1 0 1436 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1607101874
transform -1 0 1532 0 1 4305
box -2 -3 98 103
use AOI21X1  AOI21X1_263
timestamp 1607101874
transform 1 0 1532 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_581
timestamp 1607101874
transform 1 0 1564 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1421
timestamp 1607101874
transform 1 0 1596 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_417
timestamp 1607101874
transform 1 0 1628 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1420
timestamp 1607101874
transform -1 0 1756 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_414
timestamp 1607101874
transform 1 0 1756 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_223
timestamp 1607101874
transform -1 0 1884 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_3_0
timestamp 1607101874
transform 1 0 1884 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_3_1
timestamp 1607101874
transform 1 0 1892 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_217
timestamp 1607101874
transform 1 0 1900 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_216
timestamp 1607101874
transform 1 0 1932 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_902
timestamp 1607101874
transform 1 0 1964 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_913
timestamp 1607101874
transform 1 0 2060 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_553
timestamp 1607101874
transform -1 0 2188 0 1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_101
timestamp 1607101874
transform -1 0 2236 0 1 4305
box -2 -3 50 103
use INVX1  INVX1_114
timestamp 1607101874
transform 1 0 2236 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_406
timestamp 1607101874
transform 1 0 2252 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_236
timestamp 1607101874
transform 1 0 2348 0 1 4305
box -2 -3 18 103
use FILL  FILL_43_4_0
timestamp 1607101874
transform -1 0 2372 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_4_1
timestamp 1607101874
transform -1 0 2380 0 1 4305
box -2 -3 10 103
use MUX2X1  MUX2X1_342
timestamp 1607101874
transform -1 0 2428 0 1 4305
box -2 -3 50 103
use AOI21X1  AOI21X1_472
timestamp 1607101874
transform -1 0 2460 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_853
timestamp 1607101874
transform -1 0 2492 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_573
timestamp 1607101874
transform -1 0 2524 0 1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_103
timestamp 1607101874
transform -1 0 2572 0 1 4305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1607101874
transform -1 0 2668 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1428
timestamp 1607101874
transform -1 0 2700 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1429
timestamp 1607101874
transform -1 0 2732 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_574
timestamp 1607101874
transform 1 0 2732 0 1 4305
box -2 -3 34 103
use OAI22X1  OAI22X1_4
timestamp 1607101874
transform -1 0 2804 0 1 4305
box -2 -3 42 103
use AOI21X1  AOI21X1_261
timestamp 1607101874
transform 1 0 2804 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_151
timestamp 1607101874
transform 1 0 2836 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_5_0
timestamp 1607101874
transform 1 0 2868 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_5_1
timestamp 1607101874
transform 1 0 2876 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1607101874
transform 1 0 2884 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_110
timestamp 1607101874
transform 1 0 2980 0 1 4305
box -2 -3 18 103
use MUX2X1  MUX2X1_97
timestamp 1607101874
transform -1 0 3044 0 1 4305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_907
timestamp 1607101874
transform 1 0 3044 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_669
timestamp 1607101874
transform 1 0 3140 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_922
timestamp 1607101874
transform -1 0 3268 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_290
timestamp 1607101874
transform -1 0 3364 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1446
timestamp 1607101874
transform -1 0 3396 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_6_0
timestamp 1607101874
transform -1 0 3404 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_6_1
timestamp 1607101874
transform -1 0 3412 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_1447
timestamp 1607101874
transform -1 0 3444 0 1 4305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_83
timestamp 1607101874
transform -1 0 3516 0 1 4305
box -2 -3 74 103
use OAI21X1  OAI21X1_255
timestamp 1607101874
transform 1 0 3516 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_254
timestamp 1607101874
transform 1 0 3548 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_950
timestamp 1607101874
transform -1 0 3676 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_293
timestamp 1607101874
transform 1 0 3676 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1453
timestamp 1607101874
transform 1 0 3772 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1452
timestamp 1607101874
transform 1 0 3804 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_433
timestamp 1607101874
transform 1 0 3836 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_327
timestamp 1607101874
transform 1 0 3868 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_617
timestamp 1607101874
transform -1 0 3916 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_7_0
timestamp 1607101874
transform 1 0 3916 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_7_1
timestamp 1607101874
transform 1 0 3924 0 1 4305
box -2 -3 10 103
use MUX2X1  MUX2X1_299
timestamp 1607101874
transform 1 0 3932 0 1 4305
box -2 -3 50 103
use OAI21X1  OAI21X1_941
timestamp 1607101874
transform -1 0 4012 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_940
timestamp 1607101874
transform 1 0 4012 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_478
timestamp 1607101874
transform 1 0 4044 0 1 4305
box -2 -3 26 103
use MUX2X1  MUX2X1_296
timestamp 1607101874
transform 1 0 4068 0 1 4305
box -2 -3 50 103
use INVX1  INVX1_367
timestamp 1607101874
transform -1 0 4132 0 1 4305
box -2 -3 18 103
use MUX2X1  MUX2X1_358
timestamp 1607101874
transform 1 0 4132 0 1 4305
box -2 -3 50 103
use NAND2X1  NAND2X1_239
timestamp 1607101874
transform 1 0 4180 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_599
timestamp 1607101874
transform 1 0 4204 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_711
timestamp 1607101874
transform -1 0 4260 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_468
timestamp 1607101874
transform 1 0 4260 0 1 4305
box -2 -3 98 103
use NOR2X1  NOR2X1_211
timestamp 1607101874
transform 1 0 4356 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_132
timestamp 1607101874
transform -1 0 4412 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_8_0
timestamp 1607101874
transform -1 0 4420 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_8_1
timestamp 1607101874
transform -1 0 4428 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_980
timestamp 1607101874
transform -1 0 4524 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_464
timestamp 1607101874
transform -1 0 4620 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1102
timestamp 1607101874
transform 1 0 4620 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_713
timestamp 1607101874
transform 1 0 4652 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_601
timestamp 1607101874
transform -1 0 4708 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_156
timestamp 1607101874
transform 1 0 4708 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_956
timestamp 1607101874
transform 1 0 4740 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_755
timestamp 1607101874
transform -1 0 4868 0 1 4305
box -2 -3 98 103
use MUX2X1  MUX2X1_373
timestamp 1607101874
transform 1 0 4868 0 1 4305
box -2 -3 50 103
use INVX1  INVX1_378
timestamp 1607101874
transform -1 0 4932 0 1 4305
box -2 -3 18 103
use FILL  FILL_43_9_0
timestamp 1607101874
transform -1 0 4940 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_9_1
timestamp 1607101874
transform -1 0 4948 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_473
timestamp 1607101874
transform -1 0 5044 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_872
timestamp 1607101874
transform -1 0 5076 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_669
timestamp 1607101874
transform -1 0 5172 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_396
timestamp 1607101874
transform -1 0 5204 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1607101874
transform 1 0 5204 0 1 4305
box -2 -3 98 103
use FILL  FILL_44_1
timestamp 1607101874
transform 1 0 5300 0 1 4305
box -2 -3 10 103
use NAND2X1  NAND2X1_122
timestamp 1607101874
transform 1 0 4 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_486
timestamp 1607101874
transform 1 0 28 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_336
timestamp 1607101874
transform 1 0 60 0 -1 4505
box -2 -3 26 103
use NAND3X1  NAND3X1_62
timestamp 1607101874
transform 1 0 84 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_242
timestamp 1607101874
transform 1 0 116 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_243
timestamp 1607101874
transform -1 0 180 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_199
timestamp 1607101874
transform 1 0 180 0 -1 4505
box -2 -3 18 103
use NOR3X1  NOR3X1_13
timestamp 1607101874
transform 1 0 196 0 -1 4505
box -2 -3 66 103
use OAI21X1  OAI21X1_492
timestamp 1607101874
transform -1 0 292 0 -1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_54
timestamp 1607101874
transform -1 0 324 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_0_0
timestamp 1607101874
transform -1 0 332 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_0_1
timestamp 1607101874
transform -1 0 340 0 -1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_241
timestamp 1607101874
transform -1 0 372 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_323
timestamp 1607101874
transform -1 0 396 0 -1 4505
box -2 -3 26 103
use NAND3X1  NAND3X1_64
timestamp 1607101874
transform -1 0 428 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_227
timestamp 1607101874
transform 1 0 428 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1607101874
transform -1 0 492 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_328
timestamp 1607101874
transform -1 0 516 0 -1 4505
box -2 -3 26 103
use NAND3X1  NAND3X1_39
timestamp 1607101874
transform 1 0 516 0 -1 4505
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1607101874
transform -1 0 588 0 -1 4505
box -2 -3 42 103
use NOR2X1  NOR2X1_327
timestamp 1607101874
transform 1 0 588 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_490
timestamp 1607101874
transform -1 0 644 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_480
timestamp 1607101874
transform -1 0 676 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_129
timestamp 1607101874
transform -1 0 700 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_478
timestamp 1607101874
transform -1 0 732 0 -1 4505
box -2 -3 34 103
use NOR3X1  NOR3X1_10
timestamp 1607101874
transform -1 0 796 0 -1 4505
box -2 -3 66 103
use AOI22X1  AOI22X1_9
timestamp 1607101874
transform 1 0 796 0 -1 4505
box -2 -3 42 103
use FILL  FILL_44_1_0
timestamp 1607101874
transform -1 0 844 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_1_1
timestamp 1607101874
transform -1 0 852 0 -1 4505
box -2 -3 10 103
use NAND3X1  NAND3X1_66
timestamp 1607101874
transform -1 0 884 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_533
timestamp 1607101874
transform 1 0 884 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_347
timestamp 1607101874
transform -1 0 940 0 -1 4505
box -2 -3 26 103
use NAND3X1  NAND3X1_35
timestamp 1607101874
transform 1 0 940 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_219
timestamp 1607101874
transform -1 0 1004 0 -1 4505
box -2 -3 34 103
use NOR3X1  NOR3X1_8
timestamp 1607101874
transform -1 0 1068 0 -1 4505
box -2 -3 66 103
use AOI21X1  AOI21X1_217
timestamp 1607101874
transform -1 0 1100 0 -1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1607101874
transform 1 0 1100 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_218
timestamp 1607101874
transform -1 0 1164 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_140
timestamp 1607101874
transform -1 0 1188 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_446
timestamp 1607101874
transform -1 0 1220 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_99
timestamp 1607101874
transform -1 0 1244 0 -1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_302
timestamp 1607101874
transform 1 0 1244 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_202
timestamp 1607101874
transform -1 0 1300 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_357
timestamp 1607101874
transform -1 0 1324 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_206
timestamp 1607101874
transform -1 0 1356 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_2_0
timestamp 1607101874
transform -1 0 1364 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_2_1
timestamp 1607101874
transform -1 0 1372 0 -1 4505
box -2 -3 10 103
use NAND2X1  NAND2X1_101
timestamp 1607101874
transform -1 0 1396 0 -1 4505
box -2 -3 26 103
use INVX8  INVX8_11
timestamp 1607101874
transform 1 0 1396 0 -1 4505
box -2 -3 42 103
use AOI21X1  AOI21X1_99
timestamp 1607101874
transform 1 0 1436 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1607101874
transform -1 0 1492 0 -1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_903
timestamp 1607101874
transform 1 0 1492 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1113
timestamp 1607101874
transform -1 0 1620 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_102
timestamp 1607101874
transform 1 0 1620 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_167
timestamp 1607101874
transform -1 0 1676 0 -1 4505
box -2 -3 26 103
use BUFX4  BUFX4_208
timestamp 1607101874
transform -1 0 1708 0 -1 4505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1607101874
transform -1 0 1780 0 -1 4505
box -2 -3 74 103
use NAND2X1  NAND2X1_217
timestamp 1607101874
transform 1 0 1780 0 -1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_162
timestamp 1607101874
transform 1 0 1804 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_98
timestamp 1607101874
transform -1 0 1860 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_3_0
timestamp 1607101874
transform 1 0 1860 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_3_1
timestamp 1607101874
transform 1 0 1868 0 -1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_899
timestamp 1607101874
transform 1 0 1876 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_286
timestamp 1607101874
transform 1 0 1972 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_690
timestamp 1607101874
transform 1 0 1988 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_218
timestamp 1607101874
transform 1 0 2020 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_691
timestamp 1607101874
transform -1 0 2076 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_340
timestamp 1607101874
transform 1 0 2076 0 -1 4505
box -2 -3 50 103
use INVX1  INVX1_240
timestamp 1607101874
transform -1 0 2140 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1607101874
transform -1 0 2236 0 -1 4505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_29
timestamp 1607101874
transform 1 0 2236 0 -1 4505
box -2 -3 74 103
use INVX1  INVX1_420
timestamp 1607101874
transform 1 0 2308 0 -1 4505
box -2 -3 18 103
use MUX2X1  MUX2X1_345
timestamp 1607101874
transform -1 0 2372 0 -1 4505
box -2 -3 50 103
use NOR2X1  NOR2X1_83
timestamp 1607101874
transform 1 0 2372 0 -1 4505
box -2 -3 26 103
use FILL  FILL_44_4_0
timestamp 1607101874
transform 1 0 2396 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_4_1
timestamp 1607101874
transform 1 0 2404 0 -1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_499
timestamp 1607101874
transform 1 0 2412 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1209
timestamp 1607101874
transform -1 0 2476 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_116
timestamp 1607101874
transform -1 0 2492 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_923
timestamp 1607101874
transform -1 0 2588 0 -1 4505
box -2 -3 98 103
use MUX2X1  MUX2X1_104
timestamp 1607101874
transform 1 0 2588 0 -1 4505
box -2 -3 50 103
use INVX1  INVX1_117
timestamp 1607101874
transform -1 0 2652 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_851
timestamp 1607101874
transform 1 0 2652 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_399
timestamp 1607101874
transform -1 0 2708 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_463
timestamp 1607101874
transform 1 0 2708 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_577
timestamp 1607101874
transform 1 0 2740 0 -1 4505
box -2 -3 34 103
use AND2X2  AND2X2_29
timestamp 1607101874
transform -1 0 2804 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1086
timestamp 1607101874
transform -1 0 2836 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_284
timestamp 1607101874
transform 1 0 2836 0 -1 4505
box -2 -3 50 103
use INVX1  INVX1_411
timestamp 1607101874
transform -1 0 2900 0 -1 4505
box -2 -3 18 103
use FILL  FILL_44_5_0
timestamp 1607101874
transform -1 0 2908 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_5_1
timestamp 1607101874
transform -1 0 2916 0 -1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_381
timestamp 1607101874
transform -1 0 3012 0 -1 4505
box -2 -3 98 103
use MUX2X1  MUX2X1_303
timestamp 1607101874
transform -1 0 3060 0 -1 4505
box -2 -3 50 103
use NOR2X1  NOR2X1_388
timestamp 1607101874
transform 1 0 3060 0 -1 4505
box -2 -3 26 103
use INVX1  INVX1_366
timestamp 1607101874
transform -1 0 3100 0 -1 4505
box -2 -3 18 103
use AOI21X1  AOI21X1_303
timestamp 1607101874
transform -1 0 3132 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_389
timestamp 1607101874
transform -1 0 3156 0 -1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_211
timestamp 1607101874
transform 1 0 3156 0 -1 4505
box -2 -3 26 103
use OAI22X1  OAI22X1_11
timestamp 1607101874
transform 1 0 3180 0 -1 4505
box -2 -3 42 103
use OAI21X1  OAI21X1_668
timestamp 1607101874
transform -1 0 3252 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_947
timestamp 1607101874
transform -1 0 3348 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_248
timestamp 1607101874
transform -1 0 3380 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_249
timestamp 1607101874
transform -1 0 3412 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 4505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_10
timestamp 1607101874
transform 1 0 3428 0 -1 4505
box -2 -3 74 103
use BUFX4  BUFX4_434
timestamp 1607101874
transform 1 0 3500 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_117
timestamp 1607101874
transform 1 0 3532 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_190
timestamp 1607101874
transform -1 0 3588 0 -1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_954
timestamp 1607101874
transform 1 0 3588 0 -1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_618
timestamp 1607101874
transform 1 0 3684 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_116
timestamp 1607101874
transform 1 0 3708 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_953
timestamp 1607101874
transform -1 0 3836 0 -1 4505
box -2 -3 98 103
use AOI21X1  AOI21X1_454
timestamp 1607101874
transform 1 0 3836 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1063
timestamp 1607101874
transform 1 0 3868 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_7_0
timestamp 1607101874
transform 1 0 3900 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_7_1
timestamp 1607101874
transform 1 0 3908 0 -1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_368
timestamp 1607101874
transform 1 0 3916 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_368
timestamp 1607101874
transform 1 0 4012 0 -1 4505
box -2 -3 18 103
use BUFX4  BUFX4_340
timestamp 1607101874
transform 1 0 4028 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_211
timestamp 1607101874
transform -1 0 4108 0 -1 4505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1607101874
transform -1 0 4204 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_317
timestamp 1607101874
transform -1 0 4220 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_275
timestamp 1607101874
transform -1 0 4316 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_772
timestamp 1607101874
transform 1 0 4316 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_362
timestamp 1607101874
transform 1 0 4348 0 -1 4505
box -2 -3 50 103
use OAI21X1  OAI21X1_596
timestamp 1607101874
transform 1 0 4396 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_8_0
timestamp 1607101874
transform -1 0 4436 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_8_1
timestamp 1607101874
transform -1 0 4444 0 -1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_274
timestamp 1607101874
transform -1 0 4476 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_707
timestamp 1607101874
transform 1 0 4476 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_595
timestamp 1607101874
transform -1 0 4532 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_463
timestamp 1607101874
transform -1 0 4628 0 -1 4505
box -2 -3 98 103
use BUFX4  BUFX4_215
timestamp 1607101874
transform 1 0 4628 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1100
timestamp 1607101874
transform -1 0 4692 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_373
timestamp 1607101874
transform -1 0 4788 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_954
timestamp 1607101874
transform 1 0 4788 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_376
timestamp 1607101874
transform -1 0 4836 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_1194
timestamp 1607101874
transform -1 0 4868 0 -1 4505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_1
timestamp 1607101874
transform -1 0 4940 0 -1 4505
box -2 -3 74 103
use FILL  FILL_44_9_0
timestamp 1607101874
transform -1 0 4948 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_9_1
timestamp 1607101874
transform -1 0 4956 0 -1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_415
timestamp 1607101874
transform -1 0 4988 0 -1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_597
timestamp 1607101874
transform -1 0 5020 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_465
timestamp 1607101874
transform -1 0 5116 0 -1 4505
box -2 -3 98 103
use AOI21X1  AOI21X1_16
timestamp 1607101874
transform 1 0 5116 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_27
timestamp 1607101874
transform 1 0 5148 0 -1 4505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_664
timestamp 1607101874
transform -1 0 5292 0 -1 4505
box -2 -3 98 103
use FILL  FILL_45_1
timestamp 1607101874
transform -1 0 5300 0 -1 4505
box -2 -3 10 103
use FILL  FILL_45_2
timestamp 1607101874
transform -1 0 5308 0 -1 4505
box -2 -3 10 103
use INVX4  INVX4_10
timestamp 1607101874
transform -1 0 28 0 1 4505
box -2 -3 26 103
use INVX4  INVX4_12
timestamp 1607101874
transform -1 0 52 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_155
timestamp 1607101874
transform -1 0 76 0 1 4505
box -2 -3 26 103
use NAND3X1  NAND3X1_63
timestamp 1607101874
transform -1 0 108 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_404
timestamp 1607101874
transform 1 0 4 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_528
timestamp 1607101874
transform -1 0 132 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_527
timestamp 1607101874
transform -1 0 140 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_524
timestamp 1607101874
transform 1 0 140 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1607101874
transform -1 0 204 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_44
timestamp 1607101874
transform 1 0 204 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_338
timestamp 1607101874
transform 1 0 132 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_191
timestamp 1607101874
transform 1 0 156 0 -1 4705
box -2 -3 18 103
use NAND2X1  NAND2X1_116
timestamp 1607101874
transform -1 0 196 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_188
timestamp 1607101874
transform 1 0 196 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_493
timestamp 1607101874
transform 1 0 236 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_513
timestamp 1607101874
transform 1 0 268 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1607101874
transform -1 0 332 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1607101874
transform 1 0 212 0 -1 4705
box -2 -3 26 103
use NAND2X1  NAND2X1_137
timestamp 1607101874
transform -1 0 260 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_484
timestamp 1607101874
transform -1 0 292 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_0_0
timestamp 1607101874
transform 1 0 292 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_0_1
timestamp 1607101874
transform 1 0 300 0 -1 4705
box -2 -3 10 103
use FILL  FILL_45_0_0
timestamp 1607101874
transform -1 0 340 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_0_1
timestamp 1607101874
transform -1 0 348 0 1 4505
box -2 -3 10 103
use NOR2X1  NOR2X1_335
timestamp 1607101874
transform -1 0 372 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_225
timestamp 1607101874
transform 1 0 372 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_341
timestamp 1607101874
transform -1 0 428 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_403
timestamp 1607101874
transform 1 0 308 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_321
timestamp 1607101874
transform -1 0 428 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_198
timestamp 1607101874
transform -1 0 444 0 1 4505
box -2 -3 18 103
use NOR2X1  NOR2X1_340
timestamp 1607101874
transform -1 0 468 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_134
timestamp 1607101874
transform -1 0 492 0 1 4505
box -2 -3 26 103
use INVX2  INVX2_22
timestamp 1607101874
transform -1 0 508 0 1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_482
timestamp 1607101874
transform -1 0 540 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_322
timestamp 1607101874
transform 1 0 428 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_197
timestamp 1607101874
transform -1 0 468 0 -1 4705
box -2 -3 18 103
use NAND2X1  NAND2X1_133
timestamp 1607101874
transform -1 0 492 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_401
timestamp 1607101874
transform 1 0 492 0 -1 4705
box -2 -3 98 103
use OAI22X1  OAI22X1_1
timestamp 1607101874
transform 1 0 540 0 1 4505
box -2 -3 42 103
use NAND3X1  NAND3X1_41
timestamp 1607101874
transform -1 0 612 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_145
timestamp 1607101874
transform -1 0 612 0 -1 4705
box -2 -3 26 103
use NAND2X1  NAND2X1_128
timestamp 1607101874
transform 1 0 612 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_314
timestamp 1607101874
transform -1 0 660 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_313
timestamp 1607101874
transform 1 0 660 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_312
timestamp 1607101874
transform -1 0 708 0 1 4505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_6
timestamp 1607101874
transform 1 0 708 0 1 4505
box -2 -3 58 103
use NAND3X1  NAND3X1_33
timestamp 1607101874
transform 1 0 612 0 -1 4705
box -2 -3 34 103
use NAND3X1  NAND3X1_42
timestamp 1607101874
transform 1 0 644 0 -1 4705
box -2 -3 34 103
use NAND3X1  NAND3X1_43
timestamp 1607101874
transform 1 0 676 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_320
timestamp 1607101874
transform 1 0 708 0 -1 4705
box -2 -3 26 103
use NOR2X1  NOR2X1_344
timestamp 1607101874
transform -1 0 788 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_346
timestamp 1607101874
transform 1 0 788 0 1 4505
box -2 -3 26 103
use BUFX4  BUFX4_305
timestamp 1607101874
transform -1 0 764 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_534
timestamp 1607101874
transform 1 0 764 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_536
timestamp 1607101874
transform 1 0 796 0 -1 4705
box -2 -3 34 103
use NOR3X1  NOR3X1_9
timestamp 1607101874
transform 1 0 812 0 1 4505
box -2 -3 66 103
use FILL  FILL_45_1_0
timestamp 1607101874
transform 1 0 876 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_1_1
timestamp 1607101874
transform 1 0 884 0 1 4505
box -2 -3 10 103
use OAI21X1  OAI21X1_467
timestamp 1607101874
transform 1 0 892 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_535
timestamp 1607101874
transform 1 0 828 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_1_0
timestamp 1607101874
transform -1 0 868 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_1_1
timestamp 1607101874
transform -1 0 876 0 -1 4705
box -2 -3 10 103
use AOI21X1  AOI21X1_244
timestamp 1607101874
transform -1 0 908 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_537
timestamp 1607101874
transform 1 0 908 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_125
timestamp 1607101874
transform 1 0 924 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_216
timestamp 1607101874
transform 1 0 948 0 1 4505
box -2 -3 34 103
use NOR3X1  NOR3X1_3
timestamp 1607101874
transform -1 0 1044 0 1 4505
box -2 -3 66 103
use AOI21X1  AOI21X1_245
timestamp 1607101874
transform 1 0 940 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_468
timestamp 1607101874
transform -1 0 1004 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1607101874
transform -1 0 1028 0 -1 4705
box -2 -3 26 103
use NAND2X1  NAND2X1_105
timestamp 1607101874
transform -1 0 1068 0 1 4505
box -2 -3 26 103
use OR2X2  OR2X2_2
timestamp 1607101874
transform 1 0 1068 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1607101874
transform -1 0 1132 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1607101874
transform 1 0 1028 0 -1 4705
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1607101874
transform 1 0 1060 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_187
timestamp 1607101874
transform -1 0 1108 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_440
timestamp 1607101874
transform -1 0 1140 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1607101874
transform 1 0 1132 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_447
timestamp 1607101874
transform -1 0 1188 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_444
timestamp 1607101874
transform -1 0 1220 0 1 4505
box -2 -3 34 103
use INVX2  INVX2_26
timestamp 1607101874
transform -1 0 1156 0 -1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_345
timestamp 1607101874
transform -1 0 1180 0 -1 4705
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1607101874
transform -1 0 1212 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_445
timestamp 1607101874
transform -1 0 1244 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1607101874
transform -1 0 1244 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_299
timestamp 1607101874
transform 1 0 1244 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_438
timestamp 1607101874
transform 1 0 1268 0 1 4505
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1607101874
transform -1 0 1332 0 1 4505
box -2 -3 34 103
use AOI22X1  AOI22X1_1
timestamp 1607101874
transform 1 0 1244 0 -1 4705
box -2 -3 42 103
use OAI21X1  OAI21X1_532
timestamp 1607101874
transform -1 0 1316 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_354
timestamp 1607101874
transform -1 0 1340 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_216
timestamp 1607101874
transform 1 0 1340 0 -1 4705
box -2 -3 18 103
use AND2X2  AND2X2_1
timestamp 1607101874
transform -1 0 1364 0 1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_203
timestamp 1607101874
transform -1 0 1404 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_2_1
timestamp 1607101874
transform -1 0 1372 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_2_0
timestamp 1607101874
transform -1 0 1364 0 -1 4705
box -2 -3 10 103
use AOI21X1  AOI21X1_204
timestamp 1607101874
transform -1 0 1412 0 1 4505
box -2 -3 34 103
use FILL  FILL_45_2_1
timestamp 1607101874
transform -1 0 1380 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_2_0
timestamp 1607101874
transform -1 0 1372 0 1 4505
box -2 -3 10 103
use NAND3X1  NAND3X1_5
timestamp 1607101874
transform 1 0 1404 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_100
timestamp 1607101874
transform -1 0 1436 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_439
timestamp 1607101874
transform -1 0 1468 0 1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_275
timestamp 1607101874
transform 1 0 1468 0 1 4505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1607101874
transform 1 0 1516 0 1 4505
box -2 -3 98 103
use OR2X2  OR2X2_1
timestamp 1607101874
transform -1 0 1468 0 -1 4705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_45
timestamp 1607101874
transform -1 0 1540 0 -1 4705
box -2 -3 74 103
use INVX1  INVX1_220
timestamp 1607101874
transform 1 0 1612 0 1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1607101874
transform 1 0 1540 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_906
timestamp 1607101874
transform 1 0 1628 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_242
timestamp 1607101874
transform 1 0 1636 0 -1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_880
timestamp 1607101874
transform 1 0 1652 0 -1 4705
box -2 -3 98 103
use BUFX4  BUFX4_474
timestamp 1607101874
transform 1 0 1724 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1607101874
transform 1 0 1756 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1206
timestamp 1607101874
transform -1 0 1812 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_898
timestamp 1607101874
transform -1 0 1908 0 1 4505
box -2 -3 98 103
use AOI21X1  AOI21X1_91
timestamp 1607101874
transform 1 0 1748 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_154
timestamp 1607101874
transform -1 0 1804 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_879
timestamp 1607101874
transform 1 0 1804 0 -1 4705
box -2 -3 98 103
use FILL  FILL_45_3_0
timestamp 1607101874
transform 1 0 1908 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_3_1
timestamp 1607101874
transform 1 0 1916 0 1 4505
box -2 -3 10 103
use FILL  FILL_46_3_0
timestamp 1607101874
transform 1 0 1900 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_3_1
timestamp 1607101874
transform 1 0 1908 0 -1 4705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_12
timestamp 1607101874
transform 1 0 1916 0 -1 4705
box -2 -3 74 103
use AOI21X1  AOI21X1_525
timestamp 1607101874
transform 1 0 1924 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_637
timestamp 1607101874
transform -1 0 1980 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1607101874
transform -1 0 2076 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_108
timestamp 1607101874
transform 1 0 1988 0 -1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_95
timestamp 1607101874
transform 1 0 2004 0 -1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_378
timestamp 1607101874
transform 1 0 2076 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1186
timestamp 1607101874
transform -1 0 2084 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_495
timestamp 1607101874
transform 1 0 2084 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_459
timestamp 1607101874
transform 1 0 2116 0 -1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_640
timestamp 1607101874
transform 1 0 2172 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_528
timestamp 1607101874
transform -1 0 2228 0 1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_353
timestamp 1607101874
transform -1 0 2180 0 -1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1607101874
transform 1 0 2180 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_409
timestamp 1607101874
transform 1 0 2228 0 1 4505
box -2 -3 98 103
use BUFX4  BUFX4_342
timestamp 1607101874
transform -1 0 2356 0 1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_584
timestamp 1607101874
transform 1 0 2276 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_696
timestamp 1607101874
transform 1 0 2308 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_44
timestamp 1607101874
transform 1 0 2356 0 1 4505
box -2 -3 34 103
use FILL  FILL_45_4_0
timestamp 1607101874
transform -1 0 2396 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_4_1
timestamp 1607101874
transform -1 0 2404 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_730
timestamp 1607101874
transform -1 0 2500 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_910
timestamp 1607101874
transform 1 0 2332 0 -1 4705
box -2 -3 98 103
use MUX2X1  MUX2X1_100
timestamp 1607101874
transform 1 0 2500 0 1 4505
box -2 -3 50 103
use FILL  FILL_46_4_0
timestamp 1607101874
transform 1 0 2428 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_4_1
timestamp 1607101874
transform 1 0 2436 0 -1 4705
box -2 -3 10 103
use NOR2X1  NOR2X1_178
timestamp 1607101874
transform 1 0 2444 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_113
timestamp 1607101874
transform 1 0 2468 0 -1 4705
box -2 -3 18 103
use AOI21X1  AOI21X1_582
timestamp 1607101874
transform 1 0 2484 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_694
timestamp 1607101874
transform -1 0 2540 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1607101874
transform 1 0 2548 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_698
timestamp 1607101874
transform -1 0 2564 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_586
timestamp 1607101874
transform -1 0 2596 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_266
timestamp 1607101874
transform 1 0 2596 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_924
timestamp 1607101874
transform -1 0 2740 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_362
timestamp 1607101874
transform 1 0 2692 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_369
timestamp 1607101874
transform 1 0 2740 0 1 4505
box -2 -3 26 103
use MUX2X1  MUX2X1_350
timestamp 1607101874
transform 1 0 2764 0 1 4505
box -2 -3 50 103
use AOI21X1  AOI21X1_254
timestamp 1607101874
transform 1 0 2812 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_229
timestamp 1607101874
transform 1 0 2788 0 -1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_301
timestamp 1607101874
transform -1 0 2852 0 -1 4705
box -2 -3 50 103
use OAI21X1  OAI21X1_1251
timestamp 1607101874
transform -1 0 2884 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_238
timestamp 1607101874
transform -1 0 2884 0 1 4505
box -2 -3 18 103
use NOR2X1  NOR2X1_365
timestamp 1607101874
transform -1 0 2868 0 1 4505
box -2 -3 26 103
use NOR2X1  NOR2X1_386
timestamp 1607101874
transform 1 0 2932 0 -1 4705
box -2 -3 26 103
use BUFX4  BUFX4_344
timestamp 1607101874
transform -1 0 2932 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_5_1
timestamp 1607101874
transform -1 0 2900 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_5_0
timestamp 1607101874
transform -1 0 2892 0 -1 4705
box -2 -3 10 103
use FILL  FILL_45_5_1
timestamp 1607101874
transform -1 0 2900 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_5_0
timestamp 1607101874
transform -1 0 2892 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1607101874
transform -1 0 2996 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_563
timestamp 1607101874
transform 1 0 2996 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_364
timestamp 1607101874
transform 1 0 3020 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_939
timestamp 1607101874
transform 1 0 2956 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_951
timestamp 1607101874
transform -1 0 3212 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_123
timestamp 1607101874
transform 1 0 3052 0 -1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_110
timestamp 1607101874
transform -1 0 3116 0 -1 4705
box -2 -3 50 103
use BUFX4  BUFX4_359
timestamp 1607101874
transform 1 0 3116 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1607101874
transform 1 0 3212 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_188
timestamp 1607101874
transform 1 0 3148 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_115
timestamp 1607101874
transform -1 0 3204 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_667
timestamp 1607101874
transform -1 0 3236 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1607101874
transform 1 0 3244 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_250
timestamp 1607101874
transform 1 0 3268 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_251
timestamp 1607101874
transform -1 0 3332 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_948
timestamp 1607101874
transform 1 0 3332 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_462
timestamp 1607101874
transform 1 0 3236 0 -1 4705
box -2 -3 26 103
use MUX2X1  MUX2X1_117
timestamp 1607101874
transform 1 0 3260 0 -1 4705
box -2 -3 50 103
use INVX1  INVX1_130
timestamp 1607101874
transform -1 0 3324 0 -1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_619
timestamp 1607101874
transform 1 0 3324 0 -1 4705
box -2 -3 26 103
use FILL  FILL_45_6_0
timestamp 1607101874
transform 1 0 3428 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_6_1
timestamp 1607101874
transform 1 0 3436 0 1 4505
box -2 -3 10 103
use NOR2X1  NOR2X1_620
timestamp 1607101874
transform 1 0 3348 0 -1 4705
box -2 -3 26 103
use OAI22X1  OAI22X1_90
timestamp 1607101874
transform -1 0 3412 0 -1 4705
box -2 -3 42 103
use FILL  FILL_46_6_0
timestamp 1607101874
transform 1 0 3412 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_6_1
timestamp 1607101874
transform 1 0 3420 0 -1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1249
timestamp 1607101874
transform 1 0 3428 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_461
timestamp 1607101874
transform 1 0 3444 0 1 4505
box -2 -3 26 103
use OAI22X1  OAI22X1_32
timestamp 1607101874
transform -1 0 3508 0 1 4505
box -2 -3 42 103
use OAI21X1  OAI21X1_898
timestamp 1607101874
transform -1 0 3540 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_897
timestamp 1607101874
transform 1 0 3460 0 -1 4705
box -2 -3 34 103
use MUX2X1  MUX2X1_116
timestamp 1607101874
transform 1 0 3492 0 -1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_449
timestamp 1607101874
transform 1 0 3540 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_381
timestamp 1607101874
transform 1 0 3636 0 1 4505
box -2 -3 18 103
use INVX1  INVX1_129
timestamp 1607101874
transform -1 0 3556 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1061
timestamp 1607101874
transform 1 0 3556 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_326
timestamp 1607101874
transform -1 0 3612 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_1252
timestamp 1607101874
transform 1 0 3612 0 -1 4705
box -2 -3 34 103
use MUX2X1  MUX2X1_363
timestamp 1607101874
transform -1 0 3700 0 1 4505
box -2 -3 50 103
use AOI21X1  AOI21X1_418
timestamp 1607101874
transform 1 0 3700 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_189
timestamp 1607101874
transform -1 0 3756 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_968
timestamp 1607101874
transform 1 0 3644 0 -1 4705
box -2 -3 98 103
use MUX2X1  MUX2X1_115
timestamp 1607101874
transform 1 0 3740 0 -1 4705
box -2 -3 50 103
use NOR2X1  NOR2X1_514
timestamp 1607101874
transform 1 0 3756 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_253
timestamp 1607101874
transform 1 0 3780 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_252
timestamp 1607101874
transform 1 0 3812 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_128
timestamp 1607101874
transform -1 0 3804 0 -1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_465
timestamp 1607101874
transform 1 0 3804 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_941
timestamp 1607101874
transform 1 0 3828 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_900
timestamp 1607101874
transform 1 0 3844 0 1 4505
box -2 -3 34 103
use OAI22X1  OAI22X1_47
timestamp 1607101874
transform 1 0 3876 0 1 4505
box -2 -3 42 103
use FILL  FILL_45_7_0
timestamp 1607101874
transform 1 0 3916 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_7_1
timestamp 1607101874
transform 1 0 3924 0 1 4505
box -2 -3 10 103
use NOR2X1  NOR2X1_513
timestamp 1607101874
transform 1 0 3932 0 1 4505
box -2 -3 26 103
use FILL  FILL_46_7_0
timestamp 1607101874
transform 1 0 3924 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_7_1
timestamp 1607101874
transform 1 0 3932 0 -1 4705
box -2 -3 10 103
use INVX1  INVX1_125
timestamp 1607101874
transform 1 0 3940 0 -1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_949
timestamp 1607101874
transform 1 0 3956 0 1 4505
box -2 -3 98 103
use MUX2X1  MUX2X1_112
timestamp 1607101874
transform -1 0 4004 0 -1 4705
box -2 -3 50 103
use AOI21X1  AOI21X1_593
timestamp 1607101874
transform 1 0 4004 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_705
timestamp 1607101874
transform -1 0 4060 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_960
timestamp 1607101874
transform 1 0 4052 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_512
timestamp 1607101874
transform -1 0 4108 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1444
timestamp 1607101874
transform 1 0 4108 0 1 4505
box -2 -3 34 103
use OAI22X1  OAI22X1_33
timestamp 1607101874
transform 1 0 4140 0 1 4505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_453
timestamp 1607101874
transform -1 0 4156 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_464
timestamp 1607101874
transform 1 0 4180 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1445
timestamp 1607101874
transform -1 0 4236 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_511
timestamp 1607101874
transform 1 0 4236 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_285
timestamp 1607101874
transform -1 0 4252 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_902
timestamp 1607101874
transform -1 0 4292 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_315
timestamp 1607101874
transform -1 0 4308 0 1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_448
timestamp 1607101874
transform -1 0 4404 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_957
timestamp 1607101874
transform 1 0 4252 0 -1 4705
box -2 -3 98 103
use BUFX4  BUFX4_341
timestamp 1607101874
transform -1 0 4436 0 1 4505
box -2 -3 34 103
use FILL  FILL_45_8_0
timestamp 1607101874
transform -1 0 4444 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_8_1
timestamp 1607101874
transform -1 0 4452 0 1 4505
box -2 -3 10 103
use NOR2X1  NOR2X1_207
timestamp 1607101874
transform -1 0 4372 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_129
timestamp 1607101874
transform -1 0 4404 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_8_0
timestamp 1607101874
transform -1 0 4412 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_8_1
timestamp 1607101874
transform -1 0 4420 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_976
timestamp 1607101874
transform -1 0 4516 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_217
timestamp 1607101874
transform -1 0 4476 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_137
timestamp 1607101874
transform -1 0 4508 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_986
timestamp 1607101874
transform -1 0 4604 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_209
timestamp 1607101874
transform -1 0 4540 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_978
timestamp 1607101874
transform 1 0 4540 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1244
timestamp 1607101874
transform 1 0 4604 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_714
timestamp 1607101874
transform -1 0 4668 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1101
timestamp 1607101874
transform 1 0 4636 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_408
timestamp 1607101874
transform 1 0 4668 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_712
timestamp 1607101874
transform -1 0 4724 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_899
timestamp 1607101874
transform -1 0 4756 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_97
timestamp 1607101874
transform -1 0 4692 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_52
timestamp 1607101874
transform -1 0 4724 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_767
timestamp 1607101874
transform -1 0 4820 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_652
timestamp 1607101874
transform 1 0 4756 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_540
timestamp 1607101874
transform -1 0 4812 0 1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_370
timestamp 1607101874
transform 1 0 4812 0 1 4505
box -2 -3 50 103
use BUFX4  BUFX4_370
timestamp 1607101874
transform -1 0 4852 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_580
timestamp 1607101874
transform 1 0 4860 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_469
timestamp 1607101874
transform 1 0 4884 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_100
timestamp 1607101874
transform 1 0 4852 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_55
timestamp 1607101874
transform -1 0 4908 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_9_0
timestamp 1607101874
transform -1 0 4916 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_9_1
timestamp 1607101874
transform -1 0 4924 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_770
timestamp 1607101874
transform -1 0 5020 0 -1 4705
box -2 -3 98 103
use FILL  FILL_45_9_0
timestamp 1607101874
transform -1 0 4988 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_9_1
timestamp 1607101874
transform -1 0 4996 0 1 4505
box -2 -3 10 103
use OAI21X1  OAI21X1_54
timestamp 1607101874
transform -1 0 5028 0 1 4505
box -2 -3 34 103
use BUFX4  BUFX4_355
timestamp 1607101874
transform -1 0 5060 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1238
timestamp 1607101874
transform -1 0 5052 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_196
timestamp 1607101874
transform 1 0 5052 0 -1 4705
box -2 -3 34 103
use BUFX4  BUFX4_368
timestamp 1607101874
transform 1 0 5060 0 1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_383
timestamp 1607101874
transform -1 0 5124 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_807
timestamp 1607101874
transform -1 0 5156 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_293
timestamp 1607101874
transform 1 0 5084 0 -1 4705
box -2 -3 26 103
use MUX2X1  MUX2X1_28
timestamp 1607101874
transform -1 0 5156 0 -1 4705
box -2 -3 50 103
use AOI21X1  AOI21X1_354
timestamp 1607101874
transform -1 0 5188 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_41
timestamp 1607101874
transform 1 0 5188 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_668
timestamp 1607101874
transform -1 0 5308 0 1 4505
box -2 -3 98 103
use MUX2X1  MUX2X1_167
timestamp 1607101874
transform 1 0 5156 0 -1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1607101874
transform -1 0 5300 0 -1 4705
box -2 -3 98 103
use FILL  FILL_47_1
timestamp 1607101874
transform -1 0 5308 0 -1 4705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_1
timestamp 1607101874
transform -1 0 60 0 1 4705
box -2 -3 58 103
use NAND2X1  NAND2X1_136
timestamp 1607101874
transform 1 0 60 0 1 4705
box -2 -3 26 103
use INVX1  INVX1_200
timestamp 1607101874
transform 1 0 84 0 1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_325
timestamp 1607101874
transform 1 0 100 0 1 4705
box -2 -3 26 103
use NAND3X1  NAND3X1_49
timestamp 1607101874
transform 1 0 124 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_497
timestamp 1607101874
transform 1 0 156 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_156
timestamp 1607101874
transform 1 0 188 0 1 4705
box -2 -3 26 103
use NAND2X1  NAND2X1_151
timestamp 1607101874
transform 1 0 212 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_400
timestamp 1607101874
transform 1 0 236 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_0_0
timestamp 1607101874
transform 1 0 332 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_0_1
timestamp 1607101874
transform 1 0 340 0 1 4705
box -2 -3 10 103
use NAND2X1  NAND2X1_152
timestamp 1607101874
transform 1 0 348 0 1 4705
box -2 -3 26 103
use NAND3X1  NAND3X1_48
timestamp 1607101874
transform -1 0 404 0 1 4705
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1607101874
transform -1 0 436 0 1 4705
box -2 -3 34 103
use INVX4  INVX4_11
timestamp 1607101874
transform 1 0 436 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_230
timestamp 1607101874
transform 1 0 460 0 1 4705
box -2 -3 34 103
use INVX2  INVX2_25
timestamp 1607101874
transform 1 0 492 0 1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_502
timestamp 1607101874
transform 1 0 508 0 1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_229
timestamp 1607101874
transform 1 0 540 0 1 4705
box -2 -3 34 103
use INVX2  INVX2_24
timestamp 1607101874
transform -1 0 588 0 1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_517
timestamp 1607101874
transform 1 0 588 0 1 4705
box -2 -3 34 103
use INVX1  INVX1_209
timestamp 1607101874
transform -1 0 636 0 1 4705
box -2 -3 18 103
use INVX2  INVX2_20
timestamp 1607101874
transform 1 0 636 0 1 4705
box -2 -3 18 103
use NAND3X1  NAND3X1_47
timestamp 1607101874
transform -1 0 684 0 1 4705
box -2 -3 34 103
use INVX1  INVX1_202
timestamp 1607101874
transform -1 0 700 0 1 4705
box -2 -3 18 103
use BUFX4  BUFX4_304
timestamp 1607101874
transform -1 0 732 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_144
timestamp 1607101874
transform -1 0 756 0 1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_516
timestamp 1607101874
transform -1 0 788 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_442
timestamp 1607101874
transform 1 0 788 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_475
timestamp 1607101874
transform 1 0 820 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_1_0
timestamp 1607101874
transform -1 0 860 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_1_1
timestamp 1607101874
transform -1 0 868 0 1 4705
box -2 -3 10 103
use AND2X2  AND2X2_2
timestamp 1607101874
transform -1 0 900 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_301
timestamp 1607101874
transform 1 0 900 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_222
timestamp 1607101874
transform -1 0 956 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_329
timestamp 1607101874
transform 1 0 956 0 1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_501
timestamp 1607101874
transform -1 0 1012 0 1 4705
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1607101874
transform -1 0 1044 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_494
timestamp 1607101874
transform -1 0 1076 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_300
timestamp 1607101874
transform -1 0 1100 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_213
timestamp 1607101874
transform 1 0 1100 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_462
timestamp 1607101874
transform 1 0 1132 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1607101874
transform -1 0 1196 0 1 4705
box -2 -3 34 103
use MUX2X1  MUX2X1_173
timestamp 1607101874
transform 1 0 1196 0 1 4705
box -2 -3 50 103
use OAI21X1  OAI21X1_441
timestamp 1607101874
transform -1 0 1276 0 1 4705
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1607101874
transform 1 0 1276 0 1 4705
box -2 -3 42 103
use NAND2X1  NAND2X1_103
timestamp 1607101874
transform -1 0 1340 0 1 4705
box -2 -3 26 103
use NAND2X1  NAND2X1_104
timestamp 1607101874
transform -1 0 1364 0 1 4705
box -2 -3 26 103
use FILL  FILL_47_2_0
timestamp 1607101874
transform -1 0 1372 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_2_1
timestamp 1607101874
transform -1 0 1380 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1607101874
transform -1 0 1476 0 1 4705
box -2 -3 98 103
use MUX2X1  MUX2X1_337
timestamp 1607101874
transform -1 0 1524 0 1 4705
box -2 -3 50 103
use MUX2X1  MUX2X1_339
timestamp 1607101874
transform -1 0 1572 0 1 4705
box -2 -3 50 103
use AOI21X1  AOI21X1_92
timestamp 1607101874
transform 1 0 1572 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_686
timestamp 1607101874
transform 1 0 1604 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_574
timestamp 1607101874
transform -1 0 1660 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_155
timestamp 1607101874
transform -1 0 1684 0 1 4705
box -2 -3 26 103
use MUX2X1  MUX2X1_42
timestamp 1607101874
transform 1 0 1684 0 1 4705
box -2 -3 50 103
use INVX1  INVX1_52
timestamp 1607101874
transform -1 0 1748 0 1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_722
timestamp 1607101874
transform -1 0 1844 0 1 4705
box -2 -3 98 103
use MUX2X1  MUX2X1_109
timestamp 1607101874
transform -1 0 1892 0 1 4705
box -2 -3 50 103
use FILL  FILL_47_3_0
timestamp 1607101874
transform 1 0 1892 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_3_1
timestamp 1607101874
transform 1 0 1900 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_875
timestamp 1607101874
transform 1 0 1908 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1607101874
transform -1 0 2100 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_852
timestamp 1607101874
transform -1 0 2132 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_576
timestamp 1607101874
transform 1 0 2132 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_183
timestamp 1607101874
transform -1 0 2188 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_113
timestamp 1607101874
transform -1 0 2220 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_531
timestamp 1607101874
transform -1 0 2244 0 1 4705
box -2 -3 26 103
use BUFX4  BUFX4_337
timestamp 1607101874
transform -1 0 2276 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_583
timestamp 1607101874
transform 1 0 2276 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_927
timestamp 1607101874
transform 1 0 2300 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_4_0
timestamp 1607101874
transform 1 0 2396 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_4_1
timestamp 1607101874
transform 1 0 2404 0 1 4705
box -2 -3 10 103
use AOI21X1  AOI21X1_109
timestamp 1607101874
transform 1 0 2412 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1607101874
transform 1 0 2444 0 1 4705
box -2 -3 98 103
use MUX2X1  MUX2X1_278
timestamp 1607101874
transform 1 0 2540 0 1 4705
box -2 -3 50 103
use INVX1  INVX1_447
timestamp 1607101874
transform -1 0 2604 0 1 4705
box -2 -3 18 103
use AOI21X1  AOI21X1_587
timestamp 1607101874
transform 1 0 2604 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_699
timestamp 1607101874
transform -1 0 2660 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_267
timestamp 1607101874
transform -1 0 2756 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_370
timestamp 1607101874
transform 1 0 2756 0 1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_538
timestamp 1607101874
transform -1 0 2884 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_650
timestamp 1607101874
transform 1 0 2884 0 1 4705
box -2 -3 26 103
use FILL  FILL_47_5_0
timestamp 1607101874
transform -1 0 2916 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_5_1
timestamp 1607101874
transform -1 0 2924 0 1 4705
box -2 -3 10 103
use NOR2X1  NOR2X1_387
timestamp 1607101874
transform -1 0 2948 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_478
timestamp 1607101874
transform 1 0 2948 0 1 4705
box -2 -3 98 103
use INVX1  INVX1_434
timestamp 1607101874
transform 1 0 3044 0 1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_377
timestamp 1607101874
transform -1 0 3108 0 1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_952
timestamp 1607101874
transform -1 0 3204 0 1 4705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_9
timestamp 1607101874
transform -1 0 3276 0 1 4705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_970
timestamp 1607101874
transform 1 0 3276 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_6_0
timestamp 1607101874
transform 1 0 3372 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_6_1
timestamp 1607101874
transform 1 0 3380 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_944
timestamp 1607101874
transform 1 0 3388 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_969
timestamp 1607101874
transform 1 0 3484 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_965
timestamp 1607101874
transform -1 0 3676 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1463
timestamp 1607101874
transform 1 0 3676 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1464
timestamp 1607101874
transform -1 0 3740 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_458
timestamp 1607101874
transform 1 0 3740 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1062
timestamp 1607101874
transform 1 0 3836 0 1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_483
timestamp 1607101874
transform 1 0 3868 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1153
timestamp 1607101874
transform -1 0 3932 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_7_0
timestamp 1607101874
transform 1 0 3932 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_7_1
timestamp 1607101874
transform 1 0 3940 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_957
timestamp 1607101874
transform 1 0 3948 0 1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_416
timestamp 1607101874
transform -1 0 4012 0 1 4705
box -2 -3 34 103
use BUFX4  BUFX4_348
timestamp 1607101874
transform -1 0 4044 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_194
timestamp 1607101874
transform -1 0 4068 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_120
timestamp 1607101874
transform -1 0 4100 0 1 4705
box -2 -3 34 103
use MUX2X1  MUX2X1_369
timestamp 1607101874
transform -1 0 4148 0 1 4705
box -2 -3 50 103
use MUX2X1  MUX2X1_359
timestamp 1607101874
transform 1 0 4148 0 1 4705
box -2 -3 50 103
use INVX1  INVX1_379
timestamp 1607101874
transform -1 0 4212 0 1 4705
box -2 -3 18 103
use NOR2X1  NOR2X1_373
timestamp 1607101874
transform -1 0 4236 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_276
timestamp 1607101874
transform -1 0 4332 0 1 4705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_102
timestamp 1607101874
transform -1 0 4404 0 1 4705
box -2 -3 74 103
use BUFX4  BUFX4_362
timestamp 1607101874
transform -1 0 4436 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_8_0
timestamp 1607101874
transform 1 0 4436 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_8_1
timestamp 1607101874
transform 1 0 4444 0 1 4705
box -2 -3 10 103
use AOI21X1  AOI21X1_131
timestamp 1607101874
transform 1 0 4452 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_713
timestamp 1607101874
transform 1 0 4484 0 1 4705
box -2 -3 34 103
use INVX1  INVX1_73
timestamp 1607101874
transform 1 0 4516 0 1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_63
timestamp 1607101874
transform -1 0 4580 0 1 4705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_775
timestamp 1607101874
transform -1 0 4676 0 1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_469
timestamp 1607101874
transform 1 0 4676 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_198
timestamp 1607101874
transform -1 0 4732 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_123
timestamp 1607101874
transform -1 0 4764 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_960
timestamp 1607101874
transform -1 0 4860 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1607101874
transform 1 0 4860 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_9_0
timestamp 1607101874
transform -1 0 4964 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_9_1
timestamp 1607101874
transform -1 0 4972 0 1 4705
box -2 -3 10 103
use AOI21X1  AOI21X1_508
timestamp 1607101874
transform -1 0 5004 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1149
timestamp 1607101874
transform -1 0 5036 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_665
timestamp 1607101874
transform -1 0 5132 0 1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_18
timestamp 1607101874
transform 1 0 5132 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1607101874
transform -1 0 5188 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_670
timestamp 1607101874
transform -1 0 5284 0 1 4705
box -2 -3 98 103
use FILL  FILL_48_1
timestamp 1607101874
transform 1 0 5284 0 1 4705
box -2 -3 10 103
use FILL  FILL_48_2
timestamp 1607101874
transform 1 0 5292 0 1 4705
box -2 -3 10 103
use FILL  FILL_48_3
timestamp 1607101874
transform 1 0 5300 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_405
timestamp 1607101874
transform -1 0 100 0 -1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_324
timestamp 1607101874
transform -1 0 124 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_526
timestamp 1607101874
transform 1 0 124 0 -1 4905
box -2 -3 34 103
use INVX1  INVX1_210
timestamp 1607101874
transform -1 0 172 0 -1 4905
box -2 -3 18 103
use AOI22X1  AOI22X1_8
timestamp 1607101874
transform -1 0 212 0 -1 4905
box -2 -3 42 103
use OAI21X1  OAI21X1_529
timestamp 1607101874
transform -1 0 244 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_523
timestamp 1607101874
transform 1 0 244 0 -1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_59
timestamp 1607101874
transform -1 0 308 0 -1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_51
timestamp 1607101874
transform 1 0 308 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_0_0
timestamp 1607101874
transform -1 0 348 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_0_1
timestamp 1607101874
transform -1 0 356 0 -1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_511
timestamp 1607101874
transform -1 0 388 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_512
timestamp 1607101874
transform 1 0 388 0 -1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_53
timestamp 1607101874
transform 1 0 420 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_518
timestamp 1607101874
transform 1 0 452 0 -1 4905
box -2 -3 34 103
use AOI22X1  AOI22X1_5
timestamp 1607101874
transform 1 0 484 0 -1 4905
box -2 -3 42 103
use NAND2X1  NAND2X1_141
timestamp 1607101874
transform -1 0 548 0 -1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_232
timestamp 1607101874
transform 1 0 548 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_507
timestamp 1607101874
transform 1 0 580 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_234
timestamp 1607101874
transform 1 0 612 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_508
timestamp 1607101874
transform -1 0 676 0 -1 4905
box -2 -3 34 103
use NOR3X1  NOR3X1_11
timestamp 1607101874
transform 1 0 676 0 -1 4905
box -2 -3 66 103
use AOI21X1  AOI21X1_235
timestamp 1607101874
transform 1 0 740 0 -1 4905
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1607101874
transform -1 0 812 0 -1 4905
box -2 -3 42 103
use OAI21X1  OAI21X1_495
timestamp 1607101874
transform -1 0 844 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_1_0
timestamp 1607101874
transform 1 0 844 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_1_1
timestamp 1607101874
transform 1 0 852 0 -1 4905
box -2 -3 10 103
use NOR2X1  NOR2X1_333
timestamp 1607101874
transform 1 0 860 0 -1 4905
box -2 -3 26 103
use NOR2X1  NOR2X1_332
timestamp 1607101874
transform -1 0 908 0 -1 4905
box -2 -3 26 103
use INVX1  INVX1_204
timestamp 1607101874
transform -1 0 924 0 -1 4905
box -2 -3 18 103
use BUFX4  BUFX4_306
timestamp 1607101874
transform 1 0 924 0 -1 4905
box -2 -3 34 103
use INVX1  INVX1_205
timestamp 1607101874
transform -1 0 972 0 -1 4905
box -2 -3 18 103
use OAI21X1  OAI21X1_496
timestamp 1607101874
transform 1 0 972 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1607101874
transform 1 0 1004 0 -1 4905
box -2 -3 26 103
use NOR2X1  NOR2X1_330
timestamp 1607101874
transform -1 0 1052 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_498
timestamp 1607101874
transform -1 0 1084 0 -1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1607101874
transform 1 0 1084 0 -1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1607101874
transform 1 0 1116 0 -1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1607101874
transform -1 0 1172 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_443
timestamp 1607101874
transform 1 0 1172 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_461
timestamp 1607101874
transform -1 0 1236 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_212
timestamp 1607101874
transform -1 0 1268 0 -1 4905
box -2 -3 34 103
use INVX2  INVX2_17
timestamp 1607101874
transform -1 0 1284 0 -1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_422
timestamp 1607101874
transform -1 0 1380 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_2_0
timestamp 1607101874
transform 1 0 1380 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_2_1
timestamp 1607101874
transform 1 0 1388 0 -1 4905
box -2 -3 10 103
use AND2X2  AND2X2_18
timestamp 1607101874
transform 1 0 1396 0 -1 4905
box -2 -3 34 103
use AND2X2  AND2X2_17
timestamp 1607101874
transform -1 0 1460 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_358
timestamp 1607101874
transform -1 0 1484 0 -1 4905
box -2 -3 26 103
use INVX4  INVX4_9
timestamp 1607101874
transform 1 0 1484 0 -1 4905
box -2 -3 26 103
use INVX1  INVX1_241
timestamp 1607101874
transform -1 0 1524 0 -1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1607101874
transform -1 0 1620 0 -1 4905
box -2 -3 98 103
use INVX8  INVX8_15
timestamp 1607101874
transform -1 0 1660 0 -1 4905
box -2 -3 42 103
use CLKBUF1  CLKBUF1_101
timestamp 1607101874
transform -1 0 1732 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_936
timestamp 1607101874
transform 1 0 1732 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_122
timestamp 1607101874
transform 1 0 1828 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_96
timestamp 1607101874
transform 1 0 1844 0 -1 4905
box -2 -3 50 103
use FILL  FILL_48_3_0
timestamp 1607101874
transform 1 0 1892 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_3_1
timestamp 1607101874
transform 1 0 1900 0 -1 4905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_86
timestamp 1607101874
transform 1 0 1908 0 -1 4905
box -2 -3 74 103
use AOI21X1  AOI21X1_110
timestamp 1607101874
transform 1 0 1980 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_179
timestamp 1607101874
transform -1 0 2036 0 -1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1607101874
transform 1 0 2036 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_239
timestamp 1607101874
transform 1 0 2132 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_354
timestamp 1607101874
transform 1 0 2148 0 -1 4905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_938
timestamp 1607101874
transform 1 0 2196 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_930
timestamp 1607101874
transform 1 0 2292 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_4_0
timestamp 1607101874
transform 1 0 2388 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_4_1
timestamp 1607101874
transform 1 0 2396 0 -1 4905
box -2 -3 10 103
use INVX1  INVX1_121
timestamp 1607101874
transform 1 0 2404 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_108
timestamp 1607101874
transform -1 0 2468 0 -1 4905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_366
timestamp 1607101874
transform 1 0 2468 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_449
timestamp 1607101874
transform 1 0 2564 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_297
timestamp 1607101874
transform -1 0 2628 0 -1 4905
box -2 -3 50 103
use NOR2X1  NOR2X1_366
timestamp 1607101874
transform -1 0 2652 0 -1 4905
box -2 -3 26 103
use NOR2X1  NOR2X1_174
timestamp 1607101874
transform -1 0 2676 0 -1 4905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_61
timestamp 1607101874
transform 1 0 2676 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_274
timestamp 1607101874
transform 1 0 2748 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_257
timestamp 1607101874
transform 1 0 2844 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_357
timestamp 1607101874
transform -1 0 2908 0 -1 4905
box -2 -3 50 103
use FILL  FILL_48_5_0
timestamp 1607101874
transform 1 0 2908 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_5_1
timestamp 1607101874
transform 1 0 2916 0 -1 4905
box -2 -3 10 103
use BUFX4  BUFX4_369
timestamp 1607101874
transform 1 0 2924 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_275
timestamp 1607101874
transform 1 0 2956 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_599
timestamp 1607101874
transform 1 0 2988 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_666
timestamp 1607101874
transform 1 0 3020 0 -1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_210
timestamp 1607101874
transform -1 0 3076 0 -1 4905
box -2 -3 26 103
use MUX2X1  MUX2X1_111
timestamp 1607101874
transform 1 0 3076 0 -1 4905
box -2 -3 50 103
use INVX1  INVX1_124
timestamp 1607101874
transform -1 0 3140 0 -1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_940
timestamp 1607101874
transform 1 0 3140 0 -1 4905
box -2 -3 98 103
use BUFX4  BUFX4_466
timestamp 1607101874
transform -1 0 3268 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_121
timestamp 1607101874
transform 1 0 3268 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_195
timestamp 1607101874
transform -1 0 3324 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_242
timestamp 1607101874
transform 1 0 3324 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_243
timestamp 1607101874
transform -1 0 3388 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_6_0
timestamp 1607101874
transform 1 0 3388 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_6_1
timestamp 1607101874
transform 1 0 3396 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_966
timestamp 1607101874
transform 1 0 3404 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_260
timestamp 1607101874
transform 1 0 3500 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_261
timestamp 1607101874
transform -1 0 3564 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_263
timestamp 1607101874
transform 1 0 3564 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_262
timestamp 1607101874
transform -1 0 3628 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_259
timestamp 1607101874
transform 1 0 3628 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_258
timestamp 1607101874
transform 1 0 3660 0 -1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_238
timestamp 1607101874
transform 1 0 3692 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_773
timestamp 1607101874
transform -1 0 3748 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1607101874
transform 1 0 3748 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_245
timestamp 1607101874
transform -1 0 3812 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_284
timestamp 1607101874
transform 1 0 3812 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_7_0
timestamp 1607101874
transform 1 0 3908 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_7_1
timestamp 1607101874
transform 1 0 3916 0 -1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_1442
timestamp 1607101874
transform 1 0 3924 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_1443
timestamp 1607101874
transform -1 0 3988 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1607101874
transform 1 0 3988 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_193
timestamp 1607101874
transform -1 0 4044 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_1060
timestamp 1607101874
transform 1 0 4044 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_124
timestamp 1607101874
transform 1 0 4076 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_199
timestamp 1607101874
transform 1 0 4108 0 -1 4905
box -2 -3 26 103
use INVX1  INVX1_254
timestamp 1607101874
transform -1 0 4148 0 -1 4905
box -2 -3 18 103
use BUFX4  BUFX4_475
timestamp 1607101874
transform 1 0 4148 0 -1 4905
box -2 -3 34 103
use MUX2X1  MUX2X1_375
timestamp 1607101874
transform -1 0 4228 0 -1 4905
box -2 -3 50 103
use INVX1  INVX1_255
timestamp 1607101874
transform -1 0 4244 0 -1 4905
box -2 -3 18 103
use NOR2X1  NOR2X1_467
timestamp 1607101874
transform -1 0 4268 0 -1 4905
box -2 -3 26 103
use NOR2X1  NOR2X1_215
timestamp 1607101874
transform -1 0 4292 0 -1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_135
timestamp 1607101874
transform -1 0 4324 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_984
timestamp 1607101874
transform -1 0 4420 0 -1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_481
timestamp 1607101874
transform -1 0 4444 0 -1 4905
box -2 -3 26 103
use FILL  FILL_48_8_0
timestamp 1607101874
transform 1 0 4444 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_8_1
timestamp 1607101874
transform 1 0 4452 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_365
timestamp 1607101874
transform 1 0 4460 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_451
timestamp 1607101874
transform 1 0 4556 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_304
timestamp 1607101874
transform -1 0 4620 0 -1 4905
box -2 -3 50 103
use MUX2X1  MUX2X1_66
timestamp 1607101874
transform 1 0 4620 0 -1 4905
box -2 -3 50 103
use INVX1  INVX1_76
timestamp 1607101874
transform -1 0 4684 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_169
timestamp 1607101874
transform 1 0 4684 0 -1 4905
box -2 -3 50 103
use INVX1  INVX1_183
timestamp 1607101874
transform -1 0 4748 0 -1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1607101874
transform -1 0 4844 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_666
timestamp 1607101874
transform 1 0 4844 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_9_0
timestamp 1607101874
transform 1 0 4940 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_9_1
timestamp 1607101874
transform 1 0 4948 0 -1 4905
box -2 -3 10 103
use INVX1  INVX1_37
timestamp 1607101874
transform 1 0 4956 0 -1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_29
timestamp 1607101874
transform -1 0 5020 0 -1 4905
box -2 -3 50 103
use AOI21X1  AOI21X1_482
timestamp 1607101874
transform 1 0 5020 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_314
timestamp 1607101874
transform -1 0 5084 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_660
timestamp 1607101874
transform -1 0 5180 0 -1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_103
timestamp 1607101874
transform 1 0 5180 0 -1 4905
box -2 -3 74 103
use OAI21X1  OAI21X1_910
timestamp 1607101874
transform 1 0 5252 0 -1 4905
box -2 -3 34 103
use BUFX2  BUFX2_8
timestamp 1607101874
transform 1 0 5284 0 -1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_394
timestamp 1607101874
transform -1 0 100 0 1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_530
timestamp 1607101874
transform -1 0 132 0 1 4905
box -2 -3 34 103
use INVX1  INVX1_211
timestamp 1607101874
transform 1 0 132 0 1 4905
box -2 -3 18 103
use NAND3X1  NAND3X1_65
timestamp 1607101874
transform 1 0 148 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_240
timestamp 1607101874
transform 1 0 180 0 1 4905
box -2 -3 34 103
use AOI22X1  AOI22X1_6
timestamp 1607101874
transform -1 0 252 0 1 4905
box -2 -3 42 103
use INVX1  INVX1_203
timestamp 1607101874
transform 1 0 252 0 1 4905
box -2 -3 18 103
use NAND3X1  NAND3X1_45
timestamp 1607101874
transform 1 0 268 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_505
timestamp 1607101874
transform 1 0 300 0 1 4905
box -2 -3 34 103
use FILL  FILL_49_0_0
timestamp 1607101874
transform -1 0 340 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_0_1
timestamp 1607101874
transform -1 0 348 0 1 4905
box -2 -3 10 103
use AOI21X1  AOI21X1_238
timestamp 1607101874
transform -1 0 380 0 1 4905
box -2 -3 34 103
use INVX1  INVX1_207
timestamp 1607101874
transform 1 0 380 0 1 4905
box -2 -3 18 103
use AOI21X1  AOI21X1_237
timestamp 1607101874
transform -1 0 428 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_515
timestamp 1607101874
transform -1 0 460 0 1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1607101874
transform 1 0 460 0 1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_334
timestamp 1607101874
transform -1 0 516 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_506
timestamp 1607101874
transform -1 0 548 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_239
timestamp 1607101874
transform -1 0 580 0 1 4905
box -2 -3 34 103
use AND2X2  AND2X2_12
timestamp 1607101874
transform -1 0 612 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_509
timestamp 1607101874
transform 1 0 612 0 1 4905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_4
timestamp 1607101874
transform -1 0 700 0 1 4905
box -2 -3 58 103
use NAND2X1  NAND2X1_143
timestamp 1607101874
transform -1 0 724 0 1 4905
box -2 -3 26 103
use NAND3X1  NAND3X1_46
timestamp 1607101874
transform 1 0 724 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_236
timestamp 1607101874
transform -1 0 788 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_525
timestamp 1607101874
transform -1 0 820 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_522
timestamp 1607101874
transform 1 0 820 0 1 4905
box -2 -3 34 103
use FILL  FILL_49_1_0
timestamp 1607101874
transform 1 0 852 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_1_1
timestamp 1607101874
transform 1 0 860 0 1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_521
timestamp 1607101874
transform 1 0 868 0 1 4905
box -2 -3 34 103
use OR2X2  OR2X2_6
timestamp 1607101874
transform -1 0 932 0 1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1607101874
transform 1 0 932 0 1 4905
box -2 -3 26 103
use AND2X2  AND2X2_10
timestamp 1607101874
transform -1 0 988 0 1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_142
timestamp 1607101874
transform -1 0 1012 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_499
timestamp 1607101874
transform -1 0 1044 0 1 4905
box -2 -3 34 103
use NAND2X1  NAND2X1_164
timestamp 1607101874
transform -1 0 1068 0 1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_423
timestamp 1607101874
transform -1 0 1164 0 1 4905
box -2 -3 98 103
use MUX2X1  MUX2X1_176
timestamp 1607101874
transform -1 0 1212 0 1 4905
box -2 -3 50 103
use NAND3X1  NAND3X1_68
timestamp 1607101874
transform -1 0 1244 0 1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_348
timestamp 1607101874
transform 1 0 1244 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_538
timestamp 1607101874
transform 1 0 1268 0 1 4905
box -2 -3 34 103
use AND2X2  AND2X2_15
timestamp 1607101874
transform 1 0 1300 0 1 4905
box -2 -3 34 103
use NAND3X1  NAND3X1_67
timestamp 1607101874
transform 1 0 1332 0 1 4905
box -2 -3 34 103
use FILL  FILL_49_2_0
timestamp 1607101874
transform 1 0 1364 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_2_1
timestamp 1607101874
transform 1 0 1372 0 1 4905
box -2 -3 10 103
use NOR2X1  NOR2X1_359
timestamp 1607101874
transform 1 0 1380 0 1 4905
box -2 -3 26 103
use AND2X2  AND2X2_19
timestamp 1607101874
transform 1 0 1404 0 1 4905
box -2 -3 34 103
use BUFX2  BUFX2_10
timestamp 1607101874
transform -1 0 1460 0 1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_393
timestamp 1607101874
transform 1 0 1460 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_391
timestamp 1607101874
transform -1 0 1652 0 1 4905
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1607101874
transform -1 0 1676 0 1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_390
timestamp 1607101874
transform -1 0 1772 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_876
timestamp 1607101874
transform 1 0 1772 0 1 4905
box -2 -3 98 103
use FILL  FILL_49_3_0
timestamp 1607101874
transform -1 0 1876 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_3_1
timestamp 1607101874
transform -1 0 1884 0 1 4905
box -2 -3 10 103
use INVX1  INVX1_109
timestamp 1607101874
transform -1 0 1900 0 1 4905
box -2 -3 18 103
use NAND2X1  NAND2X1_34
timestamp 1607101874
transform 1 0 1900 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_92
timestamp 1607101874
transform -1 0 1956 0 1 4905
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1607101874
transform 1 0 1956 0 1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_928
timestamp 1607101874
transform 1 0 1972 0 1 4905
box -2 -3 98 103
use INVX1  INVX1_235
timestamp 1607101874
transform 1 0 2068 0 1 4905
box -2 -3 18 103
use AOI21X1  AOI21X1_374
timestamp 1607101874
transform 1 0 2084 0 1 4905
box -2 -3 34 103
use MUX2X1  MUX2X1_346
timestamp 1607101874
transform -1 0 2164 0 1 4905
box -2 -3 50 103
use MUX2X1  MUX2X1_348
timestamp 1607101874
transform -1 0 2212 0 1 4905
box -2 -3 50 103
use INVX1  INVX1_419
timestamp 1607101874
transform -1 0 2228 0 1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1607101874
transform 1 0 2228 0 1 4905
box -2 -3 98 103
use AOI21X1  AOI21X1_104
timestamp 1607101874
transform 1 0 2324 0 1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_171
timestamp 1607101874
transform -1 0 2380 0 1 4905
box -2 -3 26 103
use FILL  FILL_49_4_0
timestamp 1607101874
transform 1 0 2380 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_4_1
timestamp 1607101874
transform 1 0 2388 0 1 4905
box -2 -3 10 103
use AOI21X1  AOI21X1_373
timestamp 1607101874
transform 1 0 2396 0 1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_172
timestamp 1607101874
transform 1 0 2428 0 1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_105
timestamp 1607101874
transform -1 0 2484 0 1 4905
box -2 -3 34 103
use INVX1  INVX1_115
timestamp 1607101874
transform 1 0 2484 0 1 4905
box -2 -3 18 103
use MUX2X1  MUX2X1_102
timestamp 1607101874
transform -1 0 2548 0 1 4905
box -2 -3 50 103
use OAI21X1  OAI21X1_849
timestamp 1607101874
transform 1 0 2548 0 1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_368
timestamp 1607101874
transform -1 0 2604 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_665
timestamp 1607101874
transform 1 0 2604 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_106
timestamp 1607101874
transform 1 0 2636 0 1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_919
timestamp 1607101874
transform 1 0 2668 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_955
timestamp 1607101874
transform 1 0 2764 0 1 4905
box -2 -3 98 103
use AOI21X1  AOI21X1_118
timestamp 1607101874
transform 1 0 2860 0 1 4905
box -2 -3 34 103
use FILL  FILL_49_5_0
timestamp 1607101874
transform 1 0 2892 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_5_1
timestamp 1607101874
transform 1 0 2900 0 1 4905
box -2 -3 10 103
use NOR2X1  NOR2X1_192
timestamp 1607101874
transform 1 0 2908 0 1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_602
timestamp 1607101874
transform -1 0 2964 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_277
timestamp 1607101874
transform -1 0 2996 0 1 4905
box -2 -3 34 103
use INVX1  INVX1_259
timestamp 1607101874
transform -1 0 3012 0 1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_447
timestamp 1607101874
transform -1 0 3108 0 1 4905
box -2 -3 98 103
use MUX2X1  MUX2X1_361
timestamp 1607101874
transform 1 0 3108 0 1 4905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_943
timestamp 1607101874
transform 1 0 3156 0 1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_241
timestamp 1607101874
transform 1 0 3252 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_240
timestamp 1607101874
transform -1 0 3316 0 1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_958
timestamp 1607101874
transform -1 0 3412 0 1 4905
box -2 -3 98 103
use FILL  FILL_49_6_0
timestamp 1607101874
transform -1 0 3420 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_6_1
timestamp 1607101874
transform -1 0 3428 0 1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_963
timestamp 1607101874
transform -1 0 3524 0 1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_256
timestamp 1607101874
transform -1 0 3556 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_257
timestamp 1607101874
transform -1 0 3588 0 1 4905
box -2 -3 34 103
use BUFX4  BUFX4_435
timestamp 1607101874
transform 1 0 3588 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_1460
timestamp 1607101874
transform 1 0 3620 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_1459
timestamp 1607101874
transform 1 0 3652 0 1 4905
box -2 -3 34 103
use MUX2X1  MUX2X1_360
timestamp 1607101874
transform -1 0 3732 0 1 4905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_964
timestamp 1607101874
transform 1 0 3732 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_945
timestamp 1607101874
transform -1 0 3924 0 1 4905
box -2 -3 98 103
use FILL  FILL_49_7_0
timestamp 1607101874
transform 1 0 3924 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_7_1
timestamp 1607101874
transform 1 0 3932 0 1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_956
timestamp 1607101874
transform 1 0 3940 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_961
timestamp 1607101874
transform -1 0 4132 0 1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_1440
timestamp 1607101874
transform 1 0 4132 0 1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_1441
timestamp 1607101874
transform -1 0 4196 0 1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_283
timestamp 1607101874
transform -1 0 4292 0 1 4905
box -2 -3 98 103
use AOI21X1  AOI21X1_485
timestamp 1607101874
transform 1 0 4292 0 1 4905
box -2 -3 34 103
use MUX2X1  MUX2X1_376
timestamp 1607101874
transform -1 0 4372 0 1 4905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_475
timestamp 1607101874
transform -1 0 4468 0 1 4905
box -2 -3 98 103
use FILL  FILL_49_8_0
timestamp 1607101874
transform 1 0 4468 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_8_1
timestamp 1607101874
transform 1 0 4476 0 1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_1156
timestamp 1607101874
transform 1 0 4484 0 1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_312
timestamp 1607101874
transform 1 0 4516 0 1 4905
box -2 -3 34 103
use MUX2X1  MUX2X1_59
timestamp 1607101874
transform -1 0 4596 0 1 4905
box -2 -3 50 103
use MUX2X1  MUX2X1_300
timestamp 1607101874
transform 1 0 4596 0 1 4905
box -2 -3 50 103
use INVX1  INVX1_416
timestamp 1607101874
transform -1 0 4660 0 1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_369
timestamp 1607101874
transform -1 0 4756 0 1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_706
timestamp 1607101874
transform 1 0 4756 0 1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_594
timestamp 1607101874
transform -1 0 4812 0 1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_778
timestamp 1607101874
transform 1 0 4812 0 1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_95
timestamp 1607101874
transform -1 0 4980 0 1 4905
box -2 -3 74 103
use FILL  FILL_49_9_0
timestamp 1607101874
transform -1 0 4988 0 1 4905
box -2 -3 10 103
use FILL  FILL_49_9_1
timestamp 1607101874
transform -1 0 4996 0 1 4905
box -2 -3 10 103
use INVX1  INVX1_331
timestamp 1607101874
transform -1 0 5012 0 1 4905
box -2 -3 18 103
use OAI21X1  OAI21X1_45
timestamp 1607101874
transform 1 0 5012 0 1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1607101874
transform -1 0 5140 0 1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_340
timestamp 1607101874
transform 1 0 5140 0 1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_88
timestamp 1607101874
transform -1 0 5308 0 1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_426
timestamp 1607101874
transform 1 0 4 0 -1 5105
box -2 -3 98 103
use NAND2X1  NAND2X1_158
timestamp 1607101874
transform 1 0 100 0 -1 5105
box -2 -3 26 103
use AND2X2  AND2X2_14
timestamp 1607101874
transform -1 0 156 0 -1 5105
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1607101874
transform -1 0 180 0 -1 5105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_427
timestamp 1607101874
transform 1 0 180 0 -1 5105
box -2 -3 98 103
use NAND2X1  NAND2X1_147
timestamp 1607101874
transform 1 0 276 0 -1 5105
box -2 -3 26 103
use NAND2X1  NAND2X1_148
timestamp 1607101874
transform -1 0 324 0 -1 5105
box -2 -3 26 103
use INVX1  INVX1_208
timestamp 1607101874
transform 1 0 324 0 -1 5105
box -2 -3 18 103
use FILL  FILL_50_0_0
timestamp 1607101874
transform -1 0 348 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_0_1
timestamp 1607101874
transform -1 0 356 0 -1 5105
box -2 -3 10 103
use OAI21X1  OAI21X1_510
timestamp 1607101874
transform -1 0 388 0 -1 5105
box -2 -3 34 103
use AOI21X1  AOI21X1_233
timestamp 1607101874
transform -1 0 420 0 -1 5105
box -2 -3 34 103
use AND2X2  AND2X2_11
timestamp 1607101874
transform -1 0 452 0 -1 5105
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1607101874
transform 1 0 452 0 -1 5105
box -2 -3 34 103
use OAI21X1  OAI21X1_514
timestamp 1607101874
transform -1 0 516 0 -1 5105
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1607101874
transform -1 0 540 0 -1 5105
box -2 -3 26 103
use AOI21X1  AOI21X1_231
timestamp 1607101874
transform -1 0 572 0 -1 5105
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1607101874
transform -1 0 604 0 -1 5105
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1607101874
transform -1 0 628 0 -1 5105
box -2 -3 26 103
use NOR3X1  NOR3X1_12
timestamp 1607101874
transform 1 0 628 0 -1 5105
box -2 -3 66 103
use AOI21X1  AOI21X1_228
timestamp 1607101874
transform -1 0 724 0 -1 5105
box -2 -3 34 103
use NAND2X1  NAND2X1_149
timestamp 1607101874
transform 1 0 724 0 -1 5105
box -2 -3 26 103
use OAI21X1  OAI21X1_504
timestamp 1607101874
transform 1 0 748 0 -1 5105
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1607101874
transform -1 0 804 0 -1 5105
box -2 -3 26 103
use INVX1  INVX1_206
timestamp 1607101874
transform -1 0 820 0 -1 5105
box -2 -3 18 103
use NAND2X1  NAND2X1_146
timestamp 1607101874
transform -1 0 844 0 -1 5105
box -2 -3 26 103
use FILL  FILL_50_1_0
timestamp 1607101874
transform -1 0 852 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_1_1
timestamp 1607101874
transform -1 0 860 0 -1 5105
box -2 -3 10 103
use OAI21X1  OAI21X1_500
timestamp 1607101874
transform -1 0 892 0 -1 5105
box -2 -3 34 103
use OAI21X1  OAI21X1_503
timestamp 1607101874
transform 1 0 892 0 -1 5105
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1607101874
transform 1 0 924 0 -1 5105
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1607101874
transform -1 0 972 0 -1 5105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_395
timestamp 1607101874
transform -1 0 1068 0 -1 5105
box -2 -3 98 103
use NOR2X1  NOR2X1_349
timestamp 1607101874
transform -1 0 1092 0 -1 5105
box -2 -3 26 103
use NAND2X1  NAND2X1_162
timestamp 1607101874
transform -1 0 1116 0 -1 5105
box -2 -3 26 103
use INVX2  INVX2_16
timestamp 1607101874
transform 1 0 1116 0 -1 5105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_421
timestamp 1607101874
transform -1 0 1228 0 -1 5105
box -2 -3 98 103
use NOR2X1  NOR2X1_343
timestamp 1607101874
transform 1 0 1228 0 -1 5105
box -2 -3 26 103
use NAND2X1  NAND2X1_163
timestamp 1607101874
transform 1 0 1252 0 -1 5105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_7
timestamp 1607101874
transform -1 0 1332 0 -1 5105
box -2 -3 58 103
use FILL  FILL_50_2_0
timestamp 1607101874
transform 1 0 1332 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_2_1
timestamp 1607101874
transform 1 0 1340 0 -1 5105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_392
timestamp 1607101874
transform 1 0 1348 0 -1 5105
box -2 -3 98 103
use BUFX2  BUFX2_9
timestamp 1607101874
transform 1 0 1444 0 -1 5105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_59
timestamp 1607101874
transform -1 0 1540 0 -1 5105
box -2 -3 74 103
use BUFX2  BUFX2_2
timestamp 1607101874
transform -1 0 1564 0 -1 5105
box -2 -3 26 103
use BUFX4  BUFX4_8
timestamp 1607101874
transform 1 0 1564 0 -1 5105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_27
timestamp 1607101874
transform 1 0 1596 0 -1 5105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_41
timestamp 1607101874
transform 1 0 1668 0 -1 5105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_37
timestamp 1607101874
transform 1 0 1740 0 -1 5105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_718
timestamp 1607101874
transform 1 0 1812 0 -1 5105
box -2 -3 98 103
use FILL  FILL_50_3_0
timestamp 1607101874
transform 1 0 1908 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_3_1
timestamp 1607101874
transform 1 0 1916 0 -1 5105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1607101874
transform 1 0 1924 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_920
timestamp 1607101874
transform -1 0 2116 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_912
timestamp 1607101874
transform 1 0 2116 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_959
timestamp 1607101874
transform 1 0 2212 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_914
timestamp 1607101874
transform 1 0 2308 0 -1 5105
box -2 -3 98 103
use FILL  FILL_50_4_0
timestamp 1607101874
transform -1 0 2412 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_4_1
timestamp 1607101874
transform -1 0 2420 0 -1 5105
box -2 -3 10 103
use AOI21X1  AOI21X1_122
timestamp 1607101874
transform -1 0 2452 0 -1 5105
box -2 -3 34 103
use NOR2X1  NOR2X1_197
timestamp 1607101874
transform 1 0 2452 0 -1 5105
box -2 -3 26 103
use AOI21X1  AOI21X1_125
timestamp 1607101874
transform 1 0 2476 0 -1 5105
box -2 -3 34 103
use NOR2X1  NOR2X1_200
timestamp 1607101874
transform -1 0 2532 0 -1 5105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_962
timestamp 1607101874
transform 1 0 2532 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_451
timestamp 1607101874
transform 1 0 2628 0 -1 5105
box -2 -3 98 103
use NOR2X1  NOR2X1_703
timestamp 1607101874
transform 1 0 2724 0 -1 5105
box -2 -3 26 103
use AOI21X1  AOI21X1_591
timestamp 1607101874
transform -1 0 2780 0 -1 5105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_967
timestamp 1607101874
transform 1 0 2780 0 -1 5105
box -2 -3 98 103
use INVX1  INVX1_127
timestamp 1607101874
transform 1 0 2876 0 -1 5105
box -2 -3 18 103
use FILL  FILL_50_5_0
timestamp 1607101874
transform -1 0 2900 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_5_1
timestamp 1607101874
transform -1 0 2908 0 -1 5105
box -2 -3 10 103
use MUX2X1  MUX2X1_114
timestamp 1607101874
transform -1 0 2956 0 -1 5105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_282
timestamp 1607101874
transform -1 0 3052 0 -1 5105
box -2 -3 98 103
use OAI21X1  OAI21X1_1439
timestamp 1607101874
transform 1 0 3052 0 -1 5105
box -2 -3 34 103
use OAI21X1  OAI21X1_1438
timestamp 1607101874
transform -1 0 3116 0 -1 5105
box -2 -3 34 103
use BUFX4  BUFX4_432
timestamp 1607101874
transform -1 0 3148 0 -1 5105
box -2 -3 34 103
use OAI21X1  OAI21X1_246
timestamp 1607101874
transform 1 0 3148 0 -1 5105
box -2 -3 34 103
use OAI21X1  OAI21X1_247
timestamp 1607101874
transform -1 0 3212 0 -1 5105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_946
timestamp 1607101874
transform -1 0 3308 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_277
timestamp 1607101874
transform 1 0 3308 0 -1 5105
box -2 -3 98 103
use FILL  FILL_50_6_0
timestamp 1607101874
transform 1 0 3404 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_6_1
timestamp 1607101874
transform 1 0 3412 0 -1 5105
box -2 -3 10 103
use INVX1  INVX1_427
timestamp 1607101874
transform 1 0 3420 0 -1 5105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_460
timestamp 1607101874
transform 1 0 3436 0 -1 5105
box -2 -3 98 103
use INVX1  INVX1_316
timestamp 1607101874
transform 1 0 3532 0 -1 5105
box -2 -3 18 103
use MUX2X1  MUX2X1_366
timestamp 1607101874
transform 1 0 3548 0 -1 5105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_456
timestamp 1607101874
transform 1 0 3596 0 -1 5105
box -2 -3 98 103
use MUX2X1  MUX2X1_364
timestamp 1607101874
transform -1 0 3740 0 -1 5105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_450
timestamp 1607101874
transform 1 0 3740 0 -1 5105
box -2 -3 98 103
use INVX1  INVX1_429
timestamp 1607101874
transform 1 0 3836 0 -1 5105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_49
timestamp 1607101874
transform -1 0 3924 0 -1 5105
box -2 -3 74 103
use FILL  FILL_50_7_0
timestamp 1607101874
transform 1 0 3924 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_7_1
timestamp 1607101874
transform 1 0 3932 0 -1 5105
box -2 -3 10 103
use BUFX4  BUFX4_10
timestamp 1607101874
transform 1 0 3940 0 -1 5105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_82
timestamp 1607101874
transform -1 0 4044 0 -1 5105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_467
timestamp 1607101874
transform 1 0 4044 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_477
timestamp 1607101874
transform -1 0 4236 0 -1 5105
box -2 -3 98 103
use INVX1  INVX1_377
timestamp 1607101874
transform 1 0 4236 0 -1 5105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_771
timestamp 1607101874
transform 1 0 4252 0 -1 5105
box -2 -3 98 103
use INVX1  INVX1_69
timestamp 1607101874
transform 1 0 4348 0 -1 5105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_454
timestamp 1607101874
transform 1 0 4364 0 -1 5105
box -2 -3 98 103
use FILL  FILL_50_8_0
timestamp 1607101874
transform -1 0 4468 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_8_1
timestamp 1607101874
transform -1 0 4476 0 -1 5105
box -2 -3 10 103
use INVX1  INVX1_184
timestamp 1607101874
transform -1 0 4492 0 -1 5105
box -2 -3 18 103
use INVX1  INVX1_173
timestamp 1607101874
transform 1 0 4492 0 -1 5105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_628
timestamp 1607101874
transform -1 0 4604 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1607101874
transform -1 0 4700 0 -1 5105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1607101874
transform -1 0 4796 0 -1 5105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_63
timestamp 1607101874
transform -1 0 4868 0 -1 5105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_671
timestamp 1607101874
transform 1 0 4868 0 -1 5105
box -2 -3 98 103
use FILL  FILL_50_9_0
timestamp 1607101874
transform 1 0 4964 0 -1 5105
box -2 -3 10 103
use FILL  FILL_50_9_1
timestamp 1607101874
transform 1 0 4972 0 -1 5105
box -2 -3 10 103
use OAI21X1  OAI21X1_47
timestamp 1607101874
transform 1 0 4980 0 -1 5105
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1607101874
transform -1 0 5028 0 -1 5105
box -2 -3 18 103
use OAI21X1  OAI21X1_722
timestamp 1607101874
transform -1 0 5060 0 -1 5105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_596
timestamp 1607101874
transform 1 0 5060 0 -1 5105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_66
timestamp 1607101874
transform -1 0 5228 0 -1 5105
box -2 -3 74 103
use OAI21X1  OAI21X1_909
timestamp 1607101874
transform 1 0 5228 0 -1 5105
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1607101874
transform 1 0 5260 0 -1 5105
box -2 -3 26 103
use FILL  FILL_51_1
timestamp 1607101874
transform -1 0 5292 0 -1 5105
box -2 -3 10 103
use FILL  FILL_51_2
timestamp 1607101874
transform -1 0 5300 0 -1 5105
box -2 -3 10 103
use FILL  FILL_51_3
timestamp 1607101874
transform -1 0 5308 0 -1 5105
box -2 -3 10 103
<< labels >>
flabel metal6 s 328 -30 344 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 848 -30 864 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 3458 -22 3462 7 FreeSans 24 0 0 0 clock
port 2 nsew
flabel metal3 s -26 4448 -22 4452 7 FreeSans 24 0 0 0 ped_Hori_Interrupt
port 3 nsew
flabel metal2 s 310 5128 314 5132 3 FreeSans 24 90 0 0 ped_Vert_Interrupt
port 4 nsew
flabel metal2 s 1094 5128 1098 5132 3 FreeSans 24 90 0 0 police_Interrupt
port 5 nsew
flabel metal3 s -26 3658 -22 3662 7 FreeSans 24 0 0 0 traffic_Street_0[0]
port 6 nsew
flabel metal3 s -26 3678 -22 3682 7 FreeSans 24 0 0 0 traffic_Street_0[1]
port 7 nsew
flabel metal3 s -26 3778 -22 3782 7 FreeSans 24 0 0 0 traffic_Street_0[2]
port 8 nsew
flabel metal3 s -26 3758 -22 3762 7 FreeSans 24 0 0 0 traffic_Street_0[3]
port 9 nsew
flabel metal2 s 1190 5128 1194 5132 3 FreeSans 24 90 0 0 traffic_Street_1[0]
port 10 nsew
flabel metal2 s 4526 -22 4530 -18 7 FreeSans 24 270 0 0 traffic_Street_1[1]
port 11 nsew
flabel metal3 s -26 3358 -22 3362 7 FreeSans 24 0 0 0 traffic_Street_1[2]
port 12 nsew
flabel metal2 s 1894 5128 1898 5132 3 FreeSans 24 90 0 0 traffic_Street_1[3]
port 13 nsew
flabel metal2 s 2230 -22 2234 -18 7 FreeSans 24 270 0 0 address[0]
port 14 nsew
flabel metal3 s 5334 2648 5338 2652 3 FreeSans 24 0 0 0 address[1]
port 15 nsew
flabel metal3 s 5334 2348 5338 2352 3 FreeSans 24 0 0 0 address[2]
port 16 nsew
flabel metal3 s 5334 2948 5338 2952 3 FreeSans 24 0 0 0 address[3]
port 17 nsew
flabel metal3 s 5334 2248 5338 2252 3 FreeSans 24 0 0 0 address[4]
port 18 nsew
flabel metal3 s 5334 2548 5338 2552 3 FreeSans 24 0 0 0 address[5]
port 19 nsew
flabel metal3 s 5334 2368 5338 2372 3 FreeSans 24 0 0 0 address[6]
port 20 nsew
flabel metal3 s 5334 2408 5338 2412 3 FreeSans 24 0 0 0 read_Write
port 21 nsew
flabel metal3 s 5334 948 5338 952 3 FreeSans 24 0 0 0 enable
port 22 nsew
flabel metal3 s 5334 2388 5338 2392 3 FreeSans 24 0 0 0 street
port 23 nsew
flabel metal2 s 1662 5128 1666 5132 3 FreeSans 24 90 0 0 north_South[0]
port 24 nsew
flabel metal2 s 1550 5128 1554 5132 3 FreeSans 24 90 0 0 north_South[1]
port 25 nsew
flabel metal2 s 1454 5128 1458 5132 3 FreeSans 24 90 0 0 west_East[0]
port 26 nsew
flabel metal2 s 1430 5128 1434 5132 3 FreeSans 24 90 0 0 west_East[1]
port 27 nsew
flabel metal2 s 526 5128 530 5132 3 FreeSans 24 90 0 0 pedestrian_Hori_Street
port 28 nsew
flabel metal2 s 958 5128 962 5132 3 FreeSans 24 90 0 0 pedestrian_Vert_Street
port 29 nsew
flabel metal3 s 5334 48 5338 52 3 FreeSans 24 270 0 0 traffic_Street[0]
port 30 nsew
flabel metal3 s 5334 5048 5338 5052 3 FreeSans 24 90 0 0 traffic_Street[1]
port 31 nsew
flabel metal3 s 5334 2748 5338 2752 3 FreeSans 24 0 0 0 traffic_Street[2]
port 32 nsew
flabel metal3 s 5334 4848 5338 4852 3 FreeSans 24 0 0 0 traffic_Street[3]
port 33 nsew
<< end >>
